// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     May 28 2019 00:54:18

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "Pc2drone" view "INTERFACE"

module Pc2drone (
    uart_input_pc,
    debug_CH5_31B,
    debug_CH3_20A,
    debug_CH0_16A,
    uart_input_drone,
    ppm_output,
    debug_CH6_5B,
    debug_CH2_18A,
    debug_CH4_2A,
    debug_CH1_0A,
    clk_system);

    input uart_input_pc;
    output debug_CH5_31B;
    output debug_CH3_20A;
    output debug_CH0_16A;
    input uart_input_drone;
    output ppm_output;
    output debug_CH6_5B;
    output debug_CH2_18A;
    output debug_CH4_2A;
    output debug_CH1_0A;
    input clk_system;

    wire N__94801;
    wire N__94787;
    wire N__94786;
    wire N__94785;
    wire N__94778;
    wire N__94777;
    wire N__94776;
    wire N__94769;
    wire N__94768;
    wire N__94767;
    wire N__94760;
    wire N__94759;
    wire N__94758;
    wire N__94751;
    wire N__94750;
    wire N__94749;
    wire N__94742;
    wire N__94741;
    wire N__94740;
    wire N__94733;
    wire N__94732;
    wire N__94731;
    wire N__94724;
    wire N__94723;
    wire N__94722;
    wire N__94715;
    wire N__94714;
    wire N__94713;
    wire N__94706;
    wire N__94705;
    wire N__94704;
    wire N__94687;
    wire N__94684;
    wire N__94681;
    wire N__94680;
    wire N__94679;
    wire N__94678;
    wire N__94675;
    wire N__94670;
    wire N__94665;
    wire N__94664;
    wire N__94663;
    wire N__94660;
    wire N__94657;
    wire N__94652;
    wire N__94649;
    wire N__94646;
    wire N__94643;
    wire N__94640;
    wire N__94637;
    wire N__94634;
    wire N__94629;
    wire N__94624;
    wire N__94621;
    wire N__94618;
    wire N__94617;
    wire N__94616;
    wire N__94615;
    wire N__94606;
    wire N__94603;
    wire N__94600;
    wire N__94597;
    wire N__94594;
    wire N__94591;
    wire N__94590;
    wire N__94589;
    wire N__94588;
    wire N__94587;
    wire N__94582;
    wire N__94577;
    wire N__94574;
    wire N__94571;
    wire N__94568;
    wire N__94565;
    wire N__94560;
    wire N__94557;
    wire N__94554;
    wire N__94551;
    wire N__94546;
    wire N__94543;
    wire N__94540;
    wire N__94537;
    wire N__94536;
    wire N__94535;
    wire N__94532;
    wire N__94529;
    wire N__94526;
    wire N__94521;
    wire N__94520;
    wire N__94519;
    wire N__94514;
    wire N__94509;
    wire N__94504;
    wire N__94501;
    wire N__94498;
    wire N__94495;
    wire N__94492;
    wire N__94489;
    wire N__94488;
    wire N__94487;
    wire N__94484;
    wire N__94479;
    wire N__94474;
    wire N__94471;
    wire N__94468;
    wire N__94465;
    wire N__94464;
    wire N__94463;
    wire N__94456;
    wire N__94453;
    wire N__94450;
    wire N__94447;
    wire N__94444;
    wire N__94441;
    wire N__94438;
    wire N__94435;
    wire N__94434;
    wire N__94433;
    wire N__94426;
    wire N__94423;
    wire N__94420;
    wire N__94417;
    wire N__94414;
    wire N__94411;
    wire N__94410;
    wire N__94409;
    wire N__94408;
    wire N__94407;
    wire N__94406;
    wire N__94405;
    wire N__94404;
    wire N__94403;
    wire N__94402;
    wire N__94401;
    wire N__94400;
    wire N__94399;
    wire N__94398;
    wire N__94397;
    wire N__94396;
    wire N__94395;
    wire N__94394;
    wire N__94393;
    wire N__94392;
    wire N__94391;
    wire N__94390;
    wire N__94389;
    wire N__94388;
    wire N__94387;
    wire N__94386;
    wire N__94385;
    wire N__94384;
    wire N__94383;
    wire N__94382;
    wire N__94381;
    wire N__94380;
    wire N__94379;
    wire N__94378;
    wire N__94377;
    wire N__94376;
    wire N__94375;
    wire N__94374;
    wire N__94373;
    wire N__94372;
    wire N__94371;
    wire N__94370;
    wire N__94369;
    wire N__94368;
    wire N__94367;
    wire N__94366;
    wire N__94365;
    wire N__94364;
    wire N__94363;
    wire N__94362;
    wire N__94361;
    wire N__94360;
    wire N__94359;
    wire N__94358;
    wire N__94357;
    wire N__94356;
    wire N__94355;
    wire N__94354;
    wire N__94353;
    wire N__94352;
    wire N__94351;
    wire N__94350;
    wire N__94349;
    wire N__94348;
    wire N__94347;
    wire N__94346;
    wire N__94345;
    wire N__94344;
    wire N__94343;
    wire N__94342;
    wire N__94341;
    wire N__94340;
    wire N__94339;
    wire N__94338;
    wire N__94337;
    wire N__94336;
    wire N__94335;
    wire N__94334;
    wire N__94333;
    wire N__94332;
    wire N__94331;
    wire N__94330;
    wire N__94329;
    wire N__94328;
    wire N__94327;
    wire N__94326;
    wire N__94325;
    wire N__94324;
    wire N__94323;
    wire N__94322;
    wire N__94321;
    wire N__94320;
    wire N__94319;
    wire N__94318;
    wire N__94317;
    wire N__94316;
    wire N__94315;
    wire N__94314;
    wire N__94313;
    wire N__94312;
    wire N__94311;
    wire N__94310;
    wire N__94309;
    wire N__94308;
    wire N__94307;
    wire N__94306;
    wire N__94305;
    wire N__94304;
    wire N__94303;
    wire N__94302;
    wire N__94301;
    wire N__94300;
    wire N__94299;
    wire N__94298;
    wire N__94297;
    wire N__94296;
    wire N__94295;
    wire N__94294;
    wire N__94293;
    wire N__94292;
    wire N__94291;
    wire N__94290;
    wire N__94289;
    wire N__94288;
    wire N__94287;
    wire N__94286;
    wire N__94285;
    wire N__94284;
    wire N__94283;
    wire N__94282;
    wire N__94281;
    wire N__94280;
    wire N__94279;
    wire N__94278;
    wire N__94277;
    wire N__94276;
    wire N__94275;
    wire N__94274;
    wire N__94273;
    wire N__94272;
    wire N__94271;
    wire N__94270;
    wire N__94269;
    wire N__94268;
    wire N__94267;
    wire N__94266;
    wire N__94265;
    wire N__94264;
    wire N__94263;
    wire N__94262;
    wire N__94261;
    wire N__94260;
    wire N__94259;
    wire N__94258;
    wire N__94257;
    wire N__94256;
    wire N__94255;
    wire N__94254;
    wire N__94253;
    wire N__94252;
    wire N__94251;
    wire N__94250;
    wire N__94249;
    wire N__94248;
    wire N__94247;
    wire N__94246;
    wire N__94245;
    wire N__94244;
    wire N__94243;
    wire N__94242;
    wire N__94241;
    wire N__94240;
    wire N__94239;
    wire N__94238;
    wire N__94237;
    wire N__94236;
    wire N__94235;
    wire N__94234;
    wire N__94233;
    wire N__94232;
    wire N__94231;
    wire N__94230;
    wire N__94229;
    wire N__94228;
    wire N__94227;
    wire N__94226;
    wire N__94225;
    wire N__94224;
    wire N__94223;
    wire N__94222;
    wire N__94221;
    wire N__94220;
    wire N__94219;
    wire N__94218;
    wire N__94217;
    wire N__94216;
    wire N__94215;
    wire N__94214;
    wire N__94213;
    wire N__94212;
    wire N__94211;
    wire N__94210;
    wire N__94209;
    wire N__94208;
    wire N__94207;
    wire N__94206;
    wire N__94205;
    wire N__94204;
    wire N__94203;
    wire N__94202;
    wire N__94201;
    wire N__94200;
    wire N__94199;
    wire N__94198;
    wire N__94197;
    wire N__94196;
    wire N__94195;
    wire N__94194;
    wire N__94193;
    wire N__94192;
    wire N__94191;
    wire N__94190;
    wire N__94189;
    wire N__94188;
    wire N__94187;
    wire N__94186;
    wire N__94185;
    wire N__94184;
    wire N__94183;
    wire N__94182;
    wire N__94181;
    wire N__94180;
    wire N__94179;
    wire N__94178;
    wire N__94177;
    wire N__94176;
    wire N__94175;
    wire N__94174;
    wire N__94173;
    wire N__94172;
    wire N__94171;
    wire N__94170;
    wire N__94169;
    wire N__94168;
    wire N__94167;
    wire N__94166;
    wire N__94165;
    wire N__94164;
    wire N__94163;
    wire N__94162;
    wire N__94161;
    wire N__94160;
    wire N__94159;
    wire N__94158;
    wire N__94157;
    wire N__94156;
    wire N__94155;
    wire N__94154;
    wire N__94153;
    wire N__94152;
    wire N__94151;
    wire N__94150;
    wire N__94149;
    wire N__94148;
    wire N__94147;
    wire N__94146;
    wire N__94145;
    wire N__94144;
    wire N__94143;
    wire N__94142;
    wire N__94141;
    wire N__94140;
    wire N__94139;
    wire N__94138;
    wire N__94137;
    wire N__94136;
    wire N__94135;
    wire N__94134;
    wire N__94133;
    wire N__94132;
    wire N__94131;
    wire N__94130;
    wire N__94129;
    wire N__94128;
    wire N__94127;
    wire N__94126;
    wire N__94125;
    wire N__94124;
    wire N__94123;
    wire N__94122;
    wire N__94121;
    wire N__94120;
    wire N__94119;
    wire N__94118;
    wire N__94117;
    wire N__94116;
    wire N__94115;
    wire N__94114;
    wire N__94113;
    wire N__94112;
    wire N__94111;
    wire N__94110;
    wire N__94109;
    wire N__94108;
    wire N__94107;
    wire N__94106;
    wire N__94105;
    wire N__94104;
    wire N__94103;
    wire N__94102;
    wire N__94101;
    wire N__94100;
    wire N__94099;
    wire N__94098;
    wire N__94097;
    wire N__94096;
    wire N__94095;
    wire N__94094;
    wire N__94093;
    wire N__94092;
    wire N__94091;
    wire N__94090;
    wire N__94089;
    wire N__94088;
    wire N__94087;
    wire N__94086;
    wire N__94085;
    wire N__94084;
    wire N__94083;
    wire N__94082;
    wire N__94081;
    wire N__94080;
    wire N__93415;
    wire N__93412;
    wire N__93409;
    wire N__93408;
    wire N__93407;
    wire N__93406;
    wire N__93403;
    wire N__93400;
    wire N__93399;
    wire N__93396;
    wire N__93395;
    wire N__93394;
    wire N__93391;
    wire N__93390;
    wire N__93387;
    wire N__93386;
    wire N__93383;
    wire N__93380;
    wire N__93377;
    wire N__93374;
    wire N__93371;
    wire N__93370;
    wire N__93369;
    wire N__93368;
    wire N__93367;
    wire N__93366;
    wire N__93363;
    wire N__93360;
    wire N__93357;
    wire N__93356;
    wire N__93355;
    wire N__93352;
    wire N__93347;
    wire N__93342;
    wire N__93339;
    wire N__93336;
    wire N__93333;
    wire N__93332;
    wire N__93329;
    wire N__93326;
    wire N__93323;
    wire N__93318;
    wire N__93317;
    wire N__93316;
    wire N__93315;
    wire N__93312;
    wire N__93309;
    wire N__93306;
    wire N__93303;
    wire N__93298;
    wire N__93293;
    wire N__93290;
    wire N__93287;
    wire N__93282;
    wire N__93279;
    wire N__93276;
    wire N__93273;
    wire N__93270;
    wire N__93267;
    wire N__93262;
    wire N__93259;
    wire N__93258;
    wire N__93255;
    wire N__93252;
    wire N__93249;
    wire N__93246;
    wire N__93241;
    wire N__93238;
    wire N__93235;
    wire N__93232;
    wire N__93227;
    wire N__93224;
    wire N__93221;
    wire N__93218;
    wire N__93211;
    wire N__93202;
    wire N__93199;
    wire N__93196;
    wire N__93193;
    wire N__93190;
    wire N__93187;
    wire N__93180;
    wire N__93177;
    wire N__93170;
    wire N__93163;
    wire N__93162;
    wire N__93161;
    wire N__93160;
    wire N__93159;
    wire N__93158;
    wire N__93157;
    wire N__93156;
    wire N__93155;
    wire N__93154;
    wire N__93153;
    wire N__93152;
    wire N__93151;
    wire N__93150;
    wire N__93149;
    wire N__93148;
    wire N__93147;
    wire N__93146;
    wire N__93145;
    wire N__93144;
    wire N__93143;
    wire N__93142;
    wire N__93141;
    wire N__93140;
    wire N__93139;
    wire N__93138;
    wire N__93137;
    wire N__93136;
    wire N__93135;
    wire N__93134;
    wire N__93133;
    wire N__93132;
    wire N__93131;
    wire N__93130;
    wire N__93129;
    wire N__93128;
    wire N__93127;
    wire N__93126;
    wire N__93125;
    wire N__93124;
    wire N__93123;
    wire N__93122;
    wire N__93121;
    wire N__93114;
    wire N__93109;
    wire N__93106;
    wire N__93103;
    wire N__93098;
    wire N__93095;
    wire N__93092;
    wire N__93087;
    wire N__93084;
    wire N__93081;
    wire N__93066;
    wire N__93061;
    wire N__93048;
    wire N__93031;
    wire N__93026;
    wire N__93023;
    wire N__93020;
    wire N__93017;
    wire N__93016;
    wire N__93015;
    wire N__93014;
    wire N__93013;
    wire N__93012;
    wire N__93011;
    wire N__93010;
    wire N__93009;
    wire N__93008;
    wire N__93007;
    wire N__93006;
    wire N__93005;
    wire N__93004;
    wire N__93003;
    wire N__93002;
    wire N__93001;
    wire N__93000;
    wire N__92999;
    wire N__92998;
    wire N__92997;
    wire N__92996;
    wire N__92995;
    wire N__92994;
    wire N__92993;
    wire N__92992;
    wire N__92991;
    wire N__92990;
    wire N__92989;
    wire N__92988;
    wire N__92987;
    wire N__92986;
    wire N__92985;
    wire N__92984;
    wire N__92983;
    wire N__92982;
    wire N__92981;
    wire N__92980;
    wire N__92979;
    wire N__92978;
    wire N__92977;
    wire N__92976;
    wire N__92975;
    wire N__92974;
    wire N__92973;
    wire N__92972;
    wire N__92971;
    wire N__92970;
    wire N__92969;
    wire N__92968;
    wire N__92967;
    wire N__92966;
    wire N__92965;
    wire N__92962;
    wire N__92959;
    wire N__92956;
    wire N__92953;
    wire N__92950;
    wire N__92947;
    wire N__92944;
    wire N__92941;
    wire N__92938;
    wire N__92935;
    wire N__92932;
    wire N__92929;
    wire N__92926;
    wire N__92923;
    wire N__92920;
    wire N__92917;
    wire N__92914;
    wire N__92911;
    wire N__92770;
    wire N__92767;
    wire N__92764;
    wire N__92761;
    wire N__92758;
    wire N__92755;
    wire N__92754;
    wire N__92751;
    wire N__92748;
    wire N__92747;
    wire N__92744;
    wire N__92741;
    wire N__92738;
    wire N__92733;
    wire N__92730;
    wire N__92727;
    wire N__92724;
    wire N__92719;
    wire N__92716;
    wire N__92713;
    wire N__92710;
    wire N__92709;
    wire N__92708;
    wire N__92701;
    wire N__92698;
    wire N__92695;
    wire N__92692;
    wire N__92689;
    wire N__92686;
    wire N__92683;
    wire N__92682;
    wire N__92679;
    wire N__92678;
    wire N__92677;
    wire N__92676;
    wire N__92673;
    wire N__92672;
    wire N__92669;
    wire N__92666;
    wire N__92665;
    wire N__92662;
    wire N__92661;
    wire N__92658;
    wire N__92657;
    wire N__92656;
    wire N__92655;
    wire N__92652;
    wire N__92651;
    wire N__92650;
    wire N__92649;
    wire N__92646;
    wire N__92641;
    wire N__92638;
    wire N__92635;
    wire N__92632;
    wire N__92629;
    wire N__92626;
    wire N__92623;
    wire N__92620;
    wire N__92619;
    wire N__92616;
    wire N__92613;
    wire N__92610;
    wire N__92607;
    wire N__92604;
    wire N__92601;
    wire N__92598;
    wire N__92591;
    wire N__92586;
    wire N__92583;
    wire N__92580;
    wire N__92577;
    wire N__92574;
    wire N__92567;
    wire N__92564;
    wire N__92561;
    wire N__92552;
    wire N__92545;
    wire N__92540;
    wire N__92537;
    wire N__92534;
    wire N__92531;
    wire N__92528;
    wire N__92521;
    wire N__92520;
    wire N__92519;
    wire N__92518;
    wire N__92517;
    wire N__92516;
    wire N__92515;
    wire N__92514;
    wire N__92513;
    wire N__92510;
    wire N__92509;
    wire N__92506;
    wire N__92503;
    wire N__92500;
    wire N__92495;
    wire N__92494;
    wire N__92491;
    wire N__92488;
    wire N__92485;
    wire N__92482;
    wire N__92479;
    wire N__92476;
    wire N__92475;
    wire N__92474;
    wire N__92471;
    wire N__92466;
    wire N__92465;
    wire N__92462;
    wire N__92459;
    wire N__92454;
    wire N__92451;
    wire N__92448;
    wire N__92445;
    wire N__92442;
    wire N__92439;
    wire N__92436;
    wire N__92433;
    wire N__92432;
    wire N__92431;
    wire N__92430;
    wire N__92427;
    wire N__92420;
    wire N__92417;
    wire N__92414;
    wire N__92411;
    wire N__92408;
    wire N__92405;
    wire N__92400;
    wire N__92393;
    wire N__92392;
    wire N__92391;
    wire N__92384;
    wire N__92377;
    wire N__92370;
    wire N__92365;
    wire N__92356;
    wire N__92355;
    wire N__92352;
    wire N__92349;
    wire N__92346;
    wire N__92343;
    wire N__92340;
    wire N__92337;
    wire N__92332;
    wire N__92331;
    wire N__92330;
    wire N__92329;
    wire N__92328;
    wire N__92327;
    wire N__92326;
    wire N__92323;
    wire N__92322;
    wire N__92321;
    wire N__92320;
    wire N__92319;
    wire N__92316;
    wire N__92313;
    wire N__92308;
    wire N__92305;
    wire N__92302;
    wire N__92301;
    wire N__92298;
    wire N__92295;
    wire N__92288;
    wire N__92287;
    wire N__92284;
    wire N__92283;
    wire N__92280;
    wire N__92279;
    wire N__92276;
    wire N__92273;
    wire N__92270;
    wire N__92267;
    wire N__92264;
    wire N__92259;
    wire N__92256;
    wire N__92253;
    wire N__92250;
    wire N__92247;
    wire N__92244;
    wire N__92239;
    wire N__92236;
    wire N__92235;
    wire N__92234;
    wire N__92231;
    wire N__92228;
    wire N__92225;
    wire N__92222;
    wire N__92219;
    wire N__92216;
    wire N__92213;
    wire N__92208;
    wire N__92205;
    wire N__92200;
    wire N__92193;
    wire N__92192;
    wire N__92191;
    wire N__92188;
    wire N__92183;
    wire N__92178;
    wire N__92173;
    wire N__92170;
    wire N__92165;
    wire N__92152;
    wire N__92151;
    wire N__92148;
    wire N__92145;
    wire N__92142;
    wire N__92139;
    wire N__92134;
    wire N__92131;
    wire N__92128;
    wire N__92127;
    wire N__92126;
    wire N__92125;
    wire N__92124;
    wire N__92123;
    wire N__92122;
    wire N__92119;
    wire N__92116;
    wire N__92113;
    wire N__92110;
    wire N__92107;
    wire N__92104;
    wire N__92103;
    wire N__92102;
    wire N__92101;
    wire N__92098;
    wire N__92093;
    wire N__92090;
    wire N__92087;
    wire N__92084;
    wire N__92081;
    wire N__92078;
    wire N__92075;
    wire N__92072;
    wire N__92071;
    wire N__92070;
    wire N__92067;
    wire N__92066;
    wire N__92065;
    wire N__92062;
    wire N__92059;
    wire N__92056;
    wire N__92053;
    wire N__92052;
    wire N__92047;
    wire N__92042;
    wire N__92041;
    wire N__92038;
    wire N__92035;
    wire N__92032;
    wire N__92029;
    wire N__92026;
    wire N__92023;
    wire N__92018;
    wire N__92015;
    wire N__92012;
    wire N__92009;
    wire N__92006;
    wire N__92003;
    wire N__92000;
    wire N__91997;
    wire N__91992;
    wire N__91989;
    wire N__91982;
    wire N__91973;
    wire N__91966;
    wire N__91957;
    wire N__91956;
    wire N__91953;
    wire N__91950;
    wire N__91947;
    wire N__91944;
    wire N__91939;
    wire N__91936;
    wire N__91933;
    wire N__91932;
    wire N__91929;
    wire N__91928;
    wire N__91925;
    wire N__91924;
    wire N__91921;
    wire N__91918;
    wire N__91917;
    wire N__91914;
    wire N__91911;
    wire N__91908;
    wire N__91905;
    wire N__91902;
    wire N__91897;
    wire N__91892;
    wire N__91889;
    wire N__91886;
    wire N__91883;
    wire N__91878;
    wire N__91875;
    wire N__91870;
    wire N__91867;
    wire N__91864;
    wire N__91861;
    wire N__91858;
    wire N__91857;
    wire N__91856;
    wire N__91853;
    wire N__91848;
    wire N__91845;
    wire N__91842;
    wire N__91837;
    wire N__91834;
    wire N__91831;
    wire N__91828;
    wire N__91825;
    wire N__91822;
    wire N__91819;
    wire N__91816;
    wire N__91813;
    wire N__91812;
    wire N__91811;
    wire N__91808;
    wire N__91803;
    wire N__91798;
    wire N__91795;
    wire N__91792;
    wire N__91789;
    wire N__91786;
    wire N__91783;
    wire N__91780;
    wire N__91779;
    wire N__91776;
    wire N__91775;
    wire N__91774;
    wire N__91773;
    wire N__91766;
    wire N__91763;
    wire N__91760;
    wire N__91759;
    wire N__91758;
    wire N__91757;
    wire N__91756;
    wire N__91755;
    wire N__91754;
    wire N__91751;
    wire N__91748;
    wire N__91741;
    wire N__91740;
    wire N__91737;
    wire N__91734;
    wire N__91731;
    wire N__91730;
    wire N__91727;
    wire N__91720;
    wire N__91719;
    wire N__91718;
    wire N__91717;
    wire N__91714;
    wire N__91711;
    wire N__91704;
    wire N__91699;
    wire N__91692;
    wire N__91685;
    wire N__91682;
    wire N__91679;
    wire N__91676;
    wire N__91673;
    wire N__91670;
    wire N__91667;
    wire N__91660;
    wire N__91657;
    wire N__91654;
    wire N__91651;
    wire N__91650;
    wire N__91649;
    wire N__91648;
    wire N__91647;
    wire N__91646;
    wire N__91645;
    wire N__91644;
    wire N__91643;
    wire N__91642;
    wire N__91641;
    wire N__91640;
    wire N__91639;
    wire N__91632;
    wire N__91627;
    wire N__91626;
    wire N__91625;
    wire N__91622;
    wire N__91613;
    wire N__91606;
    wire N__91601;
    wire N__91596;
    wire N__91595;
    wire N__91594;
    wire N__91591;
    wire N__91588;
    wire N__91581;
    wire N__91576;
    wire N__91571;
    wire N__91568;
    wire N__91565;
    wire N__91560;
    wire N__91557;
    wire N__91552;
    wire N__91549;
    wire N__91546;
    wire N__91543;
    wire N__91540;
    wire N__91539;
    wire N__91538;
    wire N__91531;
    wire N__91528;
    wire N__91525;
    wire N__91522;
    wire N__91519;
    wire N__91518;
    wire N__91515;
    wire N__91512;
    wire N__91509;
    wire N__91506;
    wire N__91503;
    wire N__91500;
    wire N__91495;
    wire N__91494;
    wire N__91489;
    wire N__91488;
    wire N__91485;
    wire N__91484;
    wire N__91483;
    wire N__91482;
    wire N__91481;
    wire N__91478;
    wire N__91475;
    wire N__91466;
    wire N__91459;
    wire N__91456;
    wire N__91453;
    wire N__91450;
    wire N__91447;
    wire N__91444;
    wire N__91441;
    wire N__91438;
    wire N__91437;
    wire N__91436;
    wire N__91433;
    wire N__91432;
    wire N__91431;
    wire N__91428;
    wire N__91425;
    wire N__91422;
    wire N__91417;
    wire N__91412;
    wire N__91407;
    wire N__91404;
    wire N__91401;
    wire N__91396;
    wire N__91393;
    wire N__91390;
    wire N__91387;
    wire N__91384;
    wire N__91383;
    wire N__91382;
    wire N__91381;
    wire N__91380;
    wire N__91379;
    wire N__91378;
    wire N__91377;
    wire N__91376;
    wire N__91375;
    wire N__91374;
    wire N__91371;
    wire N__91370;
    wire N__91363;
    wire N__91358;
    wire N__91357;
    wire N__91354;
    wire N__91347;
    wire N__91344;
    wire N__91339;
    wire N__91334;
    wire N__91331;
    wire N__91330;
    wire N__91329;
    wire N__91328;
    wire N__91325;
    wire N__91320;
    wire N__91317;
    wire N__91314;
    wire N__91305;
    wire N__91300;
    wire N__91297;
    wire N__91294;
    wire N__91291;
    wire N__91286;
    wire N__91283;
    wire N__91280;
    wire N__91277;
    wire N__91270;
    wire N__91267;
    wire N__91264;
    wire N__91263;
    wire N__91260;
    wire N__91257;
    wire N__91252;
    wire N__91249;
    wire N__91248;
    wire N__91247;
    wire N__91246;
    wire N__91245;
    wire N__91244;
    wire N__91243;
    wire N__91240;
    wire N__91239;
    wire N__91238;
    wire N__91233;
    wire N__91226;
    wire N__91223;
    wire N__91220;
    wire N__91215;
    wire N__91210;
    wire N__91207;
    wire N__91204;
    wire N__91199;
    wire N__91196;
    wire N__91193;
    wire N__91190;
    wire N__91183;
    wire N__91180;
    wire N__91177;
    wire N__91174;
    wire N__91171;
    wire N__91170;
    wire N__91169;
    wire N__91166;
    wire N__91161;
    wire N__91158;
    wire N__91155;
    wire N__91152;
    wire N__91149;
    wire N__91146;
    wire N__91141;
    wire N__91138;
    wire N__91135;
    wire N__91132;
    wire N__91129;
    wire N__91128;
    wire N__91127;
    wire N__91122;
    wire N__91119;
    wire N__91116;
    wire N__91113;
    wire N__91110;
    wire N__91107;
    wire N__91104;
    wire N__91099;
    wire N__91096;
    wire N__91093;
    wire N__91090;
    wire N__91087;
    wire N__91086;
    wire N__91085;
    wire N__91078;
    wire N__91075;
    wire N__91072;
    wire N__91069;
    wire N__91066;
    wire N__91063;
    wire N__91060;
    wire N__91057;
    wire N__91054;
    wire N__91051;
    wire N__91050;
    wire N__91045;
    wire N__91042;
    wire N__91039;
    wire N__91036;
    wire N__91033;
    wire N__91030;
    wire N__91027;
    wire N__91026;
    wire N__91025;
    wire N__91022;
    wire N__91021;
    wire N__91020;
    wire N__91017;
    wire N__91014;
    wire N__91007;
    wire N__91004;
    wire N__90997;
    wire N__90994;
    wire N__90991;
    wire N__90988;
    wire N__90985;
    wire N__90982;
    wire N__90979;
    wire N__90978;
    wire N__90975;
    wire N__90974;
    wire N__90973;
    wire N__90972;
    wire N__90969;
    wire N__90968;
    wire N__90967;
    wire N__90964;
    wire N__90961;
    wire N__90958;
    wire N__90955;
    wire N__90948;
    wire N__90945;
    wire N__90936;
    wire N__90931;
    wire N__90928;
    wire N__90925;
    wire N__90922;
    wire N__90919;
    wire N__90918;
    wire N__90917;
    wire N__90912;
    wire N__90911;
    wire N__90908;
    wire N__90907;
    wire N__90904;
    wire N__90901;
    wire N__90900;
    wire N__90899;
    wire N__90898;
    wire N__90893;
    wire N__90890;
    wire N__90887;
    wire N__90880;
    wire N__90877;
    wire N__90870;
    wire N__90865;
    wire N__90862;
    wire N__90859;
    wire N__90856;
    wire N__90855;
    wire N__90852;
    wire N__90851;
    wire N__90848;
    wire N__90847;
    wire N__90844;
    wire N__90841;
    wire N__90836;
    wire N__90833;
    wire N__90828;
    wire N__90823;
    wire N__90820;
    wire N__90817;
    wire N__90814;
    wire N__90813;
    wire N__90808;
    wire N__90805;
    wire N__90802;
    wire N__90799;
    wire N__90796;
    wire N__90793;
    wire N__90790;
    wire N__90789;
    wire N__90786;
    wire N__90783;
    wire N__90780;
    wire N__90777;
    wire N__90774;
    wire N__90771;
    wire N__90768;
    wire N__90765;
    wire N__90762;
    wire N__90759;
    wire N__90754;
    wire N__90751;
    wire N__90748;
    wire N__90745;
    wire N__90744;
    wire N__90741;
    wire N__90738;
    wire N__90735;
    wire N__90732;
    wire N__90727;
    wire N__90724;
    wire N__90721;
    wire N__90718;
    wire N__90715;
    wire N__90714;
    wire N__90713;
    wire N__90710;
    wire N__90707;
    wire N__90704;
    wire N__90701;
    wire N__90696;
    wire N__90693;
    wire N__90690;
    wire N__90685;
    wire N__90682;
    wire N__90681;
    wire N__90678;
    wire N__90677;
    wire N__90676;
    wire N__90675;
    wire N__90672;
    wire N__90671;
    wire N__90670;
    wire N__90669;
    wire N__90668;
    wire N__90667;
    wire N__90664;
    wire N__90663;
    wire N__90662;
    wire N__90659;
    wire N__90658;
    wire N__90657;
    wire N__90654;
    wire N__90653;
    wire N__90650;
    wire N__90649;
    wire N__90648;
    wire N__90647;
    wire N__90646;
    wire N__90645;
    wire N__90642;
    wire N__90639;
    wire N__90636;
    wire N__90629;
    wire N__90626;
    wire N__90623;
    wire N__90620;
    wire N__90617;
    wire N__90614;
    wire N__90613;
    wire N__90610;
    wire N__90607;
    wire N__90604;
    wire N__90601;
    wire N__90600;
    wire N__90597;
    wire N__90594;
    wire N__90591;
    wire N__90588;
    wire N__90585;
    wire N__90582;
    wire N__90579;
    wire N__90574;
    wire N__90567;
    wire N__90564;
    wire N__90561;
    wire N__90558;
    wire N__90555;
    wire N__90552;
    wire N__90549;
    wire N__90546;
    wire N__90545;
    wire N__90544;
    wire N__90539;
    wire N__90536;
    wire N__90533;
    wire N__90530;
    wire N__90527;
    wire N__90518;
    wire N__90515;
    wire N__90512;
    wire N__90509;
    wire N__90506;
    wire N__90499;
    wire N__90498;
    wire N__90495;
    wire N__90492;
    wire N__90489;
    wire N__90486;
    wire N__90477;
    wire N__90468;
    wire N__90465;
    wire N__90460;
    wire N__90451;
    wire N__90442;
    wire N__90441;
    wire N__90438;
    wire N__90437;
    wire N__90436;
    wire N__90435;
    wire N__90434;
    wire N__90433;
    wire N__90432;
    wire N__90431;
    wire N__90428;
    wire N__90427;
    wire N__90420;
    wire N__90419;
    wire N__90416;
    wire N__90413;
    wire N__90412;
    wire N__90409;
    wire N__90408;
    wire N__90405;
    wire N__90404;
    wire N__90401;
    wire N__90398;
    wire N__90397;
    wire N__90396;
    wire N__90395;
    wire N__90392;
    wire N__90389;
    wire N__90386;
    wire N__90383;
    wire N__90380;
    wire N__90379;
    wire N__90378;
    wire N__90377;
    wire N__90376;
    wire N__90373;
    wire N__90370;
    wire N__90367;
    wire N__90364;
    wire N__90361;
    wire N__90356;
    wire N__90351;
    wire N__90348;
    wire N__90347;
    wire N__90344;
    wire N__90343;
    wire N__90336;
    wire N__90333;
    wire N__90324;
    wire N__90321;
    wire N__90318;
    wire N__90315;
    wire N__90310;
    wire N__90303;
    wire N__90302;
    wire N__90299;
    wire N__90296;
    wire N__90293;
    wire N__90288;
    wire N__90283;
    wire N__90274;
    wire N__90269;
    wire N__90256;
    wire N__90255;
    wire N__90254;
    wire N__90253;
    wire N__90252;
    wire N__90251;
    wire N__90248;
    wire N__90247;
    wire N__90244;
    wire N__90241;
    wire N__90240;
    wire N__90239;
    wire N__90236;
    wire N__90235;
    wire N__90234;
    wire N__90231;
    wire N__90224;
    wire N__90223;
    wire N__90222;
    wire N__90221;
    wire N__90220;
    wire N__90217;
    wire N__90212;
    wire N__90211;
    wire N__90208;
    wire N__90207;
    wire N__90204;
    wire N__90201;
    wire N__90198;
    wire N__90193;
    wire N__90190;
    wire N__90185;
    wire N__90182;
    wire N__90181;
    wire N__90178;
    wire N__90175;
    wire N__90168;
    wire N__90163;
    wire N__90160;
    wire N__90157;
    wire N__90156;
    wire N__90151;
    wire N__90146;
    wire N__90139;
    wire N__90132;
    wire N__90131;
    wire N__90130;
    wire N__90127;
    wire N__90126;
    wire N__90123;
    wire N__90120;
    wire N__90117;
    wire N__90114;
    wire N__90109;
    wire N__90106;
    wire N__90103;
    wire N__90094;
    wire N__90089;
    wire N__90082;
    wire N__90079;
    wire N__90078;
    wire N__90075;
    wire N__90072;
    wire N__90069;
    wire N__90066;
    wire N__90063;
    wire N__90060;
    wire N__90055;
    wire N__90052;
    wire N__90049;
    wire N__90046;
    wire N__90045;
    wire N__90040;
    wire N__90037;
    wire N__90034;
    wire N__90031;
    wire N__90028;
    wire N__90025;
    wire N__90022;
    wire N__90019;
    wire N__90016;
    wire N__90015;
    wire N__90014;
    wire N__90011;
    wire N__90008;
    wire N__90005;
    wire N__90002;
    wire N__89999;
    wire N__89996;
    wire N__89993;
    wire N__89988;
    wire N__89983;
    wire N__89980;
    wire N__89977;
    wire N__89974;
    wire N__89971;
    wire N__89970;
    wire N__89967;
    wire N__89962;
    wire N__89959;
    wire N__89956;
    wire N__89953;
    wire N__89950;
    wire N__89947;
    wire N__89944;
    wire N__89941;
    wire N__89940;
    wire N__89937;
    wire N__89934;
    wire N__89931;
    wire N__89928;
    wire N__89923;
    wire N__89920;
    wire N__89917;
    wire N__89914;
    wire N__89911;
    wire N__89908;
    wire N__89905;
    wire N__89902;
    wire N__89901;
    wire N__89898;
    wire N__89895;
    wire N__89890;
    wire N__89887;
    wire N__89884;
    wire N__89881;
    wire N__89878;
    wire N__89875;
    wire N__89874;
    wire N__89871;
    wire N__89868;
    wire N__89863;
    wire N__89860;
    wire N__89857;
    wire N__89854;
    wire N__89851;
    wire N__89850;
    wire N__89849;
    wire N__89846;
    wire N__89843;
    wire N__89842;
    wire N__89839;
    wire N__89838;
    wire N__89837;
    wire N__89834;
    wire N__89829;
    wire N__89828;
    wire N__89823;
    wire N__89822;
    wire N__89821;
    wire N__89820;
    wire N__89819;
    wire N__89818;
    wire N__89817;
    wire N__89816;
    wire N__89815;
    wire N__89812;
    wire N__89807;
    wire N__89804;
    wire N__89801;
    wire N__89798;
    wire N__89795;
    wire N__89794;
    wire N__89793;
    wire N__89790;
    wire N__89789;
    wire N__89788;
    wire N__89787;
    wire N__89784;
    wire N__89781;
    wire N__89778;
    wire N__89775;
    wire N__89772;
    wire N__89767;
    wire N__89762;
    wire N__89759;
    wire N__89756;
    wire N__89755;
    wire N__89752;
    wire N__89749;
    wire N__89748;
    wire N__89747;
    wire N__89746;
    wire N__89743;
    wire N__89740;
    wire N__89737;
    wire N__89734;
    wire N__89731;
    wire N__89730;
    wire N__89727;
    wire N__89724;
    wire N__89721;
    wire N__89718;
    wire N__89711;
    wire N__89708;
    wire N__89705;
    wire N__89700;
    wire N__89697;
    wire N__89696;
    wire N__89693;
    wire N__89692;
    wire N__89689;
    wire N__89686;
    wire N__89683;
    wire N__89678;
    wire N__89675;
    wire N__89672;
    wire N__89665;
    wire N__89658;
    wire N__89655;
    wire N__89652;
    wire N__89649;
    wire N__89640;
    wire N__89635;
    wire N__89628;
    wire N__89623;
    wire N__89618;
    wire N__89605;
    wire N__89604;
    wire N__89603;
    wire N__89602;
    wire N__89601;
    wire N__89598;
    wire N__89593;
    wire N__89592;
    wire N__89591;
    wire N__89590;
    wire N__89587;
    wire N__89586;
    wire N__89583;
    wire N__89580;
    wire N__89577;
    wire N__89576;
    wire N__89573;
    wire N__89572;
    wire N__89569;
    wire N__89564;
    wire N__89563;
    wire N__89562;
    wire N__89559;
    wire N__89556;
    wire N__89553;
    wire N__89550;
    wire N__89547;
    wire N__89544;
    wire N__89541;
    wire N__89536;
    wire N__89535;
    wire N__89532;
    wire N__89531;
    wire N__89530;
    wire N__89527;
    wire N__89526;
    wire N__89525;
    wire N__89522;
    wire N__89521;
    wire N__89518;
    wire N__89509;
    wire N__89508;
    wire N__89503;
    wire N__89502;
    wire N__89499;
    wire N__89496;
    wire N__89495;
    wire N__89494;
    wire N__89491;
    wire N__89488;
    wire N__89485;
    wire N__89480;
    wire N__89477;
    wire N__89474;
    wire N__89469;
    wire N__89468;
    wire N__89465;
    wire N__89462;
    wire N__89459;
    wire N__89454;
    wire N__89451;
    wire N__89444;
    wire N__89439;
    wire N__89438;
    wire N__89437;
    wire N__89436;
    wire N__89433;
    wire N__89430;
    wire N__89427;
    wire N__89422;
    wire N__89411;
    wire N__89408;
    wire N__89405;
    wire N__89400;
    wire N__89391;
    wire N__89386;
    wire N__89377;
    wire N__89376;
    wire N__89375;
    wire N__89374;
    wire N__89373;
    wire N__89372;
    wire N__89369;
    wire N__89366;
    wire N__89363;
    wire N__89360;
    wire N__89355;
    wire N__89354;
    wire N__89353;
    wire N__89352;
    wire N__89351;
    wire N__89348;
    wire N__89347;
    wire N__89346;
    wire N__89345;
    wire N__89342;
    wire N__89339;
    wire N__89338;
    wire N__89335;
    wire N__89334;
    wire N__89331;
    wire N__89324;
    wire N__89321;
    wire N__89320;
    wire N__89317;
    wire N__89312;
    wire N__89311;
    wire N__89308;
    wire N__89307;
    wire N__89306;
    wire N__89301;
    wire N__89300;
    wire N__89297;
    wire N__89294;
    wire N__89293;
    wire N__89292;
    wire N__89291;
    wire N__89288;
    wire N__89287;
    wire N__89286;
    wire N__89281;
    wire N__89278;
    wire N__89275;
    wire N__89270;
    wire N__89267;
    wire N__89264;
    wire N__89259;
    wire N__89256;
    wire N__89253;
    wire N__89252;
    wire N__89247;
    wire N__89246;
    wire N__89245;
    wire N__89242;
    wire N__89239;
    wire N__89234;
    wire N__89233;
    wire N__89232;
    wire N__89229;
    wire N__89226;
    wire N__89223;
    wire N__89216;
    wire N__89213;
    wire N__89204;
    wire N__89201;
    wire N__89198;
    wire N__89193;
    wire N__89188;
    wire N__89185;
    wire N__89182;
    wire N__89179;
    wire N__89172;
    wire N__89169;
    wire N__89164;
    wire N__89163;
    wire N__89156;
    wire N__89149;
    wire N__89144;
    wire N__89139;
    wire N__89136;
    wire N__89133;
    wire N__89130;
    wire N__89127;
    wire N__89124;
    wire N__89113;
    wire N__89112;
    wire N__89111;
    wire N__89110;
    wire N__89109;
    wire N__89106;
    wire N__89103;
    wire N__89100;
    wire N__89099;
    wire N__89098;
    wire N__89097;
    wire N__89094;
    wire N__89091;
    wire N__89088;
    wire N__89083;
    wire N__89082;
    wire N__89081;
    wire N__89080;
    wire N__89079;
    wire N__89078;
    wire N__89077;
    wire N__89074;
    wire N__89073;
    wire N__89072;
    wire N__89069;
    wire N__89068;
    wire N__89067;
    wire N__89066;
    wire N__89065;
    wire N__89062;
    wire N__89059;
    wire N__89054;
    wire N__89051;
    wire N__89044;
    wire N__89043;
    wire N__89038;
    wire N__89037;
    wire N__89034;
    wire N__89029;
    wire N__89028;
    wire N__89027;
    wire N__89024;
    wire N__89021;
    wire N__89016;
    wire N__89011;
    wire N__89004;
    wire N__88999;
    wire N__88996;
    wire N__88993;
    wire N__88990;
    wire N__88985;
    wire N__88984;
    wire N__88981;
    wire N__88976;
    wire N__88973;
    wire N__88972;
    wire N__88971;
    wire N__88966;
    wire N__88961;
    wire N__88958;
    wire N__88951;
    wire N__88948;
    wire N__88943;
    wire N__88940;
    wire N__88937;
    wire N__88934;
    wire N__88931;
    wire N__88928;
    wire N__88923;
    wire N__88920;
    wire N__88917;
    wire N__88912;
    wire N__88905;
    wire N__88902;
    wire N__88895;
    wire N__88888;
    wire N__88885;
    wire N__88882;
    wire N__88881;
    wire N__88878;
    wire N__88875;
    wire N__88872;
    wire N__88869;
    wire N__88864;
    wire N__88861;
    wire N__88860;
    wire N__88859;
    wire N__88858;
    wire N__88855;
    wire N__88854;
    wire N__88851;
    wire N__88848;
    wire N__88847;
    wire N__88846;
    wire N__88843;
    wire N__88840;
    wire N__88837;
    wire N__88834;
    wire N__88831;
    wire N__88830;
    wire N__88829;
    wire N__88828;
    wire N__88825;
    wire N__88822;
    wire N__88817;
    wire N__88814;
    wire N__88813;
    wire N__88810;
    wire N__88807;
    wire N__88802;
    wire N__88799;
    wire N__88798;
    wire N__88795;
    wire N__88792;
    wire N__88789;
    wire N__88786;
    wire N__88783;
    wire N__88778;
    wire N__88775;
    wire N__88772;
    wire N__88769;
    wire N__88768;
    wire N__88767;
    wire N__88762;
    wire N__88759;
    wire N__88756;
    wire N__88751;
    wire N__88744;
    wire N__88739;
    wire N__88726;
    wire N__88723;
    wire N__88722;
    wire N__88719;
    wire N__88716;
    wire N__88713;
    wire N__88710;
    wire N__88705;
    wire N__88702;
    wire N__88701;
    wire N__88700;
    wire N__88699;
    wire N__88696;
    wire N__88695;
    wire N__88692;
    wire N__88689;
    wire N__88686;
    wire N__88685;
    wire N__88682;
    wire N__88679;
    wire N__88676;
    wire N__88673;
    wire N__88670;
    wire N__88667;
    wire N__88666;
    wire N__88665;
    wire N__88664;
    wire N__88663;
    wire N__88658;
    wire N__88655;
    wire N__88650;
    wire N__88647;
    wire N__88646;
    wire N__88643;
    wire N__88642;
    wire N__88641;
    wire N__88640;
    wire N__88637;
    wire N__88636;
    wire N__88633;
    wire N__88630;
    wire N__88627;
    wire N__88624;
    wire N__88621;
    wire N__88618;
    wire N__88615;
    wire N__88612;
    wire N__88607;
    wire N__88604;
    wire N__88601;
    wire N__88598;
    wire N__88595;
    wire N__88588;
    wire N__88585;
    wire N__88580;
    wire N__88575;
    wire N__88574;
    wire N__88571;
    wire N__88568;
    wire N__88563;
    wire N__88560;
    wire N__88555;
    wire N__88552;
    wire N__88549;
    wire N__88534;
    wire N__88531;
    wire N__88530;
    wire N__88527;
    wire N__88524;
    wire N__88521;
    wire N__88518;
    wire N__88513;
    wire N__88510;
    wire N__88509;
    wire N__88508;
    wire N__88507;
    wire N__88506;
    wire N__88505;
    wire N__88502;
    wire N__88499;
    wire N__88496;
    wire N__88493;
    wire N__88490;
    wire N__88489;
    wire N__88486;
    wire N__88483;
    wire N__88482;
    wire N__88481;
    wire N__88480;
    wire N__88477;
    wire N__88474;
    wire N__88471;
    wire N__88470;
    wire N__88467;
    wire N__88464;
    wire N__88461;
    wire N__88458;
    wire N__88457;
    wire N__88454;
    wire N__88451;
    wire N__88448;
    wire N__88445;
    wire N__88440;
    wire N__88437;
    wire N__88434;
    wire N__88431;
    wire N__88426;
    wire N__88425;
    wire N__88422;
    wire N__88419;
    wire N__88416;
    wire N__88413;
    wire N__88410;
    wire N__88407;
    wire N__88404;
    wire N__88401;
    wire N__88396;
    wire N__88393;
    wire N__88392;
    wire N__88389;
    wire N__88386;
    wire N__88381;
    wire N__88378;
    wire N__88375;
    wire N__88366;
    wire N__88363;
    wire N__88348;
    wire N__88345;
    wire N__88344;
    wire N__88341;
    wire N__88338;
    wire N__88335;
    wire N__88332;
    wire N__88327;
    wire N__88324;
    wire N__88323;
    wire N__88322;
    wire N__88321;
    wire N__88320;
    wire N__88317;
    wire N__88314;
    wire N__88311;
    wire N__88308;
    wire N__88307;
    wire N__88306;
    wire N__88305;
    wire N__88302;
    wire N__88297;
    wire N__88294;
    wire N__88291;
    wire N__88288;
    wire N__88285;
    wire N__88282;
    wire N__88281;
    wire N__88280;
    wire N__88275;
    wire N__88270;
    wire N__88267;
    wire N__88264;
    wire N__88263;
    wire N__88262;
    wire N__88261;
    wire N__88260;
    wire N__88257;
    wire N__88256;
    wire N__88255;
    wire N__88254;
    wire N__88251;
    wire N__88248;
    wire N__88245;
    wire N__88242;
    wire N__88239;
    wire N__88236;
    wire N__88231;
    wire N__88228;
    wire N__88225;
    wire N__88222;
    wire N__88219;
    wire N__88216;
    wire N__88213;
    wire N__88210;
    wire N__88207;
    wire N__88202;
    wire N__88195;
    wire N__88194;
    wire N__88191;
    wire N__88186;
    wire N__88183;
    wire N__88180;
    wire N__88175;
    wire N__88170;
    wire N__88167;
    wire N__88164;
    wire N__88157;
    wire N__88144;
    wire N__88141;
    wire N__88140;
    wire N__88137;
    wire N__88134;
    wire N__88131;
    wire N__88128;
    wire N__88123;
    wire N__88120;
    wire N__88119;
    wire N__88116;
    wire N__88113;
    wire N__88108;
    wire N__88107;
    wire N__88106;
    wire N__88103;
    wire N__88100;
    wire N__88097;
    wire N__88092;
    wire N__88091;
    wire N__88090;
    wire N__88089;
    wire N__88088;
    wire N__88087;
    wire N__88084;
    wire N__88081;
    wire N__88080;
    wire N__88079;
    wire N__88078;
    wire N__88075;
    wire N__88072;
    wire N__88069;
    wire N__88066;
    wire N__88063;
    wire N__88058;
    wire N__88055;
    wire N__88054;
    wire N__88053;
    wire N__88050;
    wire N__88047;
    wire N__88044;
    wire N__88041;
    wire N__88038;
    wire N__88035;
    wire N__88032;
    wire N__88027;
    wire N__88024;
    wire N__88021;
    wire N__88020;
    wire N__88017;
    wire N__88014;
    wire N__88009;
    wire N__87998;
    wire N__87995;
    wire N__87992;
    wire N__87991;
    wire N__87988;
    wire N__87983;
    wire N__87980;
    wire N__87975;
    wire N__87972;
    wire N__87961;
    wire N__87960;
    wire N__87955;
    wire N__87954;
    wire N__87953;
    wire N__87952;
    wire N__87951;
    wire N__87950;
    wire N__87949;
    wire N__87948;
    wire N__87947;
    wire N__87946;
    wire N__87945;
    wire N__87944;
    wire N__87943;
    wire N__87942;
    wire N__87941;
    wire N__87940;
    wire N__87937;
    wire N__87904;
    wire N__87901;
    wire N__87898;
    wire N__87895;
    wire N__87892;
    wire N__87889;
    wire N__87886;
    wire N__87883;
    wire N__87882;
    wire N__87881;
    wire N__87874;
    wire N__87871;
    wire N__87868;
    wire N__87867;
    wire N__87864;
    wire N__87861;
    wire N__87856;
    wire N__87853;
    wire N__87850;
    wire N__87849;
    wire N__87846;
    wire N__87843;
    wire N__87838;
    wire N__87835;
    wire N__87832;
    wire N__87829;
    wire N__87826;
    wire N__87823;
    wire N__87822;
    wire N__87817;
    wire N__87814;
    wire N__87811;
    wire N__87808;
    wire N__87805;
    wire N__87804;
    wire N__87803;
    wire N__87802;
    wire N__87801;
    wire N__87800;
    wire N__87797;
    wire N__87794;
    wire N__87791;
    wire N__87790;
    wire N__87787;
    wire N__87784;
    wire N__87781;
    wire N__87780;
    wire N__87779;
    wire N__87778;
    wire N__87777;
    wire N__87776;
    wire N__87775;
    wire N__87774;
    wire N__87773;
    wire N__87770;
    wire N__87767;
    wire N__87764;
    wire N__87761;
    wire N__87760;
    wire N__87757;
    wire N__87752;
    wire N__87751;
    wire N__87750;
    wire N__87749;
    wire N__87746;
    wire N__87741;
    wire N__87738;
    wire N__87733;
    wire N__87730;
    wire N__87727;
    wire N__87724;
    wire N__87719;
    wire N__87716;
    wire N__87713;
    wire N__87710;
    wire N__87707;
    wire N__87704;
    wire N__87701;
    wire N__87698;
    wire N__87695;
    wire N__87692;
    wire N__87687;
    wire N__87684;
    wire N__87681;
    wire N__87676;
    wire N__87675;
    wire N__87674;
    wire N__87671;
    wire N__87668;
    wire N__87667;
    wire N__87660;
    wire N__87653;
    wire N__87648;
    wire N__87641;
    wire N__87638;
    wire N__87635;
    wire N__87630;
    wire N__87627;
    wire N__87624;
    wire N__87619;
    wire N__87616;
    wire N__87601;
    wire N__87600;
    wire N__87597;
    wire N__87594;
    wire N__87593;
    wire N__87590;
    wire N__87587;
    wire N__87586;
    wire N__87583;
    wire N__87580;
    wire N__87577;
    wire N__87574;
    wire N__87565;
    wire N__87562;
    wire N__87561;
    wire N__87560;
    wire N__87559;
    wire N__87558;
    wire N__87555;
    wire N__87554;
    wire N__87551;
    wire N__87550;
    wire N__87547;
    wire N__87544;
    wire N__87541;
    wire N__87540;
    wire N__87537;
    wire N__87534;
    wire N__87533;
    wire N__87530;
    wire N__87529;
    wire N__87526;
    wire N__87523;
    wire N__87518;
    wire N__87515;
    wire N__87512;
    wire N__87509;
    wire N__87506;
    wire N__87503;
    wire N__87500;
    wire N__87495;
    wire N__87490;
    wire N__87487;
    wire N__87480;
    wire N__87469;
    wire N__87468;
    wire N__87465;
    wire N__87462;
    wire N__87461;
    wire N__87456;
    wire N__87453;
    wire N__87448;
    wire N__87447;
    wire N__87444;
    wire N__87443;
    wire N__87440;
    wire N__87437;
    wire N__87436;
    wire N__87435;
    wire N__87434;
    wire N__87431;
    wire N__87430;
    wire N__87429;
    wire N__87428;
    wire N__87423;
    wire N__87422;
    wire N__87419;
    wire N__87418;
    wire N__87417;
    wire N__87416;
    wire N__87411;
    wire N__87410;
    wire N__87409;
    wire N__87408;
    wire N__87405;
    wire N__87404;
    wire N__87403;
    wire N__87400;
    wire N__87399;
    wire N__87396;
    wire N__87393;
    wire N__87390;
    wire N__87389;
    wire N__87388;
    wire N__87383;
    wire N__87380;
    wire N__87377;
    wire N__87376;
    wire N__87375;
    wire N__87374;
    wire N__87371;
    wire N__87368;
    wire N__87365;
    wire N__87362;
    wire N__87359;
    wire N__87358;
    wire N__87355;
    wire N__87352;
    wire N__87349;
    wire N__87348;
    wire N__87343;
    wire N__87340;
    wire N__87337;
    wire N__87334;
    wire N__87331;
    wire N__87330;
    wire N__87329;
    wire N__87326;
    wire N__87321;
    wire N__87318;
    wire N__87313;
    wire N__87308;
    wire N__87301;
    wire N__87298;
    wire N__87295;
    wire N__87292;
    wire N__87289;
    wire N__87286;
    wire N__87283;
    wire N__87280;
    wire N__87279;
    wire N__87278;
    wire N__87273;
    wire N__87272;
    wire N__87271;
    wire N__87270;
    wire N__87265;
    wire N__87262;
    wire N__87259;
    wire N__87258;
    wire N__87253;
    wire N__87242;
    wire N__87239;
    wire N__87230;
    wire N__87227;
    wire N__87224;
    wire N__87221;
    wire N__87218;
    wire N__87213;
    wire N__87210;
    wire N__87207;
    wire N__87200;
    wire N__87195;
    wire N__87188;
    wire N__87169;
    wire N__87166;
    wire N__87165;
    wire N__87160;
    wire N__87157;
    wire N__87154;
    wire N__87153;
    wire N__87148;
    wire N__87145;
    wire N__87144;
    wire N__87143;
    wire N__87142;
    wire N__87141;
    wire N__87140;
    wire N__87139;
    wire N__87138;
    wire N__87135;
    wire N__87132;
    wire N__87129;
    wire N__87128;
    wire N__87125;
    wire N__87118;
    wire N__87115;
    wire N__87114;
    wire N__87113;
    wire N__87110;
    wire N__87107;
    wire N__87106;
    wire N__87105;
    wire N__87104;
    wire N__87103;
    wire N__87102;
    wire N__87099;
    wire N__87098;
    wire N__87095;
    wire N__87094;
    wire N__87093;
    wire N__87090;
    wire N__87089;
    wire N__87088;
    wire N__87083;
    wire N__87080;
    wire N__87077;
    wire N__87074;
    wire N__87073;
    wire N__87072;
    wire N__87069;
    wire N__87064;
    wire N__87061;
    wire N__87056;
    wire N__87055;
    wire N__87052;
    wire N__87049;
    wire N__87048;
    wire N__87047;
    wire N__87044;
    wire N__87039;
    wire N__87036;
    wire N__87035;
    wire N__87034;
    wire N__87033;
    wire N__87032;
    wire N__87031;
    wire N__87030;
    wire N__87027;
    wire N__87026;
    wire N__87025;
    wire N__87022;
    wire N__87019;
    wire N__87014;
    wire N__87011;
    wire N__87006;
    wire N__87001;
    wire N__86996;
    wire N__86993;
    wire N__86992;
    wire N__86991;
    wire N__86990;
    wire N__86985;
    wire N__86982;
    wire N__86979;
    wire N__86972;
    wire N__86971;
    wire N__86970;
    wire N__86967;
    wire N__86958;
    wire N__86953;
    wire N__86948;
    wire N__86941;
    wire N__86940;
    wire N__86939;
    wire N__86938;
    wire N__86937;
    wire N__86936;
    wire N__86935;
    wire N__86934;
    wire N__86927;
    wire N__86924;
    wire N__86915;
    wire N__86912;
    wire N__86909;
    wire N__86904;
    wire N__86903;
    wire N__86902;
    wire N__86899;
    wire N__86896;
    wire N__86891;
    wire N__86888;
    wire N__86883;
    wire N__86876;
    wire N__86871;
    wire N__86868;
    wire N__86865;
    wire N__86862;
    wire N__86855;
    wire N__86850;
    wire N__86845;
    wire N__86838;
    wire N__86831;
    wire N__86812;
    wire N__86809;
    wire N__86806;
    wire N__86803;
    wire N__86800;
    wire N__86797;
    wire N__86794;
    wire N__86791;
    wire N__86788;
    wire N__86785;
    wire N__86784;
    wire N__86783;
    wire N__86782;
    wire N__86779;
    wire N__86778;
    wire N__86777;
    wire N__86776;
    wire N__86775;
    wire N__86774;
    wire N__86771;
    wire N__86768;
    wire N__86765;
    wire N__86762;
    wire N__86761;
    wire N__86760;
    wire N__86759;
    wire N__86756;
    wire N__86755;
    wire N__86752;
    wire N__86751;
    wire N__86748;
    wire N__86745;
    wire N__86744;
    wire N__86741;
    wire N__86738;
    wire N__86735;
    wire N__86732;
    wire N__86729;
    wire N__86726;
    wire N__86723;
    wire N__86720;
    wire N__86717;
    wire N__86714;
    wire N__86711;
    wire N__86708;
    wire N__86705;
    wire N__86702;
    wire N__86699;
    wire N__86694;
    wire N__86689;
    wire N__86686;
    wire N__86683;
    wire N__86680;
    wire N__86673;
    wire N__86668;
    wire N__86663;
    wire N__86658;
    wire N__86655;
    wire N__86652;
    wire N__86649;
    wire N__86644;
    wire N__86641;
    wire N__86638;
    wire N__86635;
    wire N__86630;
    wire N__86625;
    wire N__86620;
    wire N__86617;
    wire N__86614;
    wire N__86611;
    wire N__86602;
    wire N__86601;
    wire N__86600;
    wire N__86599;
    wire N__86598;
    wire N__86597;
    wire N__86596;
    wire N__86595;
    wire N__86594;
    wire N__86593;
    wire N__86592;
    wire N__86591;
    wire N__86590;
    wire N__86589;
    wire N__86588;
    wire N__86587;
    wire N__86586;
    wire N__86585;
    wire N__86584;
    wire N__86583;
    wire N__86582;
    wire N__86581;
    wire N__86580;
    wire N__86577;
    wire N__86572;
    wire N__86567;
    wire N__86562;
    wire N__86559;
    wire N__86546;
    wire N__86543;
    wire N__86540;
    wire N__86535;
    wire N__86532;
    wire N__86529;
    wire N__86526;
    wire N__86523;
    wire N__86520;
    wire N__86519;
    wire N__86518;
    wire N__86517;
    wire N__86516;
    wire N__86515;
    wire N__86514;
    wire N__86513;
    wire N__86512;
    wire N__86511;
    wire N__86510;
    wire N__86509;
    wire N__86508;
    wire N__86507;
    wire N__86506;
    wire N__86505;
    wire N__86504;
    wire N__86503;
    wire N__86502;
    wire N__86501;
    wire N__86500;
    wire N__86499;
    wire N__86498;
    wire N__86497;
    wire N__86496;
    wire N__86495;
    wire N__86494;
    wire N__86493;
    wire N__86492;
    wire N__86491;
    wire N__86490;
    wire N__86489;
    wire N__86488;
    wire N__86487;
    wire N__86486;
    wire N__86485;
    wire N__86484;
    wire N__86483;
    wire N__86482;
    wire N__86481;
    wire N__86480;
    wire N__86479;
    wire N__86478;
    wire N__86477;
    wire N__86476;
    wire N__86475;
    wire N__86474;
    wire N__86473;
    wire N__86472;
    wire N__86471;
    wire N__86470;
    wire N__86469;
    wire N__86468;
    wire N__86467;
    wire N__86466;
    wire N__86465;
    wire N__86464;
    wire N__86463;
    wire N__86462;
    wire N__86461;
    wire N__86460;
    wire N__86459;
    wire N__86458;
    wire N__86457;
    wire N__86456;
    wire N__86455;
    wire N__86454;
    wire N__86453;
    wire N__86452;
    wire N__86451;
    wire N__86450;
    wire N__86449;
    wire N__86448;
    wire N__86447;
    wire N__86446;
    wire N__86445;
    wire N__86444;
    wire N__86443;
    wire N__86442;
    wire N__86441;
    wire N__86440;
    wire N__86439;
    wire N__86438;
    wire N__86437;
    wire N__86436;
    wire N__86435;
    wire N__86434;
    wire N__86433;
    wire N__86432;
    wire N__86431;
    wire N__86430;
    wire N__86429;
    wire N__86428;
    wire N__86427;
    wire N__86426;
    wire N__86425;
    wire N__86424;
    wire N__86423;
    wire N__86422;
    wire N__86421;
    wire N__86420;
    wire N__86419;
    wire N__86418;
    wire N__86417;
    wire N__86416;
    wire N__86415;
    wire N__86414;
    wire N__86413;
    wire N__86412;
    wire N__86411;
    wire N__86410;
    wire N__86409;
    wire N__86408;
    wire N__86407;
    wire N__86406;
    wire N__86405;
    wire N__86404;
    wire N__86403;
    wire N__86402;
    wire N__86401;
    wire N__86400;
    wire N__86399;
    wire N__86398;
    wire N__86397;
    wire N__86396;
    wire N__86395;
    wire N__86394;
    wire N__86393;
    wire N__86392;
    wire N__86391;
    wire N__86390;
    wire N__86389;
    wire N__86388;
    wire N__86387;
    wire N__86386;
    wire N__86385;
    wire N__86384;
    wire N__86383;
    wire N__86382;
    wire N__86381;
    wire N__86380;
    wire N__86379;
    wire N__86378;
    wire N__86377;
    wire N__86376;
    wire N__86375;
    wire N__86374;
    wire N__86373;
    wire N__86372;
    wire N__86371;
    wire N__86370;
    wire N__86369;
    wire N__86368;
    wire N__86367;
    wire N__86366;
    wire N__86365;
    wire N__86364;
    wire N__86363;
    wire N__86362;
    wire N__86361;
    wire N__86360;
    wire N__86359;
    wire N__86358;
    wire N__86357;
    wire N__86356;
    wire N__86355;
    wire N__86354;
    wire N__86353;
    wire N__86352;
    wire N__86349;
    wire N__86346;
    wire N__86343;
    wire N__86340;
    wire N__86337;
    wire N__86334;
    wire N__86331;
    wire N__86328;
    wire N__86325;
    wire N__86322;
    wire N__86319;
    wire N__86316;
    wire N__86313;
    wire N__86310;
    wire N__85945;
    wire N__85942;
    wire N__85939;
    wire N__85938;
    wire N__85937;
    wire N__85936;
    wire N__85935;
    wire N__85934;
    wire N__85931;
    wire N__85930;
    wire N__85929;
    wire N__85928;
    wire N__85927;
    wire N__85926;
    wire N__85925;
    wire N__85924;
    wire N__85923;
    wire N__85920;
    wire N__85919;
    wire N__85916;
    wire N__85913;
    wire N__85912;
    wire N__85911;
    wire N__85910;
    wire N__85909;
    wire N__85904;
    wire N__85901;
    wire N__85892;
    wire N__85889;
    wire N__85886;
    wire N__85883;
    wire N__85880;
    wire N__85877;
    wire N__85874;
    wire N__85871;
    wire N__85868;
    wire N__85861;
    wire N__85860;
    wire N__85857;
    wire N__85850;
    wire N__85849;
    wire N__85846;
    wire N__85843;
    wire N__85842;
    wire N__85841;
    wire N__85832;
    wire N__85825;
    wire N__85822;
    wire N__85817;
    wire N__85814;
    wire N__85809;
    wire N__85804;
    wire N__85799;
    wire N__85794;
    wire N__85783;
    wire N__85780;
    wire N__85777;
    wire N__85776;
    wire N__85775;
    wire N__85772;
    wire N__85771;
    wire N__85770;
    wire N__85769;
    wire N__85768;
    wire N__85765;
    wire N__85764;
    wire N__85763;
    wire N__85760;
    wire N__85757;
    wire N__85754;
    wire N__85751;
    wire N__85750;
    wire N__85749;
    wire N__85748;
    wire N__85747;
    wire N__85746;
    wire N__85743;
    wire N__85740;
    wire N__85739;
    wire N__85738;
    wire N__85737;
    wire N__85734;
    wire N__85733;
    wire N__85728;
    wire N__85725;
    wire N__85720;
    wire N__85717;
    wire N__85716;
    wire N__85713;
    wire N__85710;
    wire N__85707;
    wire N__85704;
    wire N__85701;
    wire N__85698;
    wire N__85695;
    wire N__85692;
    wire N__85687;
    wire N__85684;
    wire N__85681;
    wire N__85678;
    wire N__85675;
    wire N__85670;
    wire N__85667;
    wire N__85662;
    wire N__85655;
    wire N__85648;
    wire N__85645;
    wire N__85640;
    wire N__85633;
    wire N__85628;
    wire N__85625;
    wire N__85620;
    wire N__85617;
    wire N__85614;
    wire N__85609;
    wire N__85600;
    wire N__85599;
    wire N__85596;
    wire N__85593;
    wire N__85592;
    wire N__85589;
    wire N__85586;
    wire N__85583;
    wire N__85580;
    wire N__85573;
    wire N__85570;
    wire N__85567;
    wire N__85566;
    wire N__85563;
    wire N__85560;
    wire N__85557;
    wire N__85554;
    wire N__85549;
    wire N__85546;
    wire N__85543;
    wire N__85540;
    wire N__85537;
    wire N__85534;
    wire N__85531;
    wire N__85530;
    wire N__85529;
    wire N__85528;
    wire N__85527;
    wire N__85526;
    wire N__85523;
    wire N__85520;
    wire N__85517;
    wire N__85514;
    wire N__85513;
    wire N__85510;
    wire N__85509;
    wire N__85506;
    wire N__85499;
    wire N__85496;
    wire N__85493;
    wire N__85490;
    wire N__85489;
    wire N__85486;
    wire N__85485;
    wire N__85482;
    wire N__85481;
    wire N__85480;
    wire N__85477;
    wire N__85472;
    wire N__85469;
    wire N__85468;
    wire N__85465;
    wire N__85464;
    wire N__85461;
    wire N__85458;
    wire N__85457;
    wire N__85454;
    wire N__85449;
    wire N__85446;
    wire N__85445;
    wire N__85442;
    wire N__85439;
    wire N__85436;
    wire N__85433;
    wire N__85430;
    wire N__85427;
    wire N__85424;
    wire N__85421;
    wire N__85418;
    wire N__85415;
    wire N__85414;
    wire N__85411;
    wire N__85408;
    wire N__85403;
    wire N__85396;
    wire N__85389;
    wire N__85384;
    wire N__85381;
    wire N__85366;
    wire N__85363;
    wire N__85360;
    wire N__85357;
    wire N__85354;
    wire N__85351;
    wire N__85348;
    wire N__85345;
    wire N__85342;
    wire N__85339;
    wire N__85336;
    wire N__85333;
    wire N__85330;
    wire N__85327;
    wire N__85324;
    wire N__85321;
    wire N__85318;
    wire N__85315;
    wire N__85312;
    wire N__85309;
    wire N__85306;
    wire N__85303;
    wire N__85300;
    wire N__85297;
    wire N__85294;
    wire N__85291;
    wire N__85288;
    wire N__85285;
    wire N__85282;
    wire N__85279;
    wire N__85276;
    wire N__85275;
    wire N__85270;
    wire N__85267;
    wire N__85264;
    wire N__85261;
    wire N__85258;
    wire N__85255;
    wire N__85252;
    wire N__85251;
    wire N__85250;
    wire N__85247;
    wire N__85246;
    wire N__85243;
    wire N__85240;
    wire N__85237;
    wire N__85234;
    wire N__85233;
    wire N__85232;
    wire N__85229;
    wire N__85226;
    wire N__85225;
    wire N__85222;
    wire N__85217;
    wire N__85214;
    wire N__85211;
    wire N__85208;
    wire N__85205;
    wire N__85200;
    wire N__85195;
    wire N__85190;
    wire N__85187;
    wire N__85180;
    wire N__85179;
    wire N__85178;
    wire N__85175;
    wire N__85172;
    wire N__85169;
    wire N__85166;
    wire N__85165;
    wire N__85162;
    wire N__85161;
    wire N__85160;
    wire N__85159;
    wire N__85158;
    wire N__85157;
    wire N__85156;
    wire N__85153;
    wire N__85150;
    wire N__85147;
    wire N__85144;
    wire N__85141;
    wire N__85138;
    wire N__85137;
    wire N__85134;
    wire N__85133;
    wire N__85132;
    wire N__85129;
    wire N__85128;
    wire N__85127;
    wire N__85124;
    wire N__85121;
    wire N__85118;
    wire N__85117;
    wire N__85116;
    wire N__85115;
    wire N__85114;
    wire N__85111;
    wire N__85104;
    wire N__85101;
    wire N__85096;
    wire N__85091;
    wire N__85088;
    wire N__85085;
    wire N__85084;
    wire N__85081;
    wire N__85078;
    wire N__85077;
    wire N__85076;
    wire N__85073;
    wire N__85070;
    wire N__85069;
    wire N__85068;
    wire N__85067;
    wire N__85066;
    wire N__85065;
    wire N__85062;
    wire N__85055;
    wire N__85054;
    wire N__85045;
    wire N__85038;
    wire N__85035;
    wire N__85034;
    wire N__85029;
    wire N__85026;
    wire N__85025;
    wire N__85022;
    wire N__85019;
    wire N__85016;
    wire N__85013;
    wire N__85006;
    wire N__85005;
    wire N__85002;
    wire N__84997;
    wire N__84994;
    wire N__84989;
    wire N__84986;
    wire N__84983;
    wire N__84980;
    wire N__84973;
    wire N__84964;
    wire N__84959;
    wire N__84954;
    wire N__84951;
    wire N__84934;
    wire N__84933;
    wire N__84932;
    wire N__84929;
    wire N__84926;
    wire N__84923;
    wire N__84922;
    wire N__84919;
    wire N__84916;
    wire N__84915;
    wire N__84912;
    wire N__84911;
    wire N__84908;
    wire N__84905;
    wire N__84902;
    wire N__84899;
    wire N__84898;
    wire N__84897;
    wire N__84896;
    wire N__84893;
    wire N__84890;
    wire N__84887;
    wire N__84884;
    wire N__84879;
    wire N__84872;
    wire N__84867;
    wire N__84864;
    wire N__84853;
    wire N__84850;
    wire N__84847;
    wire N__84844;
    wire N__84841;
    wire N__84838;
    wire N__84837;
    wire N__84836;
    wire N__84835;
    wire N__84834;
    wire N__84833;
    wire N__84832;
    wire N__84831;
    wire N__84828;
    wire N__84827;
    wire N__84826;
    wire N__84823;
    wire N__84820;
    wire N__84817;
    wire N__84816;
    wire N__84815;
    wire N__84812;
    wire N__84809;
    wire N__84806;
    wire N__84803;
    wire N__84800;
    wire N__84797;
    wire N__84794;
    wire N__84791;
    wire N__84788;
    wire N__84787;
    wire N__84786;
    wire N__84785;
    wire N__84782;
    wire N__84777;
    wire N__84774;
    wire N__84771;
    wire N__84770;
    wire N__84769;
    wire N__84768;
    wire N__84765;
    wire N__84762;
    wire N__84761;
    wire N__84758;
    wire N__84753;
    wire N__84748;
    wire N__84745;
    wire N__84740;
    wire N__84735;
    wire N__84732;
    wire N__84729;
    wire N__84722;
    wire N__84719;
    wire N__84716;
    wire N__84713;
    wire N__84706;
    wire N__84699;
    wire N__84682;
    wire N__84679;
    wire N__84678;
    wire N__84675;
    wire N__84672;
    wire N__84671;
    wire N__84668;
    wire N__84663;
    wire N__84662;
    wire N__84661;
    wire N__84660;
    wire N__84659;
    wire N__84656;
    wire N__84653;
    wire N__84650;
    wire N__84647;
    wire N__84644;
    wire N__84641;
    wire N__84638;
    wire N__84635;
    wire N__84632;
    wire N__84629;
    wire N__84628;
    wire N__84623;
    wire N__84616;
    wire N__84613;
    wire N__84610;
    wire N__84607;
    wire N__84602;
    wire N__84595;
    wire N__84592;
    wire N__84589;
    wire N__84586;
    wire N__84583;
    wire N__84580;
    wire N__84577;
    wire N__84576;
    wire N__84575;
    wire N__84572;
    wire N__84565;
    wire N__84564;
    wire N__84563;
    wire N__84562;
    wire N__84561;
    wire N__84560;
    wire N__84557;
    wire N__84554;
    wire N__84551;
    wire N__84550;
    wire N__84549;
    wire N__84548;
    wire N__84547;
    wire N__84546;
    wire N__84545;
    wire N__84544;
    wire N__84543;
    wire N__84542;
    wire N__84541;
    wire N__84540;
    wire N__84539;
    wire N__84538;
    wire N__84537;
    wire N__84530;
    wire N__84523;
    wire N__84522;
    wire N__84521;
    wire N__84518;
    wire N__84517;
    wire N__84516;
    wire N__84515;
    wire N__84510;
    wire N__84509;
    wire N__84508;
    wire N__84505;
    wire N__84504;
    wire N__84501;
    wire N__84500;
    wire N__84493;
    wire N__84492;
    wire N__84491;
    wire N__84488;
    wire N__84487;
    wire N__84486;
    wire N__84483;
    wire N__84478;
    wire N__84477;
    wire N__84476;
    wire N__84475;
    wire N__84474;
    wire N__84473;
    wire N__84470;
    wire N__84469;
    wire N__84468;
    wire N__84465;
    wire N__84460;
    wire N__84457;
    wire N__84454;
    wire N__84451;
    wire N__84444;
    wire N__84441;
    wire N__84436;
    wire N__84435;
    wire N__84434;
    wire N__84433;
    wire N__84432;
    wire N__84429;
    wire N__84426;
    wire N__84423;
    wire N__84420;
    wire N__84419;
    wire N__84416;
    wire N__84415;
    wire N__84414;
    wire N__84413;
    wire N__84408;
    wire N__84405;
    wire N__84404;
    wire N__84403;
    wire N__84402;
    wire N__84401;
    wire N__84398;
    wire N__84395;
    wire N__84390;
    wire N__84385;
    wire N__84378;
    wire N__84375;
    wire N__84370;
    wire N__84367;
    wire N__84362;
    wire N__84355;
    wire N__84350;
    wire N__84345;
    wire N__84342;
    wire N__84339;
    wire N__84330;
    wire N__84327;
    wire N__84324;
    wire N__84323;
    wire N__84322;
    wire N__84321;
    wire N__84316;
    wire N__84313;
    wire N__84308;
    wire N__84303;
    wire N__84298;
    wire N__84287;
    wire N__84284;
    wire N__84281;
    wire N__84278;
    wire N__84267;
    wire N__84260;
    wire N__84257;
    wire N__84256;
    wire N__84255;
    wire N__84252;
    wire N__84249;
    wire N__84246;
    wire N__84233;
    wire N__84224;
    wire N__84219;
    wire N__84214;
    wire N__84199;
    wire N__84196;
    wire N__84193;
    wire N__84192;
    wire N__84189;
    wire N__84188;
    wire N__84187;
    wire N__84186;
    wire N__84183;
    wire N__84182;
    wire N__84181;
    wire N__84180;
    wire N__84179;
    wire N__84178;
    wire N__84175;
    wire N__84172;
    wire N__84169;
    wire N__84168;
    wire N__84165;
    wire N__84162;
    wire N__84159;
    wire N__84158;
    wire N__84155;
    wire N__84150;
    wire N__84147;
    wire N__84144;
    wire N__84141;
    wire N__84138;
    wire N__84135;
    wire N__84134;
    wire N__84133;
    wire N__84132;
    wire N__84129;
    wire N__84126;
    wire N__84123;
    wire N__84120;
    wire N__84119;
    wire N__84118;
    wire N__84117;
    wire N__84116;
    wire N__84113;
    wire N__84108;
    wire N__84101;
    wire N__84100;
    wire N__84097;
    wire N__84094;
    wire N__84093;
    wire N__84092;
    wire N__84091;
    wire N__84088;
    wire N__84087;
    wire N__84084;
    wire N__84083;
    wire N__84082;
    wire N__84081;
    wire N__84078;
    wire N__84073;
    wire N__84070;
    wire N__84067;
    wire N__84064;
    wire N__84063;
    wire N__84060;
    wire N__84057;
    wire N__84056;
    wire N__84053;
    wire N__84048;
    wire N__84045;
    wire N__84042;
    wire N__84039;
    wire N__84036;
    wire N__84031;
    wire N__84028;
    wire N__84027;
    wire N__84024;
    wire N__84019;
    wire N__84014;
    wire N__84011;
    wire N__84008;
    wire N__84003;
    wire N__83996;
    wire N__83993;
    wire N__83990;
    wire N__83983;
    wire N__83978;
    wire N__83973;
    wire N__83970;
    wire N__83967;
    wire N__83964;
    wire N__83959;
    wire N__83952;
    wire N__83949;
    wire N__83938;
    wire N__83935;
    wire N__83932;
    wire N__83927;
    wire N__83924;
    wire N__83921;
    wire N__83918;
    wire N__83905;
    wire N__83902;
    wire N__83901;
    wire N__83900;
    wire N__83899;
    wire N__83898;
    wire N__83895;
    wire N__83894;
    wire N__83891;
    wire N__83890;
    wire N__83889;
    wire N__83888;
    wire N__83885;
    wire N__83882;
    wire N__83879;
    wire N__83878;
    wire N__83877;
    wire N__83874;
    wire N__83871;
    wire N__83868;
    wire N__83865;
    wire N__83862;
    wire N__83859;
    wire N__83856;
    wire N__83851;
    wire N__83848;
    wire N__83845;
    wire N__83840;
    wire N__83837;
    wire N__83834;
    wire N__83831;
    wire N__83824;
    wire N__83821;
    wire N__83818;
    wire N__83815;
    wire N__83812;
    wire N__83809;
    wire N__83806;
    wire N__83803;
    wire N__83798;
    wire N__83795;
    wire N__83792;
    wire N__83787;
    wire N__83784;
    wire N__83781;
    wire N__83778;
    wire N__83775;
    wire N__83772;
    wire N__83769;
    wire N__83766;
    wire N__83763;
    wire N__83752;
    wire N__83749;
    wire N__83746;
    wire N__83743;
    wire N__83740;
    wire N__83737;
    wire N__83734;
    wire N__83731;
    wire N__83728;
    wire N__83725;
    wire N__83724;
    wire N__83723;
    wire N__83722;
    wire N__83721;
    wire N__83716;
    wire N__83709;
    wire N__83704;
    wire N__83701;
    wire N__83698;
    wire N__83695;
    wire N__83692;
    wire N__83689;
    wire N__83686;
    wire N__83683;
    wire N__83680;
    wire N__83677;
    wire N__83676;
    wire N__83675;
    wire N__83672;
    wire N__83669;
    wire N__83666;
    wire N__83663;
    wire N__83660;
    wire N__83659;
    wire N__83656;
    wire N__83651;
    wire N__83648;
    wire N__83641;
    wire N__83640;
    wire N__83639;
    wire N__83638;
    wire N__83637;
    wire N__83636;
    wire N__83635;
    wire N__83632;
    wire N__83629;
    wire N__83628;
    wire N__83625;
    wire N__83620;
    wire N__83617;
    wire N__83614;
    wire N__83611;
    wire N__83608;
    wire N__83605;
    wire N__83600;
    wire N__83597;
    wire N__83592;
    wire N__83589;
    wire N__83588;
    wire N__83585;
    wire N__83582;
    wire N__83577;
    wire N__83574;
    wire N__83571;
    wire N__83560;
    wire N__83557;
    wire N__83554;
    wire N__83551;
    wire N__83550;
    wire N__83545;
    wire N__83542;
    wire N__83539;
    wire N__83538;
    wire N__83535;
    wire N__83532;
    wire N__83527;
    wire N__83524;
    wire N__83523;
    wire N__83522;
    wire N__83519;
    wire N__83516;
    wire N__83515;
    wire N__83514;
    wire N__83511;
    wire N__83510;
    wire N__83507;
    wire N__83506;
    wire N__83497;
    wire N__83496;
    wire N__83493;
    wire N__83492;
    wire N__83491;
    wire N__83488;
    wire N__83485;
    wire N__83482;
    wire N__83481;
    wire N__83478;
    wire N__83477;
    wire N__83476;
    wire N__83475;
    wire N__83470;
    wire N__83467;
    wire N__83462;
    wire N__83459;
    wire N__83456;
    wire N__83453;
    wire N__83450;
    wire N__83447;
    wire N__83444;
    wire N__83441;
    wire N__83438;
    wire N__83435;
    wire N__83430;
    wire N__83427;
    wire N__83422;
    wire N__83419;
    wire N__83412;
    wire N__83409;
    wire N__83406;
    wire N__83403;
    wire N__83400;
    wire N__83389;
    wire N__83386;
    wire N__83383;
    wire N__83380;
    wire N__83379;
    wire N__83378;
    wire N__83377;
    wire N__83376;
    wire N__83375;
    wire N__83374;
    wire N__83371;
    wire N__83370;
    wire N__83369;
    wire N__83368;
    wire N__83367;
    wire N__83366;
    wire N__83365;
    wire N__83362;
    wire N__83359;
    wire N__83356;
    wire N__83355;
    wire N__83354;
    wire N__83351;
    wire N__83350;
    wire N__83347;
    wire N__83344;
    wire N__83341;
    wire N__83334;
    wire N__83331;
    wire N__83328;
    wire N__83325;
    wire N__83320;
    wire N__83319;
    wire N__83318;
    wire N__83315;
    wire N__83312;
    wire N__83311;
    wire N__83308;
    wire N__83305;
    wire N__83302;
    wire N__83297;
    wire N__83292;
    wire N__83289;
    wire N__83286;
    wire N__83283;
    wire N__83280;
    wire N__83275;
    wire N__83272;
    wire N__83269;
    wire N__83268;
    wire N__83267;
    wire N__83264;
    wire N__83261;
    wire N__83252;
    wire N__83249;
    wire N__83246;
    wire N__83239;
    wire N__83236;
    wire N__83233;
    wire N__83226;
    wire N__83221;
    wire N__83214;
    wire N__83203;
    wire N__83200;
    wire N__83197;
    wire N__83194;
    wire N__83191;
    wire N__83188;
    wire N__83185;
    wire N__83184;
    wire N__83183;
    wire N__83182;
    wire N__83179;
    wire N__83178;
    wire N__83177;
    wire N__83176;
    wire N__83175;
    wire N__83174;
    wire N__83171;
    wire N__83170;
    wire N__83169;
    wire N__83168;
    wire N__83167;
    wire N__83166;
    wire N__83163;
    wire N__83160;
    wire N__83157;
    wire N__83154;
    wire N__83151;
    wire N__83150;
    wire N__83147;
    wire N__83146;
    wire N__83143;
    wire N__83140;
    wire N__83133;
    wire N__83132;
    wire N__83125;
    wire N__83122;
    wire N__83119;
    wire N__83114;
    wire N__83111;
    wire N__83108;
    wire N__83105;
    wire N__83102;
    wire N__83099;
    wire N__83094;
    wire N__83091;
    wire N__83086;
    wire N__83085;
    wire N__83084;
    wire N__83083;
    wire N__83080;
    wire N__83077;
    wire N__83072;
    wire N__83069;
    wire N__83062;
    wire N__83059;
    wire N__83056;
    wire N__83049;
    wire N__83038;
    wire N__83029;
    wire N__83028;
    wire N__83027;
    wire N__83026;
    wire N__83023;
    wire N__83020;
    wire N__83019;
    wire N__83016;
    wire N__83013;
    wire N__83012;
    wire N__83011;
    wire N__83010;
    wire N__83009;
    wire N__83008;
    wire N__83003;
    wire N__83002;
    wire N__83001;
    wire N__83000;
    wire N__82999;
    wire N__82998;
    wire N__82997;
    wire N__82996;
    wire N__82993;
    wire N__82988;
    wire N__82985;
    wire N__82982;
    wire N__82979;
    wire N__82976;
    wire N__82973;
    wire N__82970;
    wire N__82967;
    wire N__82960;
    wire N__82957;
    wire N__82954;
    wire N__82951;
    wire N__82946;
    wire N__82945;
    wire N__82944;
    wire N__82943;
    wire N__82940;
    wire N__82933;
    wire N__82930;
    wire N__82925;
    wire N__82920;
    wire N__82915;
    wire N__82912;
    wire N__82905;
    wire N__82894;
    wire N__82885;
    wire N__82882;
    wire N__82879;
    wire N__82878;
    wire N__82875;
    wire N__82872;
    wire N__82867;
    wire N__82864;
    wire N__82861;
    wire N__82860;
    wire N__82859;
    wire N__82856;
    wire N__82853;
    wire N__82852;
    wire N__82851;
    wire N__82850;
    wire N__82847;
    wire N__82844;
    wire N__82841;
    wire N__82838;
    wire N__82835;
    wire N__82832;
    wire N__82829;
    wire N__82828;
    wire N__82827;
    wire N__82824;
    wire N__82821;
    wire N__82820;
    wire N__82815;
    wire N__82812;
    wire N__82809;
    wire N__82804;
    wire N__82803;
    wire N__82798;
    wire N__82795;
    wire N__82786;
    wire N__82783;
    wire N__82774;
    wire N__82773;
    wire N__82768;
    wire N__82765;
    wire N__82764;
    wire N__82763;
    wire N__82760;
    wire N__82759;
    wire N__82758;
    wire N__82757;
    wire N__82756;
    wire N__82753;
    wire N__82752;
    wire N__82751;
    wire N__82748;
    wire N__82745;
    wire N__82744;
    wire N__82743;
    wire N__82742;
    wire N__82741;
    wire N__82740;
    wire N__82739;
    wire N__82738;
    wire N__82737;
    wire N__82734;
    wire N__82731;
    wire N__82728;
    wire N__82725;
    wire N__82722;
    wire N__82719;
    wire N__82716;
    wire N__82713;
    wire N__82710;
    wire N__82707;
    wire N__82702;
    wire N__82697;
    wire N__82690;
    wire N__82689;
    wire N__82688;
    wire N__82687;
    wire N__82686;
    wire N__82685;
    wire N__82682;
    wire N__82679;
    wire N__82676;
    wire N__82671;
    wire N__82664;
    wire N__82653;
    wire N__82650;
    wire N__82647;
    wire N__82644;
    wire N__82641;
    wire N__82640;
    wire N__82639;
    wire N__82638;
    wire N__82637;
    wire N__82636;
    wire N__82635;
    wire N__82632;
    wire N__82627;
    wire N__82620;
    wire N__82615;
    wire N__82608;
    wire N__82605;
    wire N__82602;
    wire N__82597;
    wire N__82594;
    wire N__82591;
    wire N__82586;
    wire N__82583;
    wire N__82580;
    wire N__82577;
    wire N__82558;
    wire N__82555;
    wire N__82552;
    wire N__82549;
    wire N__82546;
    wire N__82545;
    wire N__82540;
    wire N__82537;
    wire N__82534;
    wire N__82533;
    wire N__82532;
    wire N__82531;
    wire N__82528;
    wire N__82523;
    wire N__82520;
    wire N__82517;
    wire N__82514;
    wire N__82511;
    wire N__82508;
    wire N__82503;
    wire N__82498;
    wire N__82497;
    wire N__82494;
    wire N__82491;
    wire N__82490;
    wire N__82487;
    wire N__82484;
    wire N__82481;
    wire N__82480;
    wire N__82479;
    wire N__82478;
    wire N__82473;
    wire N__82470;
    wire N__82463;
    wire N__82456;
    wire N__82453;
    wire N__82450;
    wire N__82447;
    wire N__82444;
    wire N__82441;
    wire N__82440;
    wire N__82435;
    wire N__82432;
    wire N__82429;
    wire N__82426;
    wire N__82423;
    wire N__82420;
    wire N__82419;
    wire N__82414;
    wire N__82411;
    wire N__82408;
    wire N__82405;
    wire N__82404;
    wire N__82403;
    wire N__82402;
    wire N__82397;
    wire N__82392;
    wire N__82387;
    wire N__82384;
    wire N__82381;
    wire N__82378;
    wire N__82375;
    wire N__82372;
    wire N__82371;
    wire N__82370;
    wire N__82369;
    wire N__82368;
    wire N__82365;
    wire N__82362;
    wire N__82355;
    wire N__82352;
    wire N__82345;
    wire N__82342;
    wire N__82341;
    wire N__82336;
    wire N__82333;
    wire N__82330;
    wire N__82327;
    wire N__82324;
    wire N__82321;
    wire N__82318;
    wire N__82317;
    wire N__82314;
    wire N__82311;
    wire N__82308;
    wire N__82305;
    wire N__82302;
    wire N__82297;
    wire N__82296;
    wire N__82293;
    wire N__82290;
    wire N__82285;
    wire N__82282;
    wire N__82279;
    wire N__82278;
    wire N__82277;
    wire N__82276;
    wire N__82271;
    wire N__82266;
    wire N__82265;
    wire N__82260;
    wire N__82259;
    wire N__82258;
    wire N__82257;
    wire N__82256;
    wire N__82255;
    wire N__82254;
    wire N__82253;
    wire N__82252;
    wire N__82249;
    wire N__82246;
    wire N__82241;
    wire N__82240;
    wire N__82237;
    wire N__82230;
    wire N__82227;
    wire N__82224;
    wire N__82217;
    wire N__82216;
    wire N__82213;
    wire N__82212;
    wire N__82211;
    wire N__82208;
    wire N__82205;
    wire N__82202;
    wire N__82197;
    wire N__82194;
    wire N__82191;
    wire N__82188;
    wire N__82187;
    wire N__82186;
    wire N__82183;
    wire N__82180;
    wire N__82177;
    wire N__82170;
    wire N__82165;
    wire N__82160;
    wire N__82147;
    wire N__82144;
    wire N__82141;
    wire N__82138;
    wire N__82135;
    wire N__82132;
    wire N__82131;
    wire N__82130;
    wire N__82129;
    wire N__82126;
    wire N__82123;
    wire N__82120;
    wire N__82117;
    wire N__82112;
    wire N__82109;
    wire N__82106;
    wire N__82103;
    wire N__82098;
    wire N__82095;
    wire N__82092;
    wire N__82087;
    wire N__82086;
    wire N__82083;
    wire N__82082;
    wire N__82079;
    wire N__82078;
    wire N__82077;
    wire N__82074;
    wire N__82071;
    wire N__82068;
    wire N__82065;
    wire N__82064;
    wire N__82061;
    wire N__82058;
    wire N__82055;
    wire N__82052;
    wire N__82051;
    wire N__82048;
    wire N__82045;
    wire N__82042;
    wire N__82037;
    wire N__82034;
    wire N__82031;
    wire N__82028;
    wire N__82025;
    wire N__82022;
    wire N__82017;
    wire N__82014;
    wire N__82011;
    wire N__82004;
    wire N__81997;
    wire N__81994;
    wire N__81991;
    wire N__81990;
    wire N__81987;
    wire N__81984;
    wire N__81981;
    wire N__81978;
    wire N__81975;
    wire N__81970;
    wire N__81967;
    wire N__81964;
    wire N__81961;
    wire N__81958;
    wire N__81957;
    wire N__81956;
    wire N__81953;
    wire N__81948;
    wire N__81945;
    wire N__81942;
    wire N__81937;
    wire N__81934;
    wire N__81931;
    wire N__81928;
    wire N__81925;
    wire N__81924;
    wire N__81923;
    wire N__81916;
    wire N__81913;
    wire N__81910;
    wire N__81907;
    wire N__81904;
    wire N__81901;
    wire N__81898;
    wire N__81897;
    wire N__81896;
    wire N__81895;
    wire N__81894;
    wire N__81891;
    wire N__81890;
    wire N__81885;
    wire N__81876;
    wire N__81873;
    wire N__81870;
    wire N__81867;
    wire N__81864;
    wire N__81859;
    wire N__81856;
    wire N__81853;
    wire N__81852;
    wire N__81849;
    wire N__81846;
    wire N__81841;
    wire N__81838;
    wire N__81835;
    wire N__81834;
    wire N__81833;
    wire N__81828;
    wire N__81827;
    wire N__81826;
    wire N__81825;
    wire N__81824;
    wire N__81823;
    wire N__81820;
    wire N__81819;
    wire N__81816;
    wire N__81811;
    wire N__81804;
    wire N__81801;
    wire N__81798;
    wire N__81793;
    wire N__81790;
    wire N__81787;
    wire N__81784;
    wire N__81779;
    wire N__81776;
    wire N__81771;
    wire N__81766;
    wire N__81763;
    wire N__81760;
    wire N__81757;
    wire N__81754;
    wire N__81751;
    wire N__81748;
    wire N__81745;
    wire N__81744;
    wire N__81743;
    wire N__81742;
    wire N__81739;
    wire N__81732;
    wire N__81727;
    wire N__81726;
    wire N__81725;
    wire N__81722;
    wire N__81719;
    wire N__81716;
    wire N__81713;
    wire N__81708;
    wire N__81703;
    wire N__81700;
    wire N__81697;
    wire N__81694;
    wire N__81691;
    wire N__81688;
    wire N__81685;
    wire N__81684;
    wire N__81683;
    wire N__81682;
    wire N__81679;
    wire N__81674;
    wire N__81671;
    wire N__81666;
    wire N__81663;
    wire N__81660;
    wire N__81655;
    wire N__81654;
    wire N__81653;
    wire N__81650;
    wire N__81649;
    wire N__81648;
    wire N__81647;
    wire N__81644;
    wire N__81641;
    wire N__81640;
    wire N__81637;
    wire N__81634;
    wire N__81631;
    wire N__81630;
    wire N__81627;
    wire N__81624;
    wire N__81621;
    wire N__81618;
    wire N__81615;
    wire N__81612;
    wire N__81609;
    wire N__81606;
    wire N__81603;
    wire N__81602;
    wire N__81599;
    wire N__81594;
    wire N__81589;
    wire N__81584;
    wire N__81581;
    wire N__81578;
    wire N__81577;
    wire N__81576;
    wire N__81575;
    wire N__81574;
    wire N__81569;
    wire N__81564;
    wire N__81561;
    wire N__81556;
    wire N__81553;
    wire N__81548;
    wire N__81535;
    wire N__81534;
    wire N__81533;
    wire N__81530;
    wire N__81527;
    wire N__81526;
    wire N__81525;
    wire N__81524;
    wire N__81521;
    wire N__81520;
    wire N__81517;
    wire N__81514;
    wire N__81511;
    wire N__81506;
    wire N__81503;
    wire N__81500;
    wire N__81499;
    wire N__81496;
    wire N__81493;
    wire N__81488;
    wire N__81487;
    wire N__81484;
    wire N__81481;
    wire N__81478;
    wire N__81475;
    wire N__81472;
    wire N__81469;
    wire N__81466;
    wire N__81459;
    wire N__81448;
    wire N__81445;
    wire N__81444;
    wire N__81443;
    wire N__81442;
    wire N__81441;
    wire N__81438;
    wire N__81435;
    wire N__81432;
    wire N__81429;
    wire N__81426;
    wire N__81425;
    wire N__81420;
    wire N__81419;
    wire N__81416;
    wire N__81411;
    wire N__81408;
    wire N__81405;
    wire N__81404;
    wire N__81403;
    wire N__81400;
    wire N__81395;
    wire N__81390;
    wire N__81387;
    wire N__81384;
    wire N__81373;
    wire N__81370;
    wire N__81367;
    wire N__81364;
    wire N__81361;
    wire N__81358;
    wire N__81355;
    wire N__81352;
    wire N__81349;
    wire N__81346;
    wire N__81343;
    wire N__81340;
    wire N__81337;
    wire N__81334;
    wire N__81333;
    wire N__81332;
    wire N__81329;
    wire N__81328;
    wire N__81327;
    wire N__81326;
    wire N__81325;
    wire N__81324;
    wire N__81323;
    wire N__81322;
    wire N__81319;
    wire N__81318;
    wire N__81315;
    wire N__81314;
    wire N__81313;
    wire N__81312;
    wire N__81311;
    wire N__81310;
    wire N__81309;
    wire N__81306;
    wire N__81301;
    wire N__81298;
    wire N__81293;
    wire N__81292;
    wire N__81287;
    wire N__81286;
    wire N__81283;
    wire N__81280;
    wire N__81277;
    wire N__81274;
    wire N__81269;
    wire N__81264;
    wire N__81261;
    wire N__81260;
    wire N__81259;
    wire N__81256;
    wire N__81253;
    wire N__81248;
    wire N__81245;
    wire N__81244;
    wire N__81243;
    wire N__81240;
    wire N__81237;
    wire N__81228;
    wire N__81221;
    wire N__81218;
    wire N__81215;
    wire N__81212;
    wire N__81205;
    wire N__81202;
    wire N__81201;
    wire N__81198;
    wire N__81195;
    wire N__81188;
    wire N__81187;
    wire N__81184;
    wire N__81175;
    wire N__81172;
    wire N__81165;
    wire N__81162;
    wire N__81157;
    wire N__81152;
    wire N__81145;
    wire N__81142;
    wire N__81139;
    wire N__81136;
    wire N__81133;
    wire N__81130;
    wire N__81127;
    wire N__81126;
    wire N__81123;
    wire N__81120;
    wire N__81117;
    wire N__81112;
    wire N__81111;
    wire N__81110;
    wire N__81107;
    wire N__81104;
    wire N__81103;
    wire N__81100;
    wire N__81099;
    wire N__81098;
    wire N__81097;
    wire N__81094;
    wire N__81091;
    wire N__81088;
    wire N__81085;
    wire N__81082;
    wire N__81081;
    wire N__81076;
    wire N__81073;
    wire N__81068;
    wire N__81067;
    wire N__81064;
    wire N__81061;
    wire N__81058;
    wire N__81055;
    wire N__81050;
    wire N__81047;
    wire N__81044;
    wire N__81041;
    wire N__81038;
    wire N__81025;
    wire N__81024;
    wire N__81023;
    wire N__81022;
    wire N__81019;
    wire N__81014;
    wire N__81013;
    wire N__81010;
    wire N__81009;
    wire N__81006;
    wire N__81003;
    wire N__81000;
    wire N__80997;
    wire N__80994;
    wire N__80991;
    wire N__80986;
    wire N__80983;
    wire N__80980;
    wire N__80979;
    wire N__80978;
    wire N__80977;
    wire N__80972;
    wire N__80967;
    wire N__80962;
    wire N__80959;
    wire N__80950;
    wire N__80949;
    wire N__80948;
    wire N__80947;
    wire N__80944;
    wire N__80941;
    wire N__80940;
    wire N__80937;
    wire N__80936;
    wire N__80935;
    wire N__80934;
    wire N__80931;
    wire N__80928;
    wire N__80923;
    wire N__80920;
    wire N__80915;
    wire N__80912;
    wire N__80909;
    wire N__80906;
    wire N__80903;
    wire N__80898;
    wire N__80895;
    wire N__80892;
    wire N__80889;
    wire N__80886;
    wire N__80883;
    wire N__80878;
    wire N__80869;
    wire N__80868;
    wire N__80867;
    wire N__80866;
    wire N__80865;
    wire N__80864;
    wire N__80863;
    wire N__80860;
    wire N__80857;
    wire N__80854;
    wire N__80853;
    wire N__80850;
    wire N__80845;
    wire N__80842;
    wire N__80839;
    wire N__80836;
    wire N__80833;
    wire N__80832;
    wire N__80829;
    wire N__80822;
    wire N__80817;
    wire N__80816;
    wire N__80813;
    wire N__80810;
    wire N__80807;
    wire N__80802;
    wire N__80799;
    wire N__80788;
    wire N__80785;
    wire N__80782;
    wire N__80779;
    wire N__80776;
    wire N__80773;
    wire N__80770;
    wire N__80769;
    wire N__80766;
    wire N__80763;
    wire N__80760;
    wire N__80755;
    wire N__80752;
    wire N__80749;
    wire N__80746;
    wire N__80743;
    wire N__80740;
    wire N__80737;
    wire N__80734;
    wire N__80733;
    wire N__80730;
    wire N__80727;
    wire N__80722;
    wire N__80719;
    wire N__80716;
    wire N__80713;
    wire N__80710;
    wire N__80707;
    wire N__80704;
    wire N__80701;
    wire N__80700;
    wire N__80699;
    wire N__80698;
    wire N__80697;
    wire N__80696;
    wire N__80695;
    wire N__80692;
    wire N__80691;
    wire N__80690;
    wire N__80685;
    wire N__80682;
    wire N__80681;
    wire N__80678;
    wire N__80677;
    wire N__80674;
    wire N__80671;
    wire N__80670;
    wire N__80669;
    wire N__80666;
    wire N__80663;
    wire N__80660;
    wire N__80659;
    wire N__80656;
    wire N__80653;
    wire N__80650;
    wire N__80649;
    wire N__80648;
    wire N__80645;
    wire N__80642;
    wire N__80639;
    wire N__80636;
    wire N__80631;
    wire N__80630;
    wire N__80629;
    wire N__80624;
    wire N__80621;
    wire N__80620;
    wire N__80619;
    wire N__80616;
    wire N__80613;
    wire N__80610;
    wire N__80607;
    wire N__80602;
    wire N__80599;
    wire N__80596;
    wire N__80593;
    wire N__80588;
    wire N__80583;
    wire N__80578;
    wire N__80573;
    wire N__80570;
    wire N__80561;
    wire N__80558;
    wire N__80555;
    wire N__80550;
    wire N__80543;
    wire N__80538;
    wire N__80527;
    wire N__80524;
    wire N__80521;
    wire N__80518;
    wire N__80515;
    wire N__80512;
    wire N__80509;
    wire N__80506;
    wire N__80503;
    wire N__80500;
    wire N__80497;
    wire N__80494;
    wire N__80491;
    wire N__80490;
    wire N__80489;
    wire N__80486;
    wire N__80483;
    wire N__80480;
    wire N__80479;
    wire N__80476;
    wire N__80473;
    wire N__80472;
    wire N__80469;
    wire N__80466;
    wire N__80465;
    wire N__80462;
    wire N__80459;
    wire N__80456;
    wire N__80455;
    wire N__80454;
    wire N__80451;
    wire N__80446;
    wire N__80443;
    wire N__80438;
    wire N__80433;
    wire N__80428;
    wire N__80419;
    wire N__80418;
    wire N__80417;
    wire N__80414;
    wire N__80411;
    wire N__80410;
    wire N__80409;
    wire N__80408;
    wire N__80407;
    wire N__80404;
    wire N__80401;
    wire N__80398;
    wire N__80395;
    wire N__80388;
    wire N__80385;
    wire N__80380;
    wire N__80377;
    wire N__80376;
    wire N__80371;
    wire N__80370;
    wire N__80369;
    wire N__80366;
    wire N__80363;
    wire N__80360;
    wire N__80357;
    wire N__80352;
    wire N__80341;
    wire N__80340;
    wire N__80339;
    wire N__80336;
    wire N__80333;
    wire N__80330;
    wire N__80325;
    wire N__80320;
    wire N__80317;
    wire N__80314;
    wire N__80313;
    wire N__80312;
    wire N__80311;
    wire N__80310;
    wire N__80307;
    wire N__80304;
    wire N__80303;
    wire N__80300;
    wire N__80297;
    wire N__80294;
    wire N__80291;
    wire N__80288;
    wire N__80287;
    wire N__80284;
    wire N__80283;
    wire N__80282;
    wire N__80281;
    wire N__80278;
    wire N__80273;
    wire N__80268;
    wire N__80265;
    wire N__80262;
    wire N__80257;
    wire N__80254;
    wire N__80253;
    wire N__80248;
    wire N__80243;
    wire N__80240;
    wire N__80237;
    wire N__80232;
    wire N__80229;
    wire N__80218;
    wire N__80217;
    wire N__80216;
    wire N__80215;
    wire N__80214;
    wire N__80213;
    wire N__80208;
    wire N__80207;
    wire N__80206;
    wire N__80205;
    wire N__80204;
    wire N__80199;
    wire N__80198;
    wire N__80195;
    wire N__80194;
    wire N__80193;
    wire N__80192;
    wire N__80189;
    wire N__80188;
    wire N__80187;
    wire N__80184;
    wire N__80179;
    wire N__80176;
    wire N__80173;
    wire N__80170;
    wire N__80167;
    wire N__80158;
    wire N__80155;
    wire N__80152;
    wire N__80149;
    wire N__80142;
    wire N__80139;
    wire N__80136;
    wire N__80135;
    wire N__80130;
    wire N__80121;
    wire N__80120;
    wire N__80119;
    wire N__80114;
    wire N__80111;
    wire N__80108;
    wire N__80105;
    wire N__80100;
    wire N__80089;
    wire N__80086;
    wire N__80083;
    wire N__80080;
    wire N__80079;
    wire N__80074;
    wire N__80073;
    wire N__80070;
    wire N__80067;
    wire N__80064;
    wire N__80059;
    wire N__80056;
    wire N__80053;
    wire N__80052;
    wire N__80051;
    wire N__80048;
    wire N__80045;
    wire N__80042;
    wire N__80039;
    wire N__80032;
    wire N__80029;
    wire N__80026;
    wire N__80023;
    wire N__80020;
    wire N__80017;
    wire N__80014;
    wire N__80013;
    wire N__80012;
    wire N__80011;
    wire N__80008;
    wire N__80005;
    wire N__80004;
    wire N__80003;
    wire N__80002;
    wire N__79999;
    wire N__79998;
    wire N__79995;
    wire N__79992;
    wire N__79989;
    wire N__79986;
    wire N__79983;
    wire N__79980;
    wire N__79977;
    wire N__79974;
    wire N__79973;
    wire N__79972;
    wire N__79971;
    wire N__79968;
    wire N__79965;
    wire N__79962;
    wire N__79957;
    wire N__79954;
    wire N__79949;
    wire N__79942;
    wire N__79939;
    wire N__79932;
    wire N__79927;
    wire N__79922;
    wire N__79915;
    wire N__79914;
    wire N__79913;
    wire N__79912;
    wire N__79909;
    wire N__79906;
    wire N__79905;
    wire N__79904;
    wire N__79903;
    wire N__79900;
    wire N__79897;
    wire N__79894;
    wire N__79891;
    wire N__79890;
    wire N__79885;
    wire N__79884;
    wire N__79883;
    wire N__79880;
    wire N__79877;
    wire N__79874;
    wire N__79871;
    wire N__79868;
    wire N__79865;
    wire N__79862;
    wire N__79857;
    wire N__79856;
    wire N__79855;
    wire N__79852;
    wire N__79847;
    wire N__79844;
    wire N__79841;
    wire N__79838;
    wire N__79835;
    wire N__79832;
    wire N__79829;
    wire N__79826;
    wire N__79821;
    wire N__79818;
    wire N__79815;
    wire N__79812;
    wire N__79809;
    wire N__79806;
    wire N__79803;
    wire N__79794;
    wire N__79783;
    wire N__79782;
    wire N__79779;
    wire N__79776;
    wire N__79773;
    wire N__79770;
    wire N__79767;
    wire N__79764;
    wire N__79759;
    wire N__79756;
    wire N__79753;
    wire N__79750;
    wire N__79747;
    wire N__79744;
    wire N__79741;
    wire N__79738;
    wire N__79737;
    wire N__79734;
    wire N__79731;
    wire N__79728;
    wire N__79725;
    wire N__79722;
    wire N__79717;
    wire N__79714;
    wire N__79711;
    wire N__79710;
    wire N__79707;
    wire N__79704;
    wire N__79701;
    wire N__79696;
    wire N__79693;
    wire N__79690;
    wire N__79687;
    wire N__79684;
    wire N__79681;
    wire N__79678;
    wire N__79675;
    wire N__79672;
    wire N__79669;
    wire N__79666;
    wire N__79663;
    wire N__79660;
    wire N__79659;
    wire N__79656;
    wire N__79655;
    wire N__79654;
    wire N__79651;
    wire N__79650;
    wire N__79647;
    wire N__79644;
    wire N__79641;
    wire N__79638;
    wire N__79635;
    wire N__79630;
    wire N__79627;
    wire N__79626;
    wire N__79625;
    wire N__79622;
    wire N__79619;
    wire N__79616;
    wire N__79613;
    wire N__79612;
    wire N__79609;
    wire N__79606;
    wire N__79603;
    wire N__79596;
    wire N__79591;
    wire N__79588;
    wire N__79579;
    wire N__79576;
    wire N__79575;
    wire N__79572;
    wire N__79569;
    wire N__79566;
    wire N__79561;
    wire N__79558;
    wire N__79555;
    wire N__79552;
    wire N__79549;
    wire N__79546;
    wire N__79543;
    wire N__79540;
    wire N__79537;
    wire N__79534;
    wire N__79531;
    wire N__79528;
    wire N__79527;
    wire N__79522;
    wire N__79519;
    wire N__79516;
    wire N__79513;
    wire N__79510;
    wire N__79507;
    wire N__79504;
    wire N__79501;
    wire N__79498;
    wire N__79495;
    wire N__79492;
    wire N__79489;
    wire N__79486;
    wire N__79483;
    wire N__79480;
    wire N__79477;
    wire N__79474;
    wire N__79471;
    wire N__79468;
    wire N__79467;
    wire N__79466;
    wire N__79463;
    wire N__79460;
    wire N__79457;
    wire N__79454;
    wire N__79453;
    wire N__79452;
    wire N__79447;
    wire N__79446;
    wire N__79445;
    wire N__79442;
    wire N__79437;
    wire N__79434;
    wire N__79429;
    wire N__79420;
    wire N__79417;
    wire N__79414;
    wire N__79411;
    wire N__79408;
    wire N__79405;
    wire N__79402;
    wire N__79399;
    wire N__79398;
    wire N__79395;
    wire N__79392;
    wire N__79387;
    wire N__79386;
    wire N__79385;
    wire N__79384;
    wire N__79381;
    wire N__79374;
    wire N__79369;
    wire N__79366;
    wire N__79363;
    wire N__79360;
    wire N__79357;
    wire N__79354;
    wire N__79351;
    wire N__79348;
    wire N__79345;
    wire N__79344;
    wire N__79341;
    wire N__79338;
    wire N__79335;
    wire N__79332;
    wire N__79327;
    wire N__79326;
    wire N__79325;
    wire N__79322;
    wire N__79317;
    wire N__79316;
    wire N__79313;
    wire N__79310;
    wire N__79307;
    wire N__79302;
    wire N__79297;
    wire N__79294;
    wire N__79291;
    wire N__79288;
    wire N__79285;
    wire N__79284;
    wire N__79279;
    wire N__79276;
    wire N__79275;
    wire N__79272;
    wire N__79269;
    wire N__79264;
    wire N__79261;
    wire N__79258;
    wire N__79255;
    wire N__79252;
    wire N__79249;
    wire N__79248;
    wire N__79243;
    wire N__79240;
    wire N__79237;
    wire N__79234;
    wire N__79231;
    wire N__79228;
    wire N__79225;
    wire N__79224;
    wire N__79223;
    wire N__79222;
    wire N__79221;
    wire N__79214;
    wire N__79209;
    wire N__79206;
    wire N__79203;
    wire N__79198;
    wire N__79195;
    wire N__79192;
    wire N__79189;
    wire N__79186;
    wire N__79185;
    wire N__79184;
    wire N__79177;
    wire N__79174;
    wire N__79173;
    wire N__79170;
    wire N__79169;
    wire N__79168;
    wire N__79165;
    wire N__79162;
    wire N__79157;
    wire N__79154;
    wire N__79149;
    wire N__79144;
    wire N__79141;
    wire N__79138;
    wire N__79135;
    wire N__79132;
    wire N__79129;
    wire N__79126;
    wire N__79123;
    wire N__79122;
    wire N__79121;
    wire N__79120;
    wire N__79119;
    wire N__79118;
    wire N__79113;
    wire N__79110;
    wire N__79107;
    wire N__79106;
    wire N__79105;
    wire N__79100;
    wire N__79095;
    wire N__79088;
    wire N__79081;
    wire N__79078;
    wire N__79075;
    wire N__79072;
    wire N__79069;
    wire N__79066;
    wire N__79063;
    wire N__79060;
    wire N__79057;
    wire N__79054;
    wire N__79053;
    wire N__79048;
    wire N__79047;
    wire N__79046;
    wire N__79043;
    wire N__79038;
    wire N__79033;
    wire N__79030;
    wire N__79027;
    wire N__79024;
    wire N__79021;
    wire N__79018;
    wire N__79015;
    wire N__79014;
    wire N__79011;
    wire N__79008;
    wire N__79005;
    wire N__79002;
    wire N__78999;
    wire N__78996;
    wire N__78993;
    wire N__78988;
    wire N__78985;
    wire N__78982;
    wire N__78979;
    wire N__78976;
    wire N__78973;
    wire N__78970;
    wire N__78967;
    wire N__78964;
    wire N__78961;
    wire N__78960;
    wire N__78959;
    wire N__78954;
    wire N__78951;
    wire N__78948;
    wire N__78945;
    wire N__78942;
    wire N__78937;
    wire N__78934;
    wire N__78931;
    wire N__78928;
    wire N__78927;
    wire N__78924;
    wire N__78921;
    wire N__78918;
    wire N__78913;
    wire N__78912;
    wire N__78907;
    wire N__78904;
    wire N__78903;
    wire N__78900;
    wire N__78897;
    wire N__78894;
    wire N__78889;
    wire N__78886;
    wire N__78885;
    wire N__78880;
    wire N__78877;
    wire N__78876;
    wire N__78871;
    wire N__78868;
    wire N__78865;
    wire N__78862;
    wire N__78859;
    wire N__78856;
    wire N__78853;
    wire N__78850;
    wire N__78847;
    wire N__78844;
    wire N__78841;
    wire N__78838;
    wire N__78835;
    wire N__78832;
    wire N__78829;
    wire N__78826;
    wire N__78823;
    wire N__78820;
    wire N__78817;
    wire N__78814;
    wire N__78811;
    wire N__78808;
    wire N__78807;
    wire N__78806;
    wire N__78805;
    wire N__78800;
    wire N__78797;
    wire N__78794;
    wire N__78791;
    wire N__78786;
    wire N__78781;
    wire N__78778;
    wire N__78775;
    wire N__78772;
    wire N__78769;
    wire N__78768;
    wire N__78767;
    wire N__78760;
    wire N__78757;
    wire N__78754;
    wire N__78751;
    wire N__78748;
    wire N__78745;
    wire N__78742;
    wire N__78739;
    wire N__78738;
    wire N__78737;
    wire N__78736;
    wire N__78733;
    wire N__78728;
    wire N__78727;
    wire N__78724;
    wire N__78719;
    wire N__78714;
    wire N__78711;
    wire N__78708;
    wire N__78703;
    wire N__78702;
    wire N__78699;
    wire N__78696;
    wire N__78695;
    wire N__78694;
    wire N__78691;
    wire N__78690;
    wire N__78689;
    wire N__78686;
    wire N__78683;
    wire N__78682;
    wire N__78679;
    wire N__78676;
    wire N__78673;
    wire N__78670;
    wire N__78667;
    wire N__78662;
    wire N__78649;
    wire N__78646;
    wire N__78643;
    wire N__78640;
    wire N__78637;
    wire N__78634;
    wire N__78631;
    wire N__78628;
    wire N__78625;
    wire N__78622;
    wire N__78621;
    wire N__78618;
    wire N__78615;
    wire N__78614;
    wire N__78613;
    wire N__78608;
    wire N__78607;
    wire N__78606;
    wire N__78603;
    wire N__78600;
    wire N__78597;
    wire N__78594;
    wire N__78591;
    wire N__78588;
    wire N__78585;
    wire N__78574;
    wire N__78571;
    wire N__78568;
    wire N__78565;
    wire N__78562;
    wire N__78559;
    wire N__78556;
    wire N__78555;
    wire N__78554;
    wire N__78553;
    wire N__78544;
    wire N__78543;
    wire N__78542;
    wire N__78539;
    wire N__78536;
    wire N__78533;
    wire N__78530;
    wire N__78527;
    wire N__78524;
    wire N__78517;
    wire N__78514;
    wire N__78511;
    wire N__78510;
    wire N__78507;
    wire N__78504;
    wire N__78503;
    wire N__78502;
    wire N__78501;
    wire N__78500;
    wire N__78499;
    wire N__78498;
    wire N__78497;
    wire N__78496;
    wire N__78491;
    wire N__78488;
    wire N__78485;
    wire N__78482;
    wire N__78477;
    wire N__78474;
    wire N__78469;
    wire N__78468;
    wire N__78465;
    wire N__78460;
    wire N__78453;
    wire N__78450;
    wire N__78447;
    wire N__78440;
    wire N__78439;
    wire N__78436;
    wire N__78433;
    wire N__78430;
    wire N__78427;
    wire N__78418;
    wire N__78417;
    wire N__78414;
    wire N__78413;
    wire N__78412;
    wire N__78409;
    wire N__78406;
    wire N__78403;
    wire N__78400;
    wire N__78397;
    wire N__78396;
    wire N__78395;
    wire N__78392;
    wire N__78391;
    wire N__78388;
    wire N__78383;
    wire N__78380;
    wire N__78377;
    wire N__78376;
    wire N__78373;
    wire N__78370;
    wire N__78367;
    wire N__78362;
    wire N__78357;
    wire N__78354;
    wire N__78351;
    wire N__78348;
    wire N__78345;
    wire N__78342;
    wire N__78337;
    wire N__78328;
    wire N__78325;
    wire N__78324;
    wire N__78323;
    wire N__78320;
    wire N__78319;
    wire N__78316;
    wire N__78313;
    wire N__78312;
    wire N__78311;
    wire N__78308;
    wire N__78307;
    wire N__78306;
    wire N__78305;
    wire N__78304;
    wire N__78301;
    wire N__78298;
    wire N__78295;
    wire N__78290;
    wire N__78287;
    wire N__78282;
    wire N__78281;
    wire N__78276;
    wire N__78275;
    wire N__78274;
    wire N__78271;
    wire N__78268;
    wire N__78263;
    wire N__78260;
    wire N__78257;
    wire N__78254;
    wire N__78251;
    wire N__78246;
    wire N__78243;
    wire N__78240;
    wire N__78237;
    wire N__78234;
    wire N__78231;
    wire N__78224;
    wire N__78221;
    wire N__78218;
    wire N__78205;
    wire N__78202;
    wire N__78199;
    wire N__78196;
    wire N__78193;
    wire N__78190;
    wire N__78187;
    wire N__78184;
    wire N__78181;
    wire N__78178;
    wire N__78175;
    wire N__78172;
    wire N__78169;
    wire N__78166;
    wire N__78163;
    wire N__78160;
    wire N__78157;
    wire N__78154;
    wire N__78151;
    wire N__78148;
    wire N__78147;
    wire N__78146;
    wire N__78143;
    wire N__78142;
    wire N__78141;
    wire N__78138;
    wire N__78137;
    wire N__78136;
    wire N__78135;
    wire N__78132;
    wire N__78131;
    wire N__78130;
    wire N__78129;
    wire N__78126;
    wire N__78123;
    wire N__78120;
    wire N__78117;
    wire N__78114;
    wire N__78111;
    wire N__78110;
    wire N__78107;
    wire N__78106;
    wire N__78105;
    wire N__78102;
    wire N__78099;
    wire N__78096;
    wire N__78093;
    wire N__78088;
    wire N__78085;
    wire N__78080;
    wire N__78077;
    wire N__78074;
    wire N__78071;
    wire N__78070;
    wire N__78067;
    wire N__78064;
    wire N__78059;
    wire N__78054;
    wire N__78051;
    wire N__78048;
    wire N__78043;
    wire N__78038;
    wire N__78035;
    wire N__78030;
    wire N__78027;
    wire N__78022;
    wire N__78015;
    wire N__78014;
    wire N__78011;
    wire N__78006;
    wire N__78001;
    wire N__77998;
    wire N__77993;
    wire N__77990;
    wire N__77983;
    wire N__77982;
    wire N__77981;
    wire N__77978;
    wire N__77975;
    wire N__77974;
    wire N__77973;
    wire N__77972;
    wire N__77969;
    wire N__77968;
    wire N__77967;
    wire N__77966;
    wire N__77963;
    wire N__77960;
    wire N__77959;
    wire N__77956;
    wire N__77953;
    wire N__77950;
    wire N__77947;
    wire N__77944;
    wire N__77939;
    wire N__77936;
    wire N__77933;
    wire N__77930;
    wire N__77927;
    wire N__77924;
    wire N__77921;
    wire N__77914;
    wire N__77911;
    wire N__77908;
    wire N__77905;
    wire N__77902;
    wire N__77895;
    wire N__77892;
    wire N__77889;
    wire N__77884;
    wire N__77881;
    wire N__77872;
    wire N__77871;
    wire N__77868;
    wire N__77867;
    wire N__77864;
    wire N__77861;
    wire N__77858;
    wire N__77857;
    wire N__77856;
    wire N__77855;
    wire N__77854;
    wire N__77853;
    wire N__77850;
    wire N__77849;
    wire N__77848;
    wire N__77845;
    wire N__77842;
    wire N__77839;
    wire N__77836;
    wire N__77831;
    wire N__77828;
    wire N__77825;
    wire N__77820;
    wire N__77817;
    wire N__77814;
    wire N__77811;
    wire N__77810;
    wire N__77807;
    wire N__77804;
    wire N__77801;
    wire N__77796;
    wire N__77793;
    wire N__77790;
    wire N__77787;
    wire N__77784;
    wire N__77783;
    wire N__77782;
    wire N__77777;
    wire N__77772;
    wire N__77763;
    wire N__77758;
    wire N__77749;
    wire N__77748;
    wire N__77747;
    wire N__77744;
    wire N__77743;
    wire N__77740;
    wire N__77739;
    wire N__77736;
    wire N__77733;
    wire N__77732;
    wire N__77729;
    wire N__77726;
    wire N__77723;
    wire N__77722;
    wire N__77719;
    wire N__77716;
    wire N__77713;
    wire N__77710;
    wire N__77705;
    wire N__77702;
    wire N__77699;
    wire N__77696;
    wire N__77691;
    wire N__77688;
    wire N__77685;
    wire N__77684;
    wire N__77683;
    wire N__77680;
    wire N__77675;
    wire N__77670;
    wire N__77665;
    wire N__77656;
    wire N__77653;
    wire N__77650;
    wire N__77647;
    wire N__77644;
    wire N__77641;
    wire N__77638;
    wire N__77635;
    wire N__77632;
    wire N__77629;
    wire N__77626;
    wire N__77623;
    wire N__77622;
    wire N__77619;
    wire N__77616;
    wire N__77613;
    wire N__77612;
    wire N__77609;
    wire N__77606;
    wire N__77605;
    wire N__77602;
    wire N__77597;
    wire N__77594;
    wire N__77587;
    wire N__77584;
    wire N__77581;
    wire N__77578;
    wire N__77575;
    wire N__77574;
    wire N__77571;
    wire N__77568;
    wire N__77563;
    wire N__77560;
    wire N__77557;
    wire N__77554;
    wire N__77551;
    wire N__77548;
    wire N__77545;
    wire N__77542;
    wire N__77539;
    wire N__77536;
    wire N__77533;
    wire N__77530;
    wire N__77527;
    wire N__77524;
    wire N__77521;
    wire N__77518;
    wire N__77515;
    wire N__77512;
    wire N__77509;
    wire N__77506;
    wire N__77503;
    wire N__77500;
    wire N__77497;
    wire N__77494;
    wire N__77491;
    wire N__77488;
    wire N__77485;
    wire N__77482;
    wire N__77481;
    wire N__77478;
    wire N__77475;
    wire N__77472;
    wire N__77469;
    wire N__77466;
    wire N__77465;
    wire N__77462;
    wire N__77459;
    wire N__77456;
    wire N__77449;
    wire N__77446;
    wire N__77443;
    wire N__77440;
    wire N__77437;
    wire N__77434;
    wire N__77431;
    wire N__77428;
    wire N__77427;
    wire N__77424;
    wire N__77421;
    wire N__77416;
    wire N__77413;
    wire N__77410;
    wire N__77407;
    wire N__77404;
    wire N__77401;
    wire N__77398;
    wire N__77395;
    wire N__77392;
    wire N__77389;
    wire N__77386;
    wire N__77385;
    wire N__77382;
    wire N__77377;
    wire N__77374;
    wire N__77371;
    wire N__77368;
    wire N__77367;
    wire N__77364;
    wire N__77361;
    wire N__77358;
    wire N__77355;
    wire N__77352;
    wire N__77347;
    wire N__77344;
    wire N__77341;
    wire N__77338;
    wire N__77335;
    wire N__77332;
    wire N__77329;
    wire N__77326;
    wire N__77323;
    wire N__77320;
    wire N__77317;
    wire N__77314;
    wire N__77311;
    wire N__77308;
    wire N__77305;
    wire N__77302;
    wire N__77299;
    wire N__77296;
    wire N__77293;
    wire N__77290;
    wire N__77287;
    wire N__77284;
    wire N__77281;
    wire N__77278;
    wire N__77275;
    wire N__77272;
    wire N__77269;
    wire N__77266;
    wire N__77263;
    wire N__77260;
    wire N__77257;
    wire N__77254;
    wire N__77251;
    wire N__77248;
    wire N__77245;
    wire N__77242;
    wire N__77239;
    wire N__77236;
    wire N__77233;
    wire N__77232;
    wire N__77231;
    wire N__77228;
    wire N__77225;
    wire N__77224;
    wire N__77223;
    wire N__77222;
    wire N__77219;
    wire N__77218;
    wire N__77215;
    wire N__77212;
    wire N__77207;
    wire N__77204;
    wire N__77201;
    wire N__77198;
    wire N__77195;
    wire N__77192;
    wire N__77189;
    wire N__77182;
    wire N__77177;
    wire N__77174;
    wire N__77171;
    wire N__77164;
    wire N__77161;
    wire N__77158;
    wire N__77155;
    wire N__77152;
    wire N__77149;
    wire N__77146;
    wire N__77143;
    wire N__77140;
    wire N__77137;
    wire N__77134;
    wire N__77131;
    wire N__77128;
    wire N__77125;
    wire N__77122;
    wire N__77119;
    wire N__77116;
    wire N__77113;
    wire N__77110;
    wire N__77107;
    wire N__77104;
    wire N__77101;
    wire N__77098;
    wire N__77095;
    wire N__77092;
    wire N__77089;
    wire N__77088;
    wire N__77085;
    wire N__77084;
    wire N__77083;
    wire N__77080;
    wire N__77079;
    wire N__77076;
    wire N__77073;
    wire N__77070;
    wire N__77067;
    wire N__77064;
    wire N__77059;
    wire N__77054;
    wire N__77047;
    wire N__77044;
    wire N__77041;
    wire N__77038;
    wire N__77035;
    wire N__77032;
    wire N__77029;
    wire N__77028;
    wire N__77025;
    wire N__77022;
    wire N__77017;
    wire N__77014;
    wire N__77011;
    wire N__77008;
    wire N__77005;
    wire N__77002;
    wire N__76999;
    wire N__76996;
    wire N__76993;
    wire N__76990;
    wire N__76987;
    wire N__76984;
    wire N__76981;
    wire N__76978;
    wire N__76975;
    wire N__76972;
    wire N__76969;
    wire N__76966;
    wire N__76963;
    wire N__76960;
    wire N__76957;
    wire N__76956;
    wire N__76955;
    wire N__76954;
    wire N__76951;
    wire N__76948;
    wire N__76945;
    wire N__76942;
    wire N__76939;
    wire N__76936;
    wire N__76933;
    wire N__76930;
    wire N__76927;
    wire N__76920;
    wire N__76915;
    wire N__76912;
    wire N__76909;
    wire N__76906;
    wire N__76903;
    wire N__76900;
    wire N__76897;
    wire N__76896;
    wire N__76895;
    wire N__76892;
    wire N__76889;
    wire N__76886;
    wire N__76881;
    wire N__76878;
    wire N__76877;
    wire N__76876;
    wire N__76875;
    wire N__76870;
    wire N__76869;
    wire N__76868;
    wire N__76867;
    wire N__76866;
    wire N__76865;
    wire N__76864;
    wire N__76861;
    wire N__76856;
    wire N__76855;
    wire N__76852;
    wire N__76849;
    wire N__76846;
    wire N__76843;
    wire N__76840;
    wire N__76837;
    wire N__76834;
    wire N__76829;
    wire N__76826;
    wire N__76821;
    wire N__76820;
    wire N__76817;
    wire N__76814;
    wire N__76805;
    wire N__76802;
    wire N__76799;
    wire N__76796;
    wire N__76793;
    wire N__76790;
    wire N__76787;
    wire N__76780;
    wire N__76773;
    wire N__76770;
    wire N__76765;
    wire N__76762;
    wire N__76759;
    wire N__76756;
    wire N__76753;
    wire N__76750;
    wire N__76747;
    wire N__76744;
    wire N__76741;
    wire N__76738;
    wire N__76735;
    wire N__76734;
    wire N__76729;
    wire N__76726;
    wire N__76725;
    wire N__76724;
    wire N__76721;
    wire N__76716;
    wire N__76711;
    wire N__76710;
    wire N__76705;
    wire N__76702;
    wire N__76699;
    wire N__76698;
    wire N__76695;
    wire N__76692;
    wire N__76689;
    wire N__76686;
    wire N__76683;
    wire N__76680;
    wire N__76675;
    wire N__76672;
    wire N__76669;
    wire N__76666;
    wire N__76663;
    wire N__76660;
    wire N__76657;
    wire N__76656;
    wire N__76655;
    wire N__76652;
    wire N__76649;
    wire N__76648;
    wire N__76647;
    wire N__76644;
    wire N__76641;
    wire N__76638;
    wire N__76635;
    wire N__76632;
    wire N__76629;
    wire N__76618;
    wire N__76615;
    wire N__76612;
    wire N__76609;
    wire N__76606;
    wire N__76603;
    wire N__76600;
    wire N__76597;
    wire N__76594;
    wire N__76591;
    wire N__76588;
    wire N__76585;
    wire N__76582;
    wire N__76579;
    wire N__76576;
    wire N__76573;
    wire N__76570;
    wire N__76567;
    wire N__76564;
    wire N__76561;
    wire N__76558;
    wire N__76555;
    wire N__76552;
    wire N__76551;
    wire N__76548;
    wire N__76545;
    wire N__76542;
    wire N__76539;
    wire N__76536;
    wire N__76535;
    wire N__76530;
    wire N__76527;
    wire N__76522;
    wire N__76519;
    wire N__76516;
    wire N__76513;
    wire N__76512;
    wire N__76511;
    wire N__76510;
    wire N__76507;
    wire N__76504;
    wire N__76499;
    wire N__76494;
    wire N__76491;
    wire N__76486;
    wire N__76485;
    wire N__76482;
    wire N__76479;
    wire N__76476;
    wire N__76471;
    wire N__76468;
    wire N__76465;
    wire N__76462;
    wire N__76459;
    wire N__76456;
    wire N__76453;
    wire N__76450;
    wire N__76449;
    wire N__76446;
    wire N__76443;
    wire N__76440;
    wire N__76439;
    wire N__76436;
    wire N__76433;
    wire N__76430;
    wire N__76427;
    wire N__76424;
    wire N__76419;
    wire N__76414;
    wire N__76411;
    wire N__76408;
    wire N__76405;
    wire N__76402;
    wire N__76399;
    wire N__76396;
    wire N__76393;
    wire N__76390;
    wire N__76387;
    wire N__76384;
    wire N__76381;
    wire N__76378;
    wire N__76375;
    wire N__76372;
    wire N__76371;
    wire N__76366;
    wire N__76363;
    wire N__76360;
    wire N__76357;
    wire N__76354;
    wire N__76353;
    wire N__76352;
    wire N__76349;
    wire N__76344;
    wire N__76341;
    wire N__76338;
    wire N__76333;
    wire N__76330;
    wire N__76327;
    wire N__76324;
    wire N__76321;
    wire N__76318;
    wire N__76317;
    wire N__76314;
    wire N__76311;
    wire N__76306;
    wire N__76303;
    wire N__76300;
    wire N__76297;
    wire N__76296;
    wire N__76291;
    wire N__76288;
    wire N__76285;
    wire N__76284;
    wire N__76283;
    wire N__76280;
    wire N__76277;
    wire N__76274;
    wire N__76273;
    wire N__76272;
    wire N__76265;
    wire N__76262;
    wire N__76259;
    wire N__76254;
    wire N__76249;
    wire N__76246;
    wire N__76243;
    wire N__76240;
    wire N__76237;
    wire N__76234;
    wire N__76231;
    wire N__76228;
    wire N__76227;
    wire N__76226;
    wire N__76223;
    wire N__76220;
    wire N__76217;
    wire N__76216;
    wire N__76213;
    wire N__76210;
    wire N__76205;
    wire N__76202;
    wire N__76197;
    wire N__76192;
    wire N__76189;
    wire N__76188;
    wire N__76185;
    wire N__76182;
    wire N__76179;
    wire N__76176;
    wire N__76171;
    wire N__76168;
    wire N__76165;
    wire N__76162;
    wire N__76159;
    wire N__76158;
    wire N__76155;
    wire N__76152;
    wire N__76147;
    wire N__76144;
    wire N__76141;
    wire N__76140;
    wire N__76137;
    wire N__76134;
    wire N__76129;
    wire N__76126;
    wire N__76123;
    wire N__76120;
    wire N__76119;
    wire N__76114;
    wire N__76111;
    wire N__76108;
    wire N__76105;
    wire N__76102;
    wire N__76099;
    wire N__76096;
    wire N__76093;
    wire N__76090;
    wire N__76087;
    wire N__76084;
    wire N__76081;
    wire N__76078;
    wire N__76075;
    wire N__76072;
    wire N__76071;
    wire N__76068;
    wire N__76065;
    wire N__76060;
    wire N__76059;
    wire N__76056;
    wire N__76053;
    wire N__76052;
    wire N__76051;
    wire N__76048;
    wire N__76045;
    wire N__76040;
    wire N__76035;
    wire N__76032;
    wire N__76027;
    wire N__76024;
    wire N__76021;
    wire N__76018;
    wire N__76015;
    wire N__76012;
    wire N__76011;
    wire N__76010;
    wire N__76009;
    wire N__76004;
    wire N__76001;
    wire N__76000;
    wire N__75999;
    wire N__75998;
    wire N__75995;
    wire N__75990;
    wire N__75983;
    wire N__75980;
    wire N__75977;
    wire N__75972;
    wire N__75967;
    wire N__75966;
    wire N__75965;
    wire N__75964;
    wire N__75963;
    wire N__75962;
    wire N__75959;
    wire N__75958;
    wire N__75957;
    wire N__75956;
    wire N__75953;
    wire N__75946;
    wire N__75943;
    wire N__75942;
    wire N__75941;
    wire N__75940;
    wire N__75939;
    wire N__75934;
    wire N__75933;
    wire N__75930;
    wire N__75927;
    wire N__75922;
    wire N__75913;
    wire N__75910;
    wire N__75909;
    wire N__75906;
    wire N__75903;
    wire N__75898;
    wire N__75895;
    wire N__75892;
    wire N__75887;
    wire N__75884;
    wire N__75877;
    wire N__75868;
    wire N__75867;
    wire N__75866;
    wire N__75865;
    wire N__75862;
    wire N__75861;
    wire N__75854;
    wire N__75851;
    wire N__75850;
    wire N__75849;
    wire N__75846;
    wire N__75843;
    wire N__75840;
    wire N__75837;
    wire N__75832;
    wire N__75829;
    wire N__75826;
    wire N__75821;
    wire N__75818;
    wire N__75813;
    wire N__75810;
    wire N__75807;
    wire N__75804;
    wire N__75801;
    wire N__75796;
    wire N__75793;
    wire N__75792;
    wire N__75791;
    wire N__75784;
    wire N__75781;
    wire N__75778;
    wire N__75775;
    wire N__75772;
    wire N__75769;
    wire N__75768;
    wire N__75767;
    wire N__75766;
    wire N__75765;
    wire N__75764;
    wire N__75761;
    wire N__75758;
    wire N__75755;
    wire N__75752;
    wire N__75749;
    wire N__75746;
    wire N__75743;
    wire N__75738;
    wire N__75735;
    wire N__75732;
    wire N__75729;
    wire N__75726;
    wire N__75723;
    wire N__75720;
    wire N__75717;
    wire N__75710;
    wire N__75707;
    wire N__75700;
    wire N__75697;
    wire N__75696;
    wire N__75695;
    wire N__75692;
    wire N__75687;
    wire N__75684;
    wire N__75681;
    wire N__75676;
    wire N__75675;
    wire N__75672;
    wire N__75671;
    wire N__75670;
    wire N__75669;
    wire N__75666;
    wire N__75661;
    wire N__75658;
    wire N__75655;
    wire N__75654;
    wire N__75653;
    wire N__75652;
    wire N__75651;
    wire N__75646;
    wire N__75641;
    wire N__75636;
    wire N__75631;
    wire N__75628;
    wire N__75625;
    wire N__75616;
    wire N__75615;
    wire N__75614;
    wire N__75611;
    wire N__75608;
    wire N__75605;
    wire N__75602;
    wire N__75599;
    wire N__75596;
    wire N__75593;
    wire N__75590;
    wire N__75587;
    wire N__75580;
    wire N__75577;
    wire N__75574;
    wire N__75571;
    wire N__75568;
    wire N__75565;
    wire N__75564;
    wire N__75561;
    wire N__75558;
    wire N__75557;
    wire N__75554;
    wire N__75551;
    wire N__75548;
    wire N__75543;
    wire N__75540;
    wire N__75537;
    wire N__75532;
    wire N__75529;
    wire N__75526;
    wire N__75523;
    wire N__75520;
    wire N__75517;
    wire N__75514;
    wire N__75511;
    wire N__75510;
    wire N__75509;
    wire N__75506;
    wire N__75501;
    wire N__75498;
    wire N__75495;
    wire N__75492;
    wire N__75489;
    wire N__75484;
    wire N__75483;
    wire N__75480;
    wire N__75477;
    wire N__75472;
    wire N__75471;
    wire N__75470;
    wire N__75467;
    wire N__75462;
    wire N__75459;
    wire N__75456;
    wire N__75451;
    wire N__75450;
    wire N__75449;
    wire N__75446;
    wire N__75443;
    wire N__75440;
    wire N__75437;
    wire N__75434;
    wire N__75431;
    wire N__75428;
    wire N__75425;
    wire N__75420;
    wire N__75417;
    wire N__75412;
    wire N__75409;
    wire N__75408;
    wire N__75407;
    wire N__75404;
    wire N__75399;
    wire N__75396;
    wire N__75393;
    wire N__75390;
    wire N__75387;
    wire N__75382;
    wire N__75381;
    wire N__75380;
    wire N__75377;
    wire N__75372;
    wire N__75369;
    wire N__75366;
    wire N__75363;
    wire N__75360;
    wire N__75355;
    wire N__75354;
    wire N__75353;
    wire N__75350;
    wire N__75345;
    wire N__75342;
    wire N__75339;
    wire N__75336;
    wire N__75333;
    wire N__75328;
    wire N__75327;
    wire N__75326;
    wire N__75325;
    wire N__75324;
    wire N__75323;
    wire N__75322;
    wire N__75321;
    wire N__75320;
    wire N__75319;
    wire N__75318;
    wire N__75317;
    wire N__75316;
    wire N__75289;
    wire N__75286;
    wire N__75283;
    wire N__75282;
    wire N__75281;
    wire N__75280;
    wire N__75277;
    wire N__75274;
    wire N__75269;
    wire N__75266;
    wire N__75261;
    wire N__75258;
    wire N__75255;
    wire N__75250;
    wire N__75247;
    wire N__75244;
    wire N__75243;
    wire N__75242;
    wire N__75239;
    wire N__75236;
    wire N__75233;
    wire N__75226;
    wire N__75225;
    wire N__75224;
    wire N__75219;
    wire N__75216;
    wire N__75213;
    wire N__75210;
    wire N__75207;
    wire N__75204;
    wire N__75201;
    wire N__75196;
    wire N__75193;
    wire N__75192;
    wire N__75189;
    wire N__75188;
    wire N__75185;
    wire N__75182;
    wire N__75177;
    wire N__75172;
    wire N__75171;
    wire N__75170;
    wire N__75167;
    wire N__75162;
    wire N__75157;
    wire N__75154;
    wire N__75151;
    wire N__75148;
    wire N__75145;
    wire N__75144;
    wire N__75141;
    wire N__75138;
    wire N__75137;
    wire N__75136;
    wire N__75131;
    wire N__75126;
    wire N__75123;
    wire N__75120;
    wire N__75115;
    wire N__75112;
    wire N__75111;
    wire N__75110;
    wire N__75109;
    wire N__75108;
    wire N__75105;
    wire N__75102;
    wire N__75101;
    wire N__75100;
    wire N__75095;
    wire N__75092;
    wire N__75087;
    wire N__75082;
    wire N__75073;
    wire N__75070;
    wire N__75067;
    wire N__75064;
    wire N__75061;
    wire N__75058;
    wire N__75057;
    wire N__75056;
    wire N__75055;
    wire N__75052;
    wire N__75047;
    wire N__75044;
    wire N__75041;
    wire N__75036;
    wire N__75031;
    wire N__75028;
    wire N__75027;
    wire N__75026;
    wire N__75025;
    wire N__75024;
    wire N__75021;
    wire N__75020;
    wire N__75017;
    wire N__75014;
    wire N__75013;
    wire N__75008;
    wire N__75005;
    wire N__75002;
    wire N__74999;
    wire N__74994;
    wire N__74983;
    wire N__74980;
    wire N__74977;
    wire N__74974;
    wire N__74971;
    wire N__74968;
    wire N__74967;
    wire N__74966;
    wire N__74965;
    wire N__74964;
    wire N__74963;
    wire N__74962;
    wire N__74959;
    wire N__74958;
    wire N__74955;
    wire N__74952;
    wire N__74949;
    wire N__74946;
    wire N__74943;
    wire N__74942;
    wire N__74939;
    wire N__74936;
    wire N__74935;
    wire N__74932;
    wire N__74929;
    wire N__74920;
    wire N__74917;
    wire N__74914;
    wire N__74911;
    wire N__74908;
    wire N__74905;
    wire N__74902;
    wire N__74897;
    wire N__74890;
    wire N__74885;
    wire N__74882;
    wire N__74875;
    wire N__74872;
    wire N__74871;
    wire N__74868;
    wire N__74865;
    wire N__74862;
    wire N__74859;
    wire N__74858;
    wire N__74857;
    wire N__74856;
    wire N__74853;
    wire N__74850;
    wire N__74849;
    wire N__74846;
    wire N__74843;
    wire N__74840;
    wire N__74839;
    wire N__74836;
    wire N__74833;
    wire N__74830;
    wire N__74827;
    wire N__74824;
    wire N__74821;
    wire N__74818;
    wire N__74815;
    wire N__74814;
    wire N__74811;
    wire N__74806;
    wire N__74803;
    wire N__74800;
    wire N__74795;
    wire N__74792;
    wire N__74791;
    wire N__74788;
    wire N__74783;
    wire N__74776;
    wire N__74773;
    wire N__74768;
    wire N__74761;
    wire N__74758;
    wire N__74755;
    wire N__74752;
    wire N__74749;
    wire N__74746;
    wire N__74743;
    wire N__74740;
    wire N__74737;
    wire N__74734;
    wire N__74731;
    wire N__74728;
    wire N__74725;
    wire N__74722;
    wire N__74721;
    wire N__74718;
    wire N__74717;
    wire N__74716;
    wire N__74713;
    wire N__74710;
    wire N__74707;
    wire N__74704;
    wire N__74699;
    wire N__74692;
    wire N__74691;
    wire N__74690;
    wire N__74687;
    wire N__74684;
    wire N__74681;
    wire N__74678;
    wire N__74677;
    wire N__74674;
    wire N__74671;
    wire N__74668;
    wire N__74665;
    wire N__74662;
    wire N__74655;
    wire N__74652;
    wire N__74649;
    wire N__74644;
    wire N__74641;
    wire N__74638;
    wire N__74635;
    wire N__74632;
    wire N__74629;
    wire N__74626;
    wire N__74623;
    wire N__74620;
    wire N__74617;
    wire N__74614;
    wire N__74611;
    wire N__74608;
    wire N__74605;
    wire N__74602;
    wire N__74599;
    wire N__74596;
    wire N__74593;
    wire N__74590;
    wire N__74589;
    wire N__74588;
    wire N__74585;
    wire N__74580;
    wire N__74577;
    wire N__74574;
    wire N__74569;
    wire N__74568;
    wire N__74565;
    wire N__74564;
    wire N__74561;
    wire N__74558;
    wire N__74555;
    wire N__74552;
    wire N__74545;
    wire N__74542;
    wire N__74539;
    wire N__74536;
    wire N__74533;
    wire N__74530;
    wire N__74527;
    wire N__74524;
    wire N__74521;
    wire N__74518;
    wire N__74515;
    wire N__74514;
    wire N__74511;
    wire N__74508;
    wire N__74507;
    wire N__74506;
    wire N__74505;
    wire N__74504;
    wire N__74503;
    wire N__74500;
    wire N__74497;
    wire N__74496;
    wire N__74495;
    wire N__74494;
    wire N__74491;
    wire N__74488;
    wire N__74485;
    wire N__74480;
    wire N__74477;
    wire N__74474;
    wire N__74473;
    wire N__74470;
    wire N__74465;
    wire N__74460;
    wire N__74457;
    wire N__74454;
    wire N__74451;
    wire N__74448;
    wire N__74445;
    wire N__74442;
    wire N__74439;
    wire N__74432;
    wire N__74429;
    wire N__74426;
    wire N__74421;
    wire N__74418;
    wire N__74415;
    wire N__74404;
    wire N__74401;
    wire N__74398;
    wire N__74395;
    wire N__74392;
    wire N__74391;
    wire N__74390;
    wire N__74383;
    wire N__74380;
    wire N__74377;
    wire N__74374;
    wire N__74373;
    wire N__74372;
    wire N__74371;
    wire N__74368;
    wire N__74363;
    wire N__74360;
    wire N__74357;
    wire N__74356;
    wire N__74353;
    wire N__74350;
    wire N__74347;
    wire N__74344;
    wire N__74339;
    wire N__74332;
    wire N__74329;
    wire N__74326;
    wire N__74323;
    wire N__74320;
    wire N__74319;
    wire N__74318;
    wire N__74317;
    wire N__74314;
    wire N__74313;
    wire N__74312;
    wire N__74311;
    wire N__74308;
    wire N__74305;
    wire N__74304;
    wire N__74301;
    wire N__74300;
    wire N__74297;
    wire N__74294;
    wire N__74289;
    wire N__74284;
    wire N__74277;
    wire N__74274;
    wire N__74271;
    wire N__74270;
    wire N__74267;
    wire N__74266;
    wire N__74261;
    wire N__74258;
    wire N__74255;
    wire N__74252;
    wire N__74249;
    wire N__74246;
    wire N__74243;
    wire N__74232;
    wire N__74229;
    wire N__74224;
    wire N__74221;
    wire N__74218;
    wire N__74215;
    wire N__74214;
    wire N__74211;
    wire N__74208;
    wire N__74207;
    wire N__74202;
    wire N__74199;
    wire N__74194;
    wire N__74191;
    wire N__74188;
    wire N__74185;
    wire N__74184;
    wire N__74183;
    wire N__74180;
    wire N__74177;
    wire N__74176;
    wire N__74175;
    wire N__74172;
    wire N__74171;
    wire N__74168;
    wire N__74165;
    wire N__74164;
    wire N__74161;
    wire N__74158;
    wire N__74153;
    wire N__74150;
    wire N__74147;
    wire N__74146;
    wire N__74143;
    wire N__74138;
    wire N__74135;
    wire N__74134;
    wire N__74133;
    wire N__74132;
    wire N__74129;
    wire N__74126;
    wire N__74123;
    wire N__74116;
    wire N__74113;
    wire N__74108;
    wire N__74097;
    wire N__74094;
    wire N__74089;
    wire N__74086;
    wire N__74083;
    wire N__74082;
    wire N__74081;
    wire N__74078;
    wire N__74077;
    wire N__74076;
    wire N__74073;
    wire N__74070;
    wire N__74067;
    wire N__74066;
    wire N__74063;
    wire N__74062;
    wire N__74059;
    wire N__74056;
    wire N__74053;
    wire N__74052;
    wire N__74051;
    wire N__74048;
    wire N__74045;
    wire N__74042;
    wire N__74039;
    wire N__74034;
    wire N__74031;
    wire N__74026;
    wire N__74023;
    wire N__74020;
    wire N__74017;
    wire N__74012;
    wire N__74005;
    wire N__74002;
    wire N__73993;
    wire N__73990;
    wire N__73987;
    wire N__73984;
    wire N__73983;
    wire N__73980;
    wire N__73977;
    wire N__73972;
    wire N__73969;
    wire N__73966;
    wire N__73963;
    wire N__73960;
    wire N__73957;
    wire N__73954;
    wire N__73951;
    wire N__73948;
    wire N__73945;
    wire N__73942;
    wire N__73939;
    wire N__73936;
    wire N__73933;
    wire N__73930;
    wire N__73927;
    wire N__73924;
    wire N__73921;
    wire N__73918;
    wire N__73915;
    wire N__73912;
    wire N__73909;
    wire N__73908;
    wire N__73907;
    wire N__73906;
    wire N__73903;
    wire N__73900;
    wire N__73899;
    wire N__73898;
    wire N__73897;
    wire N__73896;
    wire N__73895;
    wire N__73894;
    wire N__73893;
    wire N__73888;
    wire N__73887;
    wire N__73884;
    wire N__73881;
    wire N__73876;
    wire N__73873;
    wire N__73864;
    wire N__73861;
    wire N__73860;
    wire N__73857;
    wire N__73854;
    wire N__73851;
    wire N__73848;
    wire N__73845;
    wire N__73840;
    wire N__73837;
    wire N__73834;
    wire N__73831;
    wire N__73828;
    wire N__73825;
    wire N__73820;
    wire N__73815;
    wire N__73810;
    wire N__73801;
    wire N__73798;
    wire N__73797;
    wire N__73796;
    wire N__73795;
    wire N__73794;
    wire N__73793;
    wire N__73790;
    wire N__73787;
    wire N__73782;
    wire N__73779;
    wire N__73776;
    wire N__73773;
    wire N__73770;
    wire N__73769;
    wire N__73766;
    wire N__73763;
    wire N__73760;
    wire N__73757;
    wire N__73754;
    wire N__73751;
    wire N__73744;
    wire N__73741;
    wire N__73738;
    wire N__73735;
    wire N__73732;
    wire N__73729;
    wire N__73726;
    wire N__73717;
    wire N__73714;
    wire N__73713;
    wire N__73710;
    wire N__73707;
    wire N__73702;
    wire N__73699;
    wire N__73698;
    wire N__73695;
    wire N__73692;
    wire N__73687;
    wire N__73686;
    wire N__73681;
    wire N__73678;
    wire N__73675;
    wire N__73672;
    wire N__73669;
    wire N__73666;
    wire N__73663;
    wire N__73660;
    wire N__73657;
    wire N__73654;
    wire N__73653;
    wire N__73650;
    wire N__73647;
    wire N__73642;
    wire N__73639;
    wire N__73636;
    wire N__73633;
    wire N__73632;
    wire N__73631;
    wire N__73628;
    wire N__73625;
    wire N__73622;
    wire N__73619;
    wire N__73616;
    wire N__73609;
    wire N__73606;
    wire N__73603;
    wire N__73600;
    wire N__73597;
    wire N__73594;
    wire N__73593;
    wire N__73590;
    wire N__73587;
    wire N__73584;
    wire N__73579;
    wire N__73576;
    wire N__73573;
    wire N__73570;
    wire N__73567;
    wire N__73564;
    wire N__73561;
    wire N__73558;
    wire N__73555;
    wire N__73552;
    wire N__73549;
    wire N__73546;
    wire N__73543;
    wire N__73542;
    wire N__73537;
    wire N__73534;
    wire N__73531;
    wire N__73528;
    wire N__73525;
    wire N__73522;
    wire N__73519;
    wire N__73516;
    wire N__73513;
    wire N__73510;
    wire N__73507;
    wire N__73504;
    wire N__73501;
    wire N__73498;
    wire N__73495;
    wire N__73492;
    wire N__73489;
    wire N__73486;
    wire N__73483;
    wire N__73480;
    wire N__73477;
    wire N__73474;
    wire N__73471;
    wire N__73468;
    wire N__73465;
    wire N__73462;
    wire N__73459;
    wire N__73456;
    wire N__73453;
    wire N__73450;
    wire N__73449;
    wire N__73446;
    wire N__73443;
    wire N__73438;
    wire N__73435;
    wire N__73432;
    wire N__73429;
    wire N__73428;
    wire N__73425;
    wire N__73422;
    wire N__73417;
    wire N__73414;
    wire N__73411;
    wire N__73408;
    wire N__73405;
    wire N__73404;
    wire N__73401;
    wire N__73398;
    wire N__73395;
    wire N__73390;
    wire N__73387;
    wire N__73384;
    wire N__73383;
    wire N__73380;
    wire N__73379;
    wire N__73376;
    wire N__73373;
    wire N__73368;
    wire N__73367;
    wire N__73364;
    wire N__73361;
    wire N__73358;
    wire N__73355;
    wire N__73350;
    wire N__73345;
    wire N__73342;
    wire N__73339;
    wire N__73336;
    wire N__73333;
    wire N__73330;
    wire N__73327;
    wire N__73324;
    wire N__73321;
    wire N__73318;
    wire N__73315;
    wire N__73312;
    wire N__73311;
    wire N__73308;
    wire N__73305;
    wire N__73300;
    wire N__73297;
    wire N__73294;
    wire N__73291;
    wire N__73288;
    wire N__73285;
    wire N__73282;
    wire N__73279;
    wire N__73276;
    wire N__73275;
    wire N__73272;
    wire N__73269;
    wire N__73266;
    wire N__73261;
    wire N__73258;
    wire N__73255;
    wire N__73252;
    wire N__73249;
    wire N__73246;
    wire N__73243;
    wire N__73240;
    wire N__73237;
    wire N__73234;
    wire N__73231;
    wire N__73230;
    wire N__73227;
    wire N__73224;
    wire N__73219;
    wire N__73216;
    wire N__73213;
    wire N__73210;
    wire N__73207;
    wire N__73204;
    wire N__73201;
    wire N__73198;
    wire N__73195;
    wire N__73192;
    wire N__73189;
    wire N__73186;
    wire N__73183;
    wire N__73180;
    wire N__73177;
    wire N__73176;
    wire N__73175;
    wire N__73172;
    wire N__73167;
    wire N__73164;
    wire N__73161;
    wire N__73156;
    wire N__73153;
    wire N__73152;
    wire N__73149;
    wire N__73146;
    wire N__73143;
    wire N__73140;
    wire N__73137;
    wire N__73134;
    wire N__73131;
    wire N__73128;
    wire N__73123;
    wire N__73122;
    wire N__73117;
    wire N__73114;
    wire N__73111;
    wire N__73108;
    wire N__73105;
    wire N__73102;
    wire N__73099;
    wire N__73098;
    wire N__73097;
    wire N__73096;
    wire N__73093;
    wire N__73090;
    wire N__73085;
    wire N__73078;
    wire N__73077;
    wire N__73074;
    wire N__73073;
    wire N__73070;
    wire N__73065;
    wire N__73064;
    wire N__73059;
    wire N__73056;
    wire N__73051;
    wire N__73048;
    wire N__73045;
    wire N__73042;
    wire N__73039;
    wire N__73036;
    wire N__73033;
    wire N__73032;
    wire N__73031;
    wire N__73030;
    wire N__73029;
    wire N__73026;
    wire N__73025;
    wire N__73020;
    wire N__73011;
    wire N__73006;
    wire N__73003;
    wire N__73000;
    wire N__72997;
    wire N__72994;
    wire N__72991;
    wire N__72990;
    wire N__72989;
    wire N__72986;
    wire N__72983;
    wire N__72978;
    wire N__72973;
    wire N__72970;
    wire N__72967;
    wire N__72964;
    wire N__72963;
    wire N__72960;
    wire N__72957;
    wire N__72952;
    wire N__72951;
    wire N__72950;
    wire N__72949;
    wire N__72948;
    wire N__72947;
    wire N__72944;
    wire N__72941;
    wire N__72940;
    wire N__72937;
    wire N__72934;
    wire N__72931;
    wire N__72930;
    wire N__72929;
    wire N__72928;
    wire N__72927;
    wire N__72926;
    wire N__72925;
    wire N__72924;
    wire N__72923;
    wire N__72920;
    wire N__72917;
    wire N__72914;
    wire N__72909;
    wire N__72904;
    wire N__72901;
    wire N__72896;
    wire N__72893;
    wire N__72890;
    wire N__72887;
    wire N__72880;
    wire N__72875;
    wire N__72870;
    wire N__72867;
    wire N__72864;
    wire N__72857;
    wire N__72854;
    wire N__72849;
    wire N__72844;
    wire N__72835;
    wire N__72832;
    wire N__72831;
    wire N__72830;
    wire N__72825;
    wire N__72822;
    wire N__72819;
    wire N__72814;
    wire N__72811;
    wire N__72810;
    wire N__72807;
    wire N__72804;
    wire N__72801;
    wire N__72798;
    wire N__72795;
    wire N__72790;
    wire N__72787;
    wire N__72784;
    wire N__72781;
    wire N__72778;
    wire N__72775;
    wire N__72772;
    wire N__72771;
    wire N__72768;
    wire N__72765;
    wire N__72762;
    wire N__72757;
    wire N__72756;
    wire N__72751;
    wire N__72750;
    wire N__72749;
    wire N__72748;
    wire N__72745;
    wire N__72738;
    wire N__72733;
    wire N__72730;
    wire N__72727;
    wire N__72726;
    wire N__72723;
    wire N__72720;
    wire N__72715;
    wire N__72712;
    wire N__72709;
    wire N__72706;
    wire N__72703;
    wire N__72702;
    wire N__72699;
    wire N__72696;
    wire N__72693;
    wire N__72690;
    wire N__72685;
    wire N__72682;
    wire N__72679;
    wire N__72676;
    wire N__72673;
    wire N__72670;
    wire N__72667;
    wire N__72664;
    wire N__72661;
    wire N__72660;
    wire N__72659;
    wire N__72656;
    wire N__72653;
    wire N__72650;
    wire N__72647;
    wire N__72640;
    wire N__72637;
    wire N__72634;
    wire N__72631;
    wire N__72630;
    wire N__72629;
    wire N__72626;
    wire N__72621;
    wire N__72616;
    wire N__72615;
    wire N__72612;
    wire N__72609;
    wire N__72604;
    wire N__72603;
    wire N__72600;
    wire N__72597;
    wire N__72594;
    wire N__72589;
    wire N__72586;
    wire N__72585;
    wire N__72580;
    wire N__72579;
    wire N__72576;
    wire N__72573;
    wire N__72568;
    wire N__72567;
    wire N__72566;
    wire N__72565;
    wire N__72562;
    wire N__72559;
    wire N__72556;
    wire N__72553;
    wire N__72550;
    wire N__72547;
    wire N__72544;
    wire N__72541;
    wire N__72536;
    wire N__72529;
    wire N__72526;
    wire N__72525;
    wire N__72524;
    wire N__72521;
    wire N__72518;
    wire N__72515;
    wire N__72512;
    wire N__72505;
    wire N__72502;
    wire N__72499;
    wire N__72496;
    wire N__72493;
    wire N__72490;
    wire N__72489;
    wire N__72484;
    wire N__72481;
    wire N__72478;
    wire N__72475;
    wire N__72474;
    wire N__72469;
    wire N__72468;
    wire N__72465;
    wire N__72462;
    wire N__72457;
    wire N__72454;
    wire N__72451;
    wire N__72448;
    wire N__72445;
    wire N__72442;
    wire N__72441;
    wire N__72438;
    wire N__72435;
    wire N__72432;
    wire N__72429;
    wire N__72424;
    wire N__72421;
    wire N__72418;
    wire N__72415;
    wire N__72412;
    wire N__72409;
    wire N__72408;
    wire N__72407;
    wire N__72402;
    wire N__72399;
    wire N__72396;
    wire N__72393;
    wire N__72390;
    wire N__72385;
    wire N__72382;
    wire N__72379;
    wire N__72376;
    wire N__72375;
    wire N__72370;
    wire N__72367;
    wire N__72364;
    wire N__72361;
    wire N__72358;
    wire N__72355;
    wire N__72352;
    wire N__72351;
    wire N__72348;
    wire N__72345;
    wire N__72340;
    wire N__72337;
    wire N__72336;
    wire N__72333;
    wire N__72330;
    wire N__72329;
    wire N__72326;
    wire N__72323;
    wire N__72320;
    wire N__72315;
    wire N__72310;
    wire N__72307;
    wire N__72304;
    wire N__72301;
    wire N__72298;
    wire N__72295;
    wire N__72292;
    wire N__72289;
    wire N__72286;
    wire N__72285;
    wire N__72280;
    wire N__72277;
    wire N__72274;
    wire N__72273;
    wire N__72272;
    wire N__72267;
    wire N__72264;
    wire N__72261;
    wire N__72256;
    wire N__72253;
    wire N__72250;
    wire N__72247;
    wire N__72244;
    wire N__72241;
    wire N__72240;
    wire N__72239;
    wire N__72238;
    wire N__72231;
    wire N__72228;
    wire N__72223;
    wire N__72220;
    wire N__72217;
    wire N__72216;
    wire N__72213;
    wire N__72210;
    wire N__72207;
    wire N__72202;
    wire N__72199;
    wire N__72198;
    wire N__72195;
    wire N__72192;
    wire N__72191;
    wire N__72188;
    wire N__72185;
    wire N__72182;
    wire N__72179;
    wire N__72174;
    wire N__72171;
    wire N__72168;
    wire N__72163;
    wire N__72160;
    wire N__72157;
    wire N__72154;
    wire N__72151;
    wire N__72148;
    wire N__72145;
    wire N__72142;
    wire N__72139;
    wire N__72136;
    wire N__72133;
    wire N__72132;
    wire N__72131;
    wire N__72128;
    wire N__72125;
    wire N__72122;
    wire N__72119;
    wire N__72116;
    wire N__72113;
    wire N__72106;
    wire N__72105;
    wire N__72102;
    wire N__72099;
    wire N__72094;
    wire N__72091;
    wire N__72088;
    wire N__72085;
    wire N__72084;
    wire N__72081;
    wire N__72078;
    wire N__72075;
    wire N__72072;
    wire N__72069;
    wire N__72066;
    wire N__72061;
    wire N__72058;
    wire N__72057;
    wire N__72056;
    wire N__72053;
    wire N__72048;
    wire N__72045;
    wire N__72042;
    wire N__72037;
    wire N__72034;
    wire N__72033;
    wire N__72030;
    wire N__72027;
    wire N__72024;
    wire N__72021;
    wire N__72016;
    wire N__72013;
    wire N__72012;
    wire N__72009;
    wire N__72006;
    wire N__72003;
    wire N__72000;
    wire N__71995;
    wire N__71992;
    wire N__71989;
    wire N__71986;
    wire N__71983;
    wire N__71980;
    wire N__71977;
    wire N__71974;
    wire N__71971;
    wire N__71970;
    wire N__71969;
    wire N__71968;
    wire N__71965;
    wire N__71960;
    wire N__71957;
    wire N__71950;
    wire N__71947;
    wire N__71946;
    wire N__71945;
    wire N__71940;
    wire N__71939;
    wire N__71936;
    wire N__71935;
    wire N__71932;
    wire N__71929;
    wire N__71924;
    wire N__71917;
    wire N__71914;
    wire N__71913;
    wire N__71912;
    wire N__71909;
    wire N__71906;
    wire N__71905;
    wire N__71904;
    wire N__71903;
    wire N__71902;
    wire N__71899;
    wire N__71892;
    wire N__71889;
    wire N__71886;
    wire N__71881;
    wire N__71878;
    wire N__71869;
    wire N__71866;
    wire N__71863;
    wire N__71860;
    wire N__71857;
    wire N__71854;
    wire N__71853;
    wire N__71848;
    wire N__71845;
    wire N__71844;
    wire N__71843;
    wire N__71842;
    wire N__71839;
    wire N__71836;
    wire N__71831;
    wire N__71824;
    wire N__71821;
    wire N__71818;
    wire N__71817;
    wire N__71816;
    wire N__71813;
    wire N__71810;
    wire N__71809;
    wire N__71806;
    wire N__71805;
    wire N__71804;
    wire N__71799;
    wire N__71796;
    wire N__71795;
    wire N__71794;
    wire N__71791;
    wire N__71788;
    wire N__71787;
    wire N__71786;
    wire N__71785;
    wire N__71782;
    wire N__71777;
    wire N__71774;
    wire N__71771;
    wire N__71766;
    wire N__71763;
    wire N__71760;
    wire N__71757;
    wire N__71748;
    wire N__71747;
    wire N__71742;
    wire N__71739;
    wire N__71734;
    wire N__71731;
    wire N__71726;
    wire N__71721;
    wire N__71716;
    wire N__71715;
    wire N__71714;
    wire N__71711;
    wire N__71708;
    wire N__71707;
    wire N__71706;
    wire N__71705;
    wire N__71704;
    wire N__71701;
    wire N__71700;
    wire N__71699;
    wire N__71696;
    wire N__71693;
    wire N__71690;
    wire N__71687;
    wire N__71684;
    wire N__71683;
    wire N__71680;
    wire N__71677;
    wire N__71674;
    wire N__71671;
    wire N__71668;
    wire N__71661;
    wire N__71658;
    wire N__71655;
    wire N__71652;
    wire N__71645;
    wire N__71640;
    wire N__71635;
    wire N__71630;
    wire N__71629;
    wire N__71628;
    wire N__71627;
    wire N__71624;
    wire N__71621;
    wire N__71618;
    wire N__71615;
    wire N__71612;
    wire N__71609;
    wire N__71596;
    wire N__71595;
    wire N__71592;
    wire N__71589;
    wire N__71586;
    wire N__71583;
    wire N__71580;
    wire N__71577;
    wire N__71574;
    wire N__71571;
    wire N__71566;
    wire N__71563;
    wire N__71562;
    wire N__71559;
    wire N__71556;
    wire N__71553;
    wire N__71552;
    wire N__71549;
    wire N__71546;
    wire N__71543;
    wire N__71540;
    wire N__71535;
    wire N__71530;
    wire N__71527;
    wire N__71524;
    wire N__71521;
    wire N__71518;
    wire N__71515;
    wire N__71512;
    wire N__71509;
    wire N__71506;
    wire N__71503;
    wire N__71500;
    wire N__71497;
    wire N__71494;
    wire N__71491;
    wire N__71488;
    wire N__71485;
    wire N__71482;
    wire N__71479;
    wire N__71476;
    wire N__71473;
    wire N__71470;
    wire N__71467;
    wire N__71464;
    wire N__71461;
    wire N__71458;
    wire N__71455;
    wire N__71452;
    wire N__71449;
    wire N__71448;
    wire N__71443;
    wire N__71440;
    wire N__71437;
    wire N__71434;
    wire N__71433;
    wire N__71432;
    wire N__71429;
    wire N__71424;
    wire N__71421;
    wire N__71418;
    wire N__71415;
    wire N__71412;
    wire N__71407;
    wire N__71406;
    wire N__71401;
    wire N__71398;
    wire N__71397;
    wire N__71394;
    wire N__71391;
    wire N__71390;
    wire N__71387;
    wire N__71384;
    wire N__71381;
    wire N__71376;
    wire N__71371;
    wire N__71370;
    wire N__71365;
    wire N__71362;
    wire N__71361;
    wire N__71360;
    wire N__71359;
    wire N__71354;
    wire N__71349;
    wire N__71344;
    wire N__71341;
    wire N__71338;
    wire N__71337;
    wire N__71336;
    wire N__71333;
    wire N__71328;
    wire N__71325;
    wire N__71320;
    wire N__71317;
    wire N__71316;
    wire N__71311;
    wire N__71308;
    wire N__71305;
    wire N__71302;
    wire N__71299;
    wire N__71296;
    wire N__71293;
    wire N__71290;
    wire N__71287;
    wire N__71286;
    wire N__71283;
    wire N__71280;
    wire N__71277;
    wire N__71274;
    wire N__71271;
    wire N__71266;
    wire N__71265;
    wire N__71260;
    wire N__71257;
    wire N__71256;
    wire N__71255;
    wire N__71252;
    wire N__71247;
    wire N__71244;
    wire N__71241;
    wire N__71236;
    wire N__71233;
    wire N__71232;
    wire N__71227;
    wire N__71224;
    wire N__71223;
    wire N__71220;
    wire N__71219;
    wire N__71216;
    wire N__71213;
    wire N__71210;
    wire N__71207;
    wire N__71202;
    wire N__71197;
    wire N__71194;
    wire N__71193;
    wire N__71188;
    wire N__71185;
    wire N__71184;
    wire N__71183;
    wire N__71180;
    wire N__71175;
    wire N__71172;
    wire N__71169;
    wire N__71164;
    wire N__71161;
    wire N__71160;
    wire N__71157;
    wire N__71154;
    wire N__71149;
    wire N__71146;
    wire N__71143;
    wire N__71142;
    wire N__71139;
    wire N__71136;
    wire N__71131;
    wire N__71128;
    wire N__71127;
    wire N__71124;
    wire N__71121;
    wire N__71116;
    wire N__71115;
    wire N__71114;
    wire N__71111;
    wire N__71106;
    wire N__71103;
    wire N__71100;
    wire N__71095;
    wire N__71092;
    wire N__71091;
    wire N__71088;
    wire N__71085;
    wire N__71082;
    wire N__71079;
    wire N__71076;
    wire N__71073;
    wire N__71068;
    wire N__71065;
    wire N__71064;
    wire N__71063;
    wire N__71062;
    wire N__71061;
    wire N__71058;
    wire N__71057;
    wire N__71052;
    wire N__71051;
    wire N__71048;
    wire N__71047;
    wire N__71046;
    wire N__71045;
    wire N__71044;
    wire N__71041;
    wire N__71040;
    wire N__71039;
    wire N__71038;
    wire N__71037;
    wire N__71034;
    wire N__71031;
    wire N__71030;
    wire N__71029;
    wire N__71028;
    wire N__71027;
    wire N__71026;
    wire N__71025;
    wire N__71024;
    wire N__71023;
    wire N__71022;
    wire N__71019;
    wire N__71018;
    wire N__71017;
    wire N__71008;
    wire N__71005;
    wire N__70998;
    wire N__70993;
    wire N__70990;
    wire N__70985;
    wire N__70984;
    wire N__70983;
    wire N__70982;
    wire N__70981;
    wire N__70980;
    wire N__70979;
    wire N__70978;
    wire N__70977;
    wire N__70974;
    wire N__70973;
    wire N__70972;
    wire N__70967;
    wire N__70966;
    wire N__70965;
    wire N__70964;
    wire N__70963;
    wire N__70962;
    wire N__70961;
    wire N__70960;
    wire N__70955;
    wire N__70948;
    wire N__70945;
    wire N__70942;
    wire N__70939;
    wire N__70938;
    wire N__70935;
    wire N__70930;
    wire N__70929;
    wire N__70926;
    wire N__70919;
    wire N__70918;
    wire N__70911;
    wire N__70906;
    wire N__70899;
    wire N__70896;
    wire N__70893;
    wire N__70890;
    wire N__70887;
    wire N__70884;
    wire N__70881;
    wire N__70880;
    wire N__70875;
    wire N__70870;
    wire N__70867;
    wire N__70864;
    wire N__70861;
    wire N__70858;
    wire N__70855;
    wire N__70852;
    wire N__70851;
    wire N__70850;
    wire N__70847;
    wire N__70844;
    wire N__70843;
    wire N__70840;
    wire N__70839;
    wire N__70838;
    wire N__70835;
    wire N__70830;
    wire N__70827;
    wire N__70820;
    wire N__70817;
    wire N__70812;
    wire N__70811;
    wire N__70810;
    wire N__70807;
    wire N__70806;
    wire N__70805;
    wire N__70804;
    wire N__70803;
    wire N__70802;
    wire N__70797;
    wire N__70796;
    wire N__70795;
    wire N__70794;
    wire N__70791;
    wire N__70788;
    wire N__70781;
    wire N__70776;
    wire N__70771;
    wire N__70766;
    wire N__70763;
    wire N__70760;
    wire N__70757;
    wire N__70754;
    wire N__70753;
    wire N__70750;
    wire N__70747;
    wire N__70740;
    wire N__70737;
    wire N__70732;
    wire N__70731;
    wire N__70730;
    wire N__70729;
    wire N__70724;
    wire N__70721;
    wire N__70716;
    wire N__70709;
    wire N__70706;
    wire N__70705;
    wire N__70704;
    wire N__70697;
    wire N__70688;
    wire N__70683;
    wire N__70674;
    wire N__70671;
    wire N__70666;
    wire N__70659;
    wire N__70652;
    wire N__70641;
    wire N__70636;
    wire N__70627;
    wire N__70612;
    wire N__70611;
    wire N__70610;
    wire N__70607;
    wire N__70606;
    wire N__70605;
    wire N__70604;
    wire N__70601;
    wire N__70596;
    wire N__70593;
    wire N__70590;
    wire N__70587;
    wire N__70584;
    wire N__70581;
    wire N__70578;
    wire N__70575;
    wire N__70572;
    wire N__70569;
    wire N__70566;
    wire N__70563;
    wire N__70560;
    wire N__70559;
    wire N__70558;
    wire N__70557;
    wire N__70554;
    wire N__70551;
    wire N__70544;
    wire N__70537;
    wire N__70534;
    wire N__70525;
    wire N__70522;
    wire N__70521;
    wire N__70520;
    wire N__70519;
    wire N__70518;
    wire N__70517;
    wire N__70516;
    wire N__70515;
    wire N__70502;
    wire N__70499;
    wire N__70498;
    wire N__70497;
    wire N__70496;
    wire N__70495;
    wire N__70492;
    wire N__70489;
    wire N__70486;
    wire N__70483;
    wire N__70482;
    wire N__70479;
    wire N__70476;
    wire N__70473;
    wire N__70470;
    wire N__70469;
    wire N__70462;
    wire N__70461;
    wire N__70458;
    wire N__70451;
    wire N__70448;
    wire N__70447;
    wire N__70444;
    wire N__70441;
    wire N__70436;
    wire N__70433;
    wire N__70430;
    wire N__70425;
    wire N__70422;
    wire N__70411;
    wire N__70410;
    wire N__70407;
    wire N__70404;
    wire N__70399;
    wire N__70396;
    wire N__70395;
    wire N__70394;
    wire N__70391;
    wire N__70386;
    wire N__70383;
    wire N__70380;
    wire N__70375;
    wire N__70372;
    wire N__70369;
    wire N__70366;
    wire N__70365;
    wire N__70362;
    wire N__70359;
    wire N__70356;
    wire N__70353;
    wire N__70350;
    wire N__70345;
    wire N__70342;
    wire N__70339;
    wire N__70336;
    wire N__70333;
    wire N__70332;
    wire N__70327;
    wire N__70324;
    wire N__70321;
    wire N__70318;
    wire N__70315;
    wire N__70314;
    wire N__70311;
    wire N__70308;
    wire N__70303;
    wire N__70300;
    wire N__70297;
    wire N__70294;
    wire N__70291;
    wire N__70288;
    wire N__70285;
    wire N__70282;
    wire N__70281;
    wire N__70278;
    wire N__70277;
    wire N__70274;
    wire N__70269;
    wire N__70268;
    wire N__70263;
    wire N__70260;
    wire N__70257;
    wire N__70252;
    wire N__70249;
    wire N__70246;
    wire N__70243;
    wire N__70240;
    wire N__70237;
    wire N__70236;
    wire N__70231;
    wire N__70228;
    wire N__70225;
    wire N__70224;
    wire N__70219;
    wire N__70216;
    wire N__70213;
    wire N__70210;
    wire N__70207;
    wire N__70204;
    wire N__70203;
    wire N__70198;
    wire N__70195;
    wire N__70192;
    wire N__70189;
    wire N__70186;
    wire N__70183;
    wire N__70182;
    wire N__70177;
    wire N__70174;
    wire N__70171;
    wire N__70170;
    wire N__70169;
    wire N__70166;
    wire N__70161;
    wire N__70158;
    wire N__70155;
    wire N__70150;
    wire N__70149;
    wire N__70146;
    wire N__70145;
    wire N__70140;
    wire N__70137;
    wire N__70132;
    wire N__70129;
    wire N__70126;
    wire N__70123;
    wire N__70120;
    wire N__70117;
    wire N__70116;
    wire N__70113;
    wire N__70110;
    wire N__70107;
    wire N__70104;
    wire N__70099;
    wire N__70096;
    wire N__70095;
    wire N__70092;
    wire N__70091;
    wire N__70084;
    wire N__70081;
    wire N__70078;
    wire N__70075;
    wire N__70072;
    wire N__70069;
    wire N__70066;
    wire N__70065;
    wire N__70062;
    wire N__70061;
    wire N__70058;
    wire N__70057;
    wire N__70054;
    wire N__70051;
    wire N__70048;
    wire N__70045;
    wire N__70042;
    wire N__70037;
    wire N__70034;
    wire N__70027;
    wire N__70024;
    wire N__70023;
    wire N__70022;
    wire N__70019;
    wire N__70016;
    wire N__70013;
    wire N__70008;
    wire N__70005;
    wire N__70002;
    wire N__70001;
    wire N__69998;
    wire N__69995;
    wire N__69992;
    wire N__69985;
    wire N__69982;
    wire N__69979;
    wire N__69976;
    wire N__69975;
    wire N__69974;
    wire N__69967;
    wire N__69964;
    wire N__69961;
    wire N__69958;
    wire N__69957;
    wire N__69954;
    wire N__69951;
    wire N__69950;
    wire N__69945;
    wire N__69942;
    wire N__69939;
    wire N__69934;
    wire N__69931;
    wire N__69930;
    wire N__69927;
    wire N__69924;
    wire N__69921;
    wire N__69916;
    wire N__69913;
    wire N__69910;
    wire N__69909;
    wire N__69908;
    wire N__69905;
    wire N__69900;
    wire N__69895;
    wire N__69894;
    wire N__69891;
    wire N__69888;
    wire N__69883;
    wire N__69882;
    wire N__69879;
    wire N__69876;
    wire N__69873;
    wire N__69870;
    wire N__69867;
    wire N__69866;
    wire N__69863;
    wire N__69860;
    wire N__69857;
    wire N__69850;
    wire N__69849;
    wire N__69846;
    wire N__69843;
    wire N__69838;
    wire N__69835;
    wire N__69832;
    wire N__69829;
    wire N__69826;
    wire N__69823;
    wire N__69820;
    wire N__69817;
    wire N__69814;
    wire N__69811;
    wire N__69808;
    wire N__69805;
    wire N__69802;
    wire N__69799;
    wire N__69796;
    wire N__69793;
    wire N__69790;
    wire N__69787;
    wire N__69784;
    wire N__69781;
    wire N__69778;
    wire N__69775;
    wire N__69772;
    wire N__69769;
    wire N__69766;
    wire N__69763;
    wire N__69760;
    wire N__69757;
    wire N__69754;
    wire N__69751;
    wire N__69748;
    wire N__69745;
    wire N__69742;
    wire N__69739;
    wire N__69736;
    wire N__69733;
    wire N__69730;
    wire N__69727;
    wire N__69724;
    wire N__69721;
    wire N__69718;
    wire N__69715;
    wire N__69712;
    wire N__69709;
    wire N__69706;
    wire N__69703;
    wire N__69702;
    wire N__69701;
    wire N__69696;
    wire N__69693;
    wire N__69690;
    wire N__69687;
    wire N__69684;
    wire N__69681;
    wire N__69676;
    wire N__69675;
    wire N__69670;
    wire N__69667;
    wire N__69664;
    wire N__69661;
    wire N__69658;
    wire N__69657;
    wire N__69654;
    wire N__69651;
    wire N__69648;
    wire N__69645;
    wire N__69640;
    wire N__69637;
    wire N__69634;
    wire N__69631;
    wire N__69628;
    wire N__69625;
    wire N__69622;
    wire N__69619;
    wire N__69616;
    wire N__69613;
    wire N__69610;
    wire N__69607;
    wire N__69604;
    wire N__69601;
    wire N__69598;
    wire N__69595;
    wire N__69594;
    wire N__69591;
    wire N__69588;
    wire N__69583;
    wire N__69582;
    wire N__69581;
    wire N__69580;
    wire N__69577;
    wire N__69574;
    wire N__69571;
    wire N__69568;
    wire N__69565;
    wire N__69562;
    wire N__69559;
    wire N__69556;
    wire N__69553;
    wire N__69552;
    wire N__69545;
    wire N__69542;
    wire N__69539;
    wire N__69532;
    wire N__69529;
    wire N__69526;
    wire N__69523;
    wire N__69520;
    wire N__69517;
    wire N__69514;
    wire N__69511;
    wire N__69508;
    wire N__69505;
    wire N__69504;
    wire N__69501;
    wire N__69498;
    wire N__69495;
    wire N__69492;
    wire N__69491;
    wire N__69486;
    wire N__69483;
    wire N__69482;
    wire N__69481;
    wire N__69478;
    wire N__69475;
    wire N__69470;
    wire N__69467;
    wire N__69464;
    wire N__69461;
    wire N__69458;
    wire N__69451;
    wire N__69448;
    wire N__69445;
    wire N__69442;
    wire N__69441;
    wire N__69438;
    wire N__69435;
    wire N__69432;
    wire N__69429;
    wire N__69424;
    wire N__69421;
    wire N__69418;
    wire N__69417;
    wire N__69416;
    wire N__69411;
    wire N__69410;
    wire N__69409;
    wire N__69408;
    wire N__69405;
    wire N__69402;
    wire N__69397;
    wire N__69394;
    wire N__69393;
    wire N__69392;
    wire N__69389;
    wire N__69386;
    wire N__69381;
    wire N__69376;
    wire N__69375;
    wire N__69374;
    wire N__69373;
    wire N__69372;
    wire N__69371;
    wire N__69368;
    wire N__69361;
    wire N__69350;
    wire N__69343;
    wire N__69342;
    wire N__69339;
    wire N__69336;
    wire N__69333;
    wire N__69330;
    wire N__69327;
    wire N__69322;
    wire N__69319;
    wire N__69316;
    wire N__69315;
    wire N__69312;
    wire N__69309;
    wire N__69304;
    wire N__69301;
    wire N__69298;
    wire N__69295;
    wire N__69292;
    wire N__69291;
    wire N__69290;
    wire N__69287;
    wire N__69282;
    wire N__69279;
    wire N__69276;
    wire N__69275;
    wire N__69274;
    wire N__69273;
    wire N__69272;
    wire N__69269;
    wire N__69266;
    wire N__69261;
    wire N__69256;
    wire N__69247;
    wire N__69246;
    wire N__69243;
    wire N__69240;
    wire N__69237;
    wire N__69234;
    wire N__69231;
    wire N__69228;
    wire N__69223;
    wire N__69222;
    wire N__69219;
    wire N__69216;
    wire N__69213;
    wire N__69210;
    wire N__69207;
    wire N__69202;
    wire N__69199;
    wire N__69198;
    wire N__69195;
    wire N__69192;
    wire N__69191;
    wire N__69190;
    wire N__69187;
    wire N__69184;
    wire N__69183;
    wire N__69182;
    wire N__69179;
    wire N__69178;
    wire N__69177;
    wire N__69174;
    wire N__69171;
    wire N__69168;
    wire N__69165;
    wire N__69162;
    wire N__69159;
    wire N__69156;
    wire N__69151;
    wire N__69150;
    wire N__69147;
    wire N__69142;
    wire N__69139;
    wire N__69132;
    wire N__69129;
    wire N__69124;
    wire N__69121;
    wire N__69118;
    wire N__69115;
    wire N__69112;
    wire N__69109;
    wire N__69106;
    wire N__69105;
    wire N__69104;
    wire N__69101;
    wire N__69098;
    wire N__69093;
    wire N__69088;
    wire N__69079;
    wire N__69078;
    wire N__69077;
    wire N__69074;
    wire N__69071;
    wire N__69068;
    wire N__69065;
    wire N__69062;
    wire N__69059;
    wire N__69056;
    wire N__69053;
    wire N__69050;
    wire N__69047;
    wire N__69046;
    wire N__69045;
    wire N__69038;
    wire N__69033;
    wire N__69030;
    wire N__69025;
    wire N__69024;
    wire N__69023;
    wire N__69022;
    wire N__69021;
    wire N__69020;
    wire N__69019;
    wire N__69018;
    wire N__69015;
    wire N__69014;
    wire N__69013;
    wire N__69012;
    wire N__69011;
    wire N__69010;
    wire N__69009;
    wire N__69008;
    wire N__69005;
    wire N__69004;
    wire N__69003;
    wire N__69002;
    wire N__68985;
    wire N__68980;
    wire N__68979;
    wire N__68976;
    wire N__68961;
    wire N__68960;
    wire N__68959;
    wire N__68958;
    wire N__68955;
    wire N__68952;
    wire N__68949;
    wire N__68946;
    wire N__68943;
    wire N__68936;
    wire N__68931;
    wire N__68928;
    wire N__68921;
    wire N__68916;
    wire N__68913;
    wire N__68912;
    wire N__68907;
    wire N__68904;
    wire N__68901;
    wire N__68896;
    wire N__68893;
    wire N__68890;
    wire N__68887;
    wire N__68884;
    wire N__68881;
    wire N__68878;
    wire N__68875;
    wire N__68872;
    wire N__68869;
    wire N__68866;
    wire N__68863;
    wire N__68860;
    wire N__68857;
    wire N__68854;
    wire N__68851;
    wire N__68848;
    wire N__68845;
    wire N__68842;
    wire N__68839;
    wire N__68836;
    wire N__68833;
    wire N__68830;
    wire N__68827;
    wire N__68824;
    wire N__68821;
    wire N__68818;
    wire N__68815;
    wire N__68812;
    wire N__68809;
    wire N__68806;
    wire N__68803;
    wire N__68800;
    wire N__68797;
    wire N__68794;
    wire N__68791;
    wire N__68788;
    wire N__68785;
    wire N__68782;
    wire N__68779;
    wire N__68776;
    wire N__68773;
    wire N__68770;
    wire N__68767;
    wire N__68764;
    wire N__68761;
    wire N__68758;
    wire N__68755;
    wire N__68752;
    wire N__68749;
    wire N__68746;
    wire N__68745;
    wire N__68742;
    wire N__68739;
    wire N__68734;
    wire N__68731;
    wire N__68728;
    wire N__68725;
    wire N__68722;
    wire N__68719;
    wire N__68716;
    wire N__68713;
    wire N__68712;
    wire N__68709;
    wire N__68706;
    wire N__68703;
    wire N__68700;
    wire N__68699;
    wire N__68696;
    wire N__68693;
    wire N__68690;
    wire N__68683;
    wire N__68680;
    wire N__68677;
    wire N__68674;
    wire N__68671;
    wire N__68670;
    wire N__68667;
    wire N__68664;
    wire N__68661;
    wire N__68658;
    wire N__68655;
    wire N__68650;
    wire N__68649;
    wire N__68646;
    wire N__68643;
    wire N__68640;
    wire N__68637;
    wire N__68634;
    wire N__68629;
    wire N__68626;
    wire N__68623;
    wire N__68622;
    wire N__68619;
    wire N__68616;
    wire N__68611;
    wire N__68608;
    wire N__68605;
    wire N__68602;
    wire N__68599;
    wire N__68596;
    wire N__68593;
    wire N__68590;
    wire N__68589;
    wire N__68588;
    wire N__68585;
    wire N__68580;
    wire N__68577;
    wire N__68574;
    wire N__68569;
    wire N__68566;
    wire N__68563;
    wire N__68562;
    wire N__68561;
    wire N__68558;
    wire N__68553;
    wire N__68548;
    wire N__68545;
    wire N__68542;
    wire N__68539;
    wire N__68538;
    wire N__68535;
    wire N__68532;
    wire N__68529;
    wire N__68524;
    wire N__68521;
    wire N__68518;
    wire N__68517;
    wire N__68512;
    wire N__68509;
    wire N__68506;
    wire N__68503;
    wire N__68502;
    wire N__68499;
    wire N__68498;
    wire N__68491;
    wire N__68488;
    wire N__68485;
    wire N__68484;
    wire N__68481;
    wire N__68478;
    wire N__68475;
    wire N__68470;
    wire N__68467;
    wire N__68464;
    wire N__68461;
    wire N__68458;
    wire N__68455;
    wire N__68452;
    wire N__68449;
    wire N__68446;
    wire N__68443;
    wire N__68440;
    wire N__68437;
    wire N__68436;
    wire N__68433;
    wire N__68430;
    wire N__68425;
    wire N__68422;
    wire N__68419;
    wire N__68416;
    wire N__68413;
    wire N__68410;
    wire N__68407;
    wire N__68404;
    wire N__68401;
    wire N__68398;
    wire N__68395;
    wire N__68392;
    wire N__68389;
    wire N__68386;
    wire N__68383;
    wire N__68380;
    wire N__68377;
    wire N__68374;
    wire N__68371;
    wire N__68370;
    wire N__68369;
    wire N__68366;
    wire N__68361;
    wire N__68358;
    wire N__68355;
    wire N__68350;
    wire N__68347;
    wire N__68344;
    wire N__68341;
    wire N__68340;
    wire N__68337;
    wire N__68334;
    wire N__68329;
    wire N__68326;
    wire N__68323;
    wire N__68320;
    wire N__68319;
    wire N__68318;
    wire N__68315;
    wire N__68310;
    wire N__68305;
    wire N__68302;
    wire N__68299;
    wire N__68296;
    wire N__68293;
    wire N__68292;
    wire N__68289;
    wire N__68286;
    wire N__68281;
    wire N__68280;
    wire N__68279;
    wire N__68276;
    wire N__68271;
    wire N__68266;
    wire N__68263;
    wire N__68260;
    wire N__68257;
    wire N__68254;
    wire N__68253;
    wire N__68252;
    wire N__68249;
    wire N__68246;
    wire N__68243;
    wire N__68240;
    wire N__68235;
    wire N__68232;
    wire N__68229;
    wire N__68224;
    wire N__68221;
    wire N__68218;
    wire N__68217;
    wire N__68214;
    wire N__68211;
    wire N__68206;
    wire N__68203;
    wire N__68200;
    wire N__68197;
    wire N__68196;
    wire N__68193;
    wire N__68190;
    wire N__68185;
    wire N__68182;
    wire N__68179;
    wire N__68176;
    wire N__68175;
    wire N__68170;
    wire N__68169;
    wire N__68166;
    wire N__68163;
    wire N__68160;
    wire N__68155;
    wire N__68154;
    wire N__68151;
    wire N__68148;
    wire N__68143;
    wire N__68142;
    wire N__68141;
    wire N__68138;
    wire N__68133;
    wire N__68128;
    wire N__68125;
    wire N__68122;
    wire N__68119;
    wire N__68118;
    wire N__68113;
    wire N__68110;
    wire N__68107;
    wire N__68104;
    wire N__68101;
    wire N__68100;
    wire N__68097;
    wire N__68094;
    wire N__68089;
    wire N__68086;
    wire N__68085;
    wire N__68084;
    wire N__68079;
    wire N__68076;
    wire N__68071;
    wire N__68068;
    wire N__68065;
    wire N__68064;
    wire N__68063;
    wire N__68060;
    wire N__68057;
    wire N__68054;
    wire N__68047;
    wire N__68044;
    wire N__68041;
    wire N__68040;
    wire N__68037;
    wire N__68036;
    wire N__68033;
    wire N__68028;
    wire N__68025;
    wire N__68022;
    wire N__68017;
    wire N__68014;
    wire N__68011;
    wire N__68008;
    wire N__68005;
    wire N__68002;
    wire N__67999;
    wire N__67996;
    wire N__67993;
    wire N__67990;
    wire N__67989;
    wire N__67986;
    wire N__67983;
    wire N__67980;
    wire N__67979;
    wire N__67976;
    wire N__67973;
    wire N__67970;
    wire N__67967;
    wire N__67960;
    wire N__67957;
    wire N__67956;
    wire N__67953;
    wire N__67950;
    wire N__67945;
    wire N__67944;
    wire N__67943;
    wire N__67940;
    wire N__67935;
    wire N__67930;
    wire N__67929;
    wire N__67924;
    wire N__67921;
    wire N__67918;
    wire N__67917;
    wire N__67916;
    wire N__67913;
    wire N__67908;
    wire N__67903;
    wire N__67900;
    wire N__67897;
    wire N__67894;
    wire N__67891;
    wire N__67890;
    wire N__67887;
    wire N__67884;
    wire N__67881;
    wire N__67880;
    wire N__67877;
    wire N__67874;
    wire N__67871;
    wire N__67864;
    wire N__67861;
    wire N__67858;
    wire N__67855;
    wire N__67852;
    wire N__67851;
    wire N__67850;
    wire N__67847;
    wire N__67842;
    wire N__67839;
    wire N__67836;
    wire N__67833;
    wire N__67830;
    wire N__67825;
    wire N__67822;
    wire N__67819;
    wire N__67816;
    wire N__67813;
    wire N__67810;
    wire N__67809;
    wire N__67806;
    wire N__67803;
    wire N__67800;
    wire N__67795;
    wire N__67792;
    wire N__67791;
    wire N__67786;
    wire N__67783;
    wire N__67782;
    wire N__67777;
    wire N__67774;
    wire N__67771;
    wire N__67770;
    wire N__67767;
    wire N__67764;
    wire N__67759;
    wire N__67756;
    wire N__67753;
    wire N__67750;
    wire N__67749;
    wire N__67746;
    wire N__67743;
    wire N__67740;
    wire N__67735;
    wire N__67732;
    wire N__67729;
    wire N__67726;
    wire N__67723;
    wire N__67720;
    wire N__67717;
    wire N__67716;
    wire N__67711;
    wire N__67708;
    wire N__67705;
    wire N__67702;
    wire N__67699;
    wire N__67698;
    wire N__67693;
    wire N__67692;
    wire N__67689;
    wire N__67688;
    wire N__67687;
    wire N__67686;
    wire N__67685;
    wire N__67684;
    wire N__67681;
    wire N__67678;
    wire N__67675;
    wire N__67672;
    wire N__67669;
    wire N__67664;
    wire N__67659;
    wire N__67648;
    wire N__67647;
    wire N__67642;
    wire N__67641;
    wire N__67640;
    wire N__67639;
    wire N__67636;
    wire N__67635;
    wire N__67634;
    wire N__67633;
    wire N__67630;
    wire N__67627;
    wire N__67624;
    wire N__67621;
    wire N__67616;
    wire N__67613;
    wire N__67600;
    wire N__67599;
    wire N__67596;
    wire N__67593;
    wire N__67588;
    wire N__67587;
    wire N__67584;
    wire N__67583;
    wire N__67580;
    wire N__67579;
    wire N__67574;
    wire N__67571;
    wire N__67568;
    wire N__67565;
    wire N__67558;
    wire N__67557;
    wire N__67554;
    wire N__67551;
    wire N__67546;
    wire N__67545;
    wire N__67544;
    wire N__67541;
    wire N__67536;
    wire N__67531;
    wire N__67528;
    wire N__67525;
    wire N__67522;
    wire N__67519;
    wire N__67516;
    wire N__67513;
    wire N__67510;
    wire N__67509;
    wire N__67506;
    wire N__67503;
    wire N__67498;
    wire N__67495;
    wire N__67492;
    wire N__67491;
    wire N__67486;
    wire N__67483;
    wire N__67482;
    wire N__67477;
    wire N__67474;
    wire N__67471;
    wire N__67468;
    wire N__67467;
    wire N__67466;
    wire N__67465;
    wire N__67460;
    wire N__67455;
    wire N__67450;
    wire N__67449;
    wire N__67448;
    wire N__67447;
    wire N__67442;
    wire N__67437;
    wire N__67432;
    wire N__67429;
    wire N__67428;
    wire N__67427;
    wire N__67426;
    wire N__67423;
    wire N__67418;
    wire N__67415;
    wire N__67408;
    wire N__67405;
    wire N__67402;
    wire N__67399;
    wire N__67396;
    wire N__67393;
    wire N__67390;
    wire N__67389;
    wire N__67386;
    wire N__67383;
    wire N__67380;
    wire N__67377;
    wire N__67372;
    wire N__67369;
    wire N__67366;
    wire N__67363;
    wire N__67360;
    wire N__67357;
    wire N__67354;
    wire N__67351;
    wire N__67348;
    wire N__67345;
    wire N__67342;
    wire N__67339;
    wire N__67336;
    wire N__67333;
    wire N__67330;
    wire N__67327;
    wire N__67324;
    wire N__67321;
    wire N__67318;
    wire N__67315;
    wire N__67312;
    wire N__67309;
    wire N__67306;
    wire N__67303;
    wire N__67300;
    wire N__67297;
    wire N__67294;
    wire N__67291;
    wire N__67288;
    wire N__67285;
    wire N__67284;
    wire N__67279;
    wire N__67276;
    wire N__67273;
    wire N__67270;
    wire N__67269;
    wire N__67264;
    wire N__67261;
    wire N__67258;
    wire N__67255;
    wire N__67252;
    wire N__67249;
    wire N__67248;
    wire N__67247;
    wire N__67240;
    wire N__67237;
    wire N__67234;
    wire N__67231;
    wire N__67228;
    wire N__67225;
    wire N__67222;
    wire N__67221;
    wire N__67218;
    wire N__67215;
    wire N__67210;
    wire N__67209;
    wire N__67206;
    wire N__67203;
    wire N__67198;
    wire N__67195;
    wire N__67194;
    wire N__67191;
    wire N__67188;
    wire N__67183;
    wire N__67180;
    wire N__67177;
    wire N__67174;
    wire N__67171;
    wire N__67168;
    wire N__67165;
    wire N__67162;
    wire N__67159;
    wire N__67156;
    wire N__67155;
    wire N__67150;
    wire N__67147;
    wire N__67144;
    wire N__67143;
    wire N__67138;
    wire N__67135;
    wire N__67134;
    wire N__67129;
    wire N__67126;
    wire N__67123;
    wire N__67120;
    wire N__67117;
    wire N__67114;
    wire N__67113;
    wire N__67108;
    wire N__67105;
    wire N__67102;
    wire N__67099;
    wire N__67098;
    wire N__67097;
    wire N__67094;
    wire N__67093;
    wire N__67092;
    wire N__67091;
    wire N__67090;
    wire N__67089;
    wire N__67088;
    wire N__67085;
    wire N__67082;
    wire N__67079;
    wire N__67078;
    wire N__67075;
    wire N__67072;
    wire N__67071;
    wire N__67070;
    wire N__67063;
    wire N__67060;
    wire N__67055;
    wire N__67052;
    wire N__67045;
    wire N__67044;
    wire N__67043;
    wire N__67040;
    wire N__67039;
    wire N__67036;
    wire N__67027;
    wire N__67024;
    wire N__67015;
    wire N__67012;
    wire N__67009;
    wire N__67004;
    wire N__66997;
    wire N__66994;
    wire N__66991;
    wire N__66990;
    wire N__66987;
    wire N__66984;
    wire N__66981;
    wire N__66978;
    wire N__66977;
    wire N__66974;
    wire N__66971;
    wire N__66968;
    wire N__66961;
    wire N__66960;
    wire N__66957;
    wire N__66954;
    wire N__66951;
    wire N__66948;
    wire N__66945;
    wire N__66942;
    wire N__66939;
    wire N__66934;
    wire N__66931;
    wire N__66928;
    wire N__66925;
    wire N__66922;
    wire N__66921;
    wire N__66920;
    wire N__66915;
    wire N__66912;
    wire N__66909;
    wire N__66906;
    wire N__66901;
    wire N__66898;
    wire N__66897;
    wire N__66896;
    wire N__66889;
    wire N__66886;
    wire N__66883;
    wire N__66880;
    wire N__66877;
    wire N__66874;
    wire N__66871;
    wire N__66868;
    wire N__66865;
    wire N__66862;
    wire N__66859;
    wire N__66856;
    wire N__66853;
    wire N__66850;
    wire N__66847;
    wire N__66844;
    wire N__66841;
    wire N__66838;
    wire N__66835;
    wire N__66834;
    wire N__66833;
    wire N__66830;
    wire N__66825;
    wire N__66820;
    wire N__66819;
    wire N__66816;
    wire N__66815;
    wire N__66812;
    wire N__66807;
    wire N__66804;
    wire N__66799;
    wire N__66798;
    wire N__66795;
    wire N__66792;
    wire N__66787;
    wire N__66784;
    wire N__66781;
    wire N__66778;
    wire N__66777;
    wire N__66774;
    wire N__66771;
    wire N__66766;
    wire N__66763;
    wire N__66760;
    wire N__66757;
    wire N__66756;
    wire N__66753;
    wire N__66750;
    wire N__66745;
    wire N__66742;
    wire N__66741;
    wire N__66740;
    wire N__66739;
    wire N__66738;
    wire N__66733;
    wire N__66726;
    wire N__66721;
    wire N__66718;
    wire N__66715;
    wire N__66712;
    wire N__66709;
    wire N__66708;
    wire N__66707;
    wire N__66706;
    wire N__66705;
    wire N__66704;
    wire N__66703;
    wire N__66696;
    wire N__66695;
    wire N__66694;
    wire N__66693;
    wire N__66692;
    wire N__66691;
    wire N__66684;
    wire N__66681;
    wire N__66678;
    wire N__66669;
    wire N__66668;
    wire N__66667;
    wire N__66664;
    wire N__66663;
    wire N__66662;
    wire N__66661;
    wire N__66658;
    wire N__66651;
    wire N__66644;
    wire N__66641;
    wire N__66636;
    wire N__66631;
    wire N__66622;
    wire N__66621;
    wire N__66618;
    wire N__66615;
    wire N__66612;
    wire N__66609;
    wire N__66606;
    wire N__66603;
    wire N__66598;
    wire N__66595;
    wire N__66592;
    wire N__66589;
    wire N__66586;
    wire N__66583;
    wire N__66580;
    wire N__66577;
    wire N__66574;
    wire N__66571;
    wire N__66568;
    wire N__66565;
    wire N__66562;
    wire N__66559;
    wire N__66558;
    wire N__66557;
    wire N__66556;
    wire N__66555;
    wire N__66552;
    wire N__66545;
    wire N__66542;
    wire N__66539;
    wire N__66532;
    wire N__66529;
    wire N__66526;
    wire N__66525;
    wire N__66520;
    wire N__66517;
    wire N__66514;
    wire N__66511;
    wire N__66510;
    wire N__66505;
    wire N__66502;
    wire N__66499;
    wire N__66496;
    wire N__66493;
    wire N__66490;
    wire N__66487;
    wire N__66484;
    wire N__66481;
    wire N__66478;
    wire N__66475;
    wire N__66472;
    wire N__66471;
    wire N__66466;
    wire N__66463;
    wire N__66460;
    wire N__66457;
    wire N__66454;
    wire N__66451;
    wire N__66448;
    wire N__66445;
    wire N__66442;
    wire N__66439;
    wire N__66436;
    wire N__66433;
    wire N__66430;
    wire N__66427;
    wire N__66424;
    wire N__66421;
    wire N__66418;
    wire N__66415;
    wire N__66412;
    wire N__66409;
    wire N__66406;
    wire N__66403;
    wire N__66400;
    wire N__66397;
    wire N__66394;
    wire N__66391;
    wire N__66388;
    wire N__66385;
    wire N__66382;
    wire N__66379;
    wire N__66376;
    wire N__66373;
    wire N__66370;
    wire N__66367;
    wire N__66366;
    wire N__66363;
    wire N__66360;
    wire N__66355;
    wire N__66352;
    wire N__66349;
    wire N__66346;
    wire N__66343;
    wire N__66340;
    wire N__66337;
    wire N__66334;
    wire N__66333;
    wire N__66332;
    wire N__66329;
    wire N__66326;
    wire N__66323;
    wire N__66316;
    wire N__66313;
    wire N__66310;
    wire N__66307;
    wire N__66304;
    wire N__66301;
    wire N__66298;
    wire N__66295;
    wire N__66292;
    wire N__66289;
    wire N__66286;
    wire N__66283;
    wire N__66282;
    wire N__66279;
    wire N__66276;
    wire N__66273;
    wire N__66270;
    wire N__66265;
    wire N__66264;
    wire N__66261;
    wire N__66258;
    wire N__66255;
    wire N__66252;
    wire N__66249;
    wire N__66246;
    wire N__66241;
    wire N__66238;
    wire N__66235;
    wire N__66232;
    wire N__66229;
    wire N__66226;
    wire N__66223;
    wire N__66220;
    wire N__66217;
    wire N__66216;
    wire N__66213;
    wire N__66210;
    wire N__66209;
    wire N__66204;
    wire N__66201;
    wire N__66196;
    wire N__66193;
    wire N__66190;
    wire N__66187;
    wire N__66184;
    wire N__66181;
    wire N__66178;
    wire N__66175;
    wire N__66172;
    wire N__66169;
    wire N__66166;
    wire N__66163;
    wire N__66160;
    wire N__66157;
    wire N__66156;
    wire N__66151;
    wire N__66148;
    wire N__66145;
    wire N__66142;
    wire N__66139;
    wire N__66136;
    wire N__66133;
    wire N__66130;
    wire N__66127;
    wire N__66124;
    wire N__66121;
    wire N__66118;
    wire N__66115;
    wire N__66112;
    wire N__66109;
    wire N__66106;
    wire N__66103;
    wire N__66100;
    wire N__66097;
    wire N__66094;
    wire N__66091;
    wire N__66088;
    wire N__66085;
    wire N__66082;
    wire N__66079;
    wire N__66076;
    wire N__66073;
    wire N__66072;
    wire N__66071;
    wire N__66068;
    wire N__66065;
    wire N__66064;
    wire N__66061;
    wire N__66058;
    wire N__66055;
    wire N__66052;
    wire N__66047;
    wire N__66042;
    wire N__66039;
    wire N__66036;
    wire N__66031;
    wire N__66028;
    wire N__66025;
    wire N__66022;
    wire N__66019;
    wire N__66016;
    wire N__66013;
    wire N__66010;
    wire N__66007;
    wire N__66004;
    wire N__66001;
    wire N__65998;
    wire N__65995;
    wire N__65992;
    wire N__65989;
    wire N__65986;
    wire N__65983;
    wire N__65980;
    wire N__65977;
    wire N__65974;
    wire N__65971;
    wire N__65968;
    wire N__65965;
    wire N__65962;
    wire N__65959;
    wire N__65956;
    wire N__65955;
    wire N__65954;
    wire N__65953;
    wire N__65950;
    wire N__65949;
    wire N__65948;
    wire N__65945;
    wire N__65942;
    wire N__65941;
    wire N__65938;
    wire N__65937;
    wire N__65936;
    wire N__65933;
    wire N__65930;
    wire N__65927;
    wire N__65924;
    wire N__65921;
    wire N__65918;
    wire N__65917;
    wire N__65914;
    wire N__65911;
    wire N__65908;
    wire N__65907;
    wire N__65904;
    wire N__65901;
    wire N__65898;
    wire N__65895;
    wire N__65890;
    wire N__65887;
    wire N__65882;
    wire N__65879;
    wire N__65878;
    wire N__65875;
    wire N__65874;
    wire N__65869;
    wire N__65868;
    wire N__65867;
    wire N__65866;
    wire N__65865;
    wire N__65864;
    wire N__65863;
    wire N__65862;
    wire N__65861;
    wire N__65860;
    wire N__65859;
    wire N__65858;
    wire N__65855;
    wire N__65854;
    wire N__65851;
    wire N__65846;
    wire N__65845;
    wire N__65842;
    wire N__65839;
    wire N__65836;
    wire N__65833;
    wire N__65830;
    wire N__65829;
    wire N__65826;
    wire N__65823;
    wire N__65822;
    wire N__65819;
    wire N__65816;
    wire N__65813;
    wire N__65810;
    wire N__65807;
    wire N__65804;
    wire N__65801;
    wire N__65798;
    wire N__65795;
    wire N__65794;
    wire N__65793;
    wire N__65792;
    wire N__65789;
    wire N__65788;
    wire N__65785;
    wire N__65784;
    wire N__65781;
    wire N__65778;
    wire N__65775;
    wire N__65772;
    wire N__65765;
    wire N__65762;
    wire N__65759;
    wire N__65756;
    wire N__65751;
    wire N__65744;
    wire N__65735;
    wire N__65728;
    wire N__65725;
    wire N__65722;
    wire N__65719;
    wire N__65716;
    wire N__65713;
    wire N__65710;
    wire N__65707;
    wire N__65706;
    wire N__65705;
    wire N__65704;
    wire N__65701;
    wire N__65700;
    wire N__65699;
    wire N__65696;
    wire N__65693;
    wire N__65690;
    wire N__65681;
    wire N__65678;
    wire N__65675;
    wire N__65670;
    wire N__65667;
    wire N__65664;
    wire N__65661;
    wire N__65658;
    wire N__65655;
    wire N__65652;
    wire N__65649;
    wire N__65646;
    wire N__65645;
    wire N__65642;
    wire N__65639;
    wire N__65638;
    wire N__65635;
    wire N__65632;
    wire N__65629;
    wire N__65628;
    wire N__65623;
    wire N__65618;
    wire N__65615;
    wire N__65612;
    wire N__65605;
    wire N__65602;
    wire N__65597;
    wire N__65592;
    wire N__65589;
    wire N__65582;
    wire N__65579;
    wire N__65576;
    wire N__65571;
    wire N__65568;
    wire N__65563;
    wire N__65560;
    wire N__65555;
    wire N__65550;
    wire N__65543;
    wire N__65540;
    wire N__65535;
    wire N__65532;
    wire N__65515;
    wire N__65512;
    wire N__65509;
    wire N__65506;
    wire N__65503;
    wire N__65500;
    wire N__65499;
    wire N__65496;
    wire N__65493;
    wire N__65490;
    wire N__65485;
    wire N__65484;
    wire N__65483;
    wire N__65482;
    wire N__65477;
    wire N__65472;
    wire N__65469;
    wire N__65468;
    wire N__65465;
    wire N__65462;
    wire N__65459;
    wire N__65456;
    wire N__65453;
    wire N__65446;
    wire N__65443;
    wire N__65442;
    wire N__65439;
    wire N__65436;
    wire N__65431;
    wire N__65428;
    wire N__65425;
    wire N__65422;
    wire N__65419;
    wire N__65416;
    wire N__65413;
    wire N__65410;
    wire N__65407;
    wire N__65404;
    wire N__65403;
    wire N__65402;
    wire N__65399;
    wire N__65394;
    wire N__65389;
    wire N__65386;
    wire N__65383;
    wire N__65380;
    wire N__65377;
    wire N__65374;
    wire N__65371;
    wire N__65368;
    wire N__65365;
    wire N__65362;
    wire N__65359;
    wire N__65356;
    wire N__65353;
    wire N__65350;
    wire N__65347;
    wire N__65344;
    wire N__65343;
    wire N__65340;
    wire N__65337;
    wire N__65334;
    wire N__65331;
    wire N__65326;
    wire N__65323;
    wire N__65320;
    wire N__65317;
    wire N__65314;
    wire N__65311;
    wire N__65308;
    wire N__65305;
    wire N__65304;
    wire N__65303;
    wire N__65300;
    wire N__65295;
    wire N__65290;
    wire N__65287;
    wire N__65286;
    wire N__65281;
    wire N__65278;
    wire N__65277;
    wire N__65274;
    wire N__65273;
    wire N__65270;
    wire N__65267;
    wire N__65264;
    wire N__65261;
    wire N__65254;
    wire N__65251;
    wire N__65248;
    wire N__65245;
    wire N__65242;
    wire N__65239;
    wire N__65236;
    wire N__65235;
    wire N__65232;
    wire N__65229;
    wire N__65228;
    wire N__65225;
    wire N__65222;
    wire N__65219;
    wire N__65212;
    wire N__65209;
    wire N__65206;
    wire N__65203;
    wire N__65200;
    wire N__65197;
    wire N__65194;
    wire N__65191;
    wire N__65188;
    wire N__65185;
    wire N__65182;
    wire N__65179;
    wire N__65176;
    wire N__65173;
    wire N__65170;
    wire N__65167;
    wire N__65164;
    wire N__65161;
    wire N__65158;
    wire N__65155;
    wire N__65152;
    wire N__65149;
    wire N__65146;
    wire N__65143;
    wire N__65140;
    wire N__65137;
    wire N__65134;
    wire N__65131;
    wire N__65130;
    wire N__65129;
    wire N__65128;
    wire N__65127;
    wire N__65126;
    wire N__65121;
    wire N__65118;
    wire N__65115;
    wire N__65112;
    wire N__65109;
    wire N__65108;
    wire N__65099;
    wire N__65096;
    wire N__65093;
    wire N__65090;
    wire N__65085;
    wire N__65080;
    wire N__65079;
    wire N__65078;
    wire N__65077;
    wire N__65076;
    wire N__65075;
    wire N__65074;
    wire N__65073;
    wire N__65072;
    wire N__65071;
    wire N__65070;
    wire N__65047;
    wire N__65044;
    wire N__65041;
    wire N__65038;
    wire N__65035;
    wire N__65032;
    wire N__65029;
    wire N__65026;
    wire N__65023;
    wire N__65020;
    wire N__65017;
    wire N__65014;
    wire N__65011;
    wire N__65008;
    wire N__65005;
    wire N__65002;
    wire N__64999;
    wire N__64996;
    wire N__64993;
    wire N__64990;
    wire N__64987;
    wire N__64984;
    wire N__64981;
    wire N__64978;
    wire N__64975;
    wire N__64972;
    wire N__64969;
    wire N__64966;
    wire N__64963;
    wire N__64960;
    wire N__64957;
    wire N__64954;
    wire N__64951;
    wire N__64948;
    wire N__64945;
    wire N__64942;
    wire N__64939;
    wire N__64936;
    wire N__64933;
    wire N__64930;
    wire N__64927;
    wire N__64924;
    wire N__64921;
    wire N__64918;
    wire N__64915;
    wire N__64912;
    wire N__64909;
    wire N__64906;
    wire N__64903;
    wire N__64900;
    wire N__64897;
    wire N__64894;
    wire N__64891;
    wire N__64888;
    wire N__64885;
    wire N__64882;
    wire N__64879;
    wire N__64878;
    wire N__64877;
    wire N__64874;
    wire N__64871;
    wire N__64868;
    wire N__64865;
    wire N__64862;
    wire N__64859;
    wire N__64856;
    wire N__64851;
    wire N__64846;
    wire N__64843;
    wire N__64840;
    wire N__64839;
    wire N__64836;
    wire N__64835;
    wire N__64834;
    wire N__64831;
    wire N__64828;
    wire N__64823;
    wire N__64820;
    wire N__64817;
    wire N__64814;
    wire N__64807;
    wire N__64804;
    wire N__64803;
    wire N__64802;
    wire N__64801;
    wire N__64798;
    wire N__64797;
    wire N__64792;
    wire N__64789;
    wire N__64784;
    wire N__64781;
    wire N__64776;
    wire N__64771;
    wire N__64768;
    wire N__64765;
    wire N__64762;
    wire N__64759;
    wire N__64756;
    wire N__64755;
    wire N__64752;
    wire N__64747;
    wire N__64744;
    wire N__64743;
    wire N__64740;
    wire N__64737;
    wire N__64734;
    wire N__64729;
    wire N__64726;
    wire N__64723;
    wire N__64720;
    wire N__64717;
    wire N__64714;
    wire N__64711;
    wire N__64708;
    wire N__64705;
    wire N__64702;
    wire N__64699;
    wire N__64696;
    wire N__64693;
    wire N__64690;
    wire N__64687;
    wire N__64684;
    wire N__64681;
    wire N__64678;
    wire N__64675;
    wire N__64672;
    wire N__64669;
    wire N__64666;
    wire N__64663;
    wire N__64660;
    wire N__64659;
    wire N__64658;
    wire N__64653;
    wire N__64650;
    wire N__64647;
    wire N__64644;
    wire N__64639;
    wire N__64636;
    wire N__64635;
    wire N__64634;
    wire N__64629;
    wire N__64628;
    wire N__64625;
    wire N__64622;
    wire N__64619;
    wire N__64616;
    wire N__64611;
    wire N__64608;
    wire N__64603;
    wire N__64600;
    wire N__64599;
    wire N__64598;
    wire N__64593;
    wire N__64592;
    wire N__64589;
    wire N__64586;
    wire N__64583;
    wire N__64580;
    wire N__64575;
    wire N__64572;
    wire N__64567;
    wire N__64564;
    wire N__64563;
    wire N__64560;
    wire N__64559;
    wire N__64556;
    wire N__64553;
    wire N__64550;
    wire N__64547;
    wire N__64544;
    wire N__64541;
    wire N__64538;
    wire N__64533;
    wire N__64528;
    wire N__64525;
    wire N__64524;
    wire N__64523;
    wire N__64520;
    wire N__64517;
    wire N__64514;
    wire N__64511;
    wire N__64508;
    wire N__64505;
    wire N__64502;
    wire N__64499;
    wire N__64494;
    wire N__64489;
    wire N__64486;
    wire N__64483;
    wire N__64480;
    wire N__64479;
    wire N__64478;
    wire N__64475;
    wire N__64470;
    wire N__64467;
    wire N__64464;
    wire N__64459;
    wire N__64456;
    wire N__64453;
    wire N__64452;
    wire N__64451;
    wire N__64448;
    wire N__64443;
    wire N__64438;
    wire N__64435;
    wire N__64432;
    wire N__64429;
    wire N__64426;
    wire N__64425;
    wire N__64424;
    wire N__64421;
    wire N__64416;
    wire N__64411;
    wire N__64408;
    wire N__64405;
    wire N__64404;
    wire N__64401;
    wire N__64398;
    wire N__64397;
    wire N__64396;
    wire N__64393;
    wire N__64390;
    wire N__64385;
    wire N__64382;
    wire N__64377;
    wire N__64374;
    wire N__64371;
    wire N__64366;
    wire N__64363;
    wire N__64362;
    wire N__64357;
    wire N__64354;
    wire N__64353;
    wire N__64352;
    wire N__64349;
    wire N__64348;
    wire N__64347;
    wire N__64346;
    wire N__64343;
    wire N__64340;
    wire N__64337;
    wire N__64330;
    wire N__64321;
    wire N__64318;
    wire N__64315;
    wire N__64312;
    wire N__64309;
    wire N__64306;
    wire N__64303;
    wire N__64300;
    wire N__64297;
    wire N__64296;
    wire N__64293;
    wire N__64290;
    wire N__64289;
    wire N__64284;
    wire N__64281;
    wire N__64276;
    wire N__64273;
    wire N__64272;
    wire N__64267;
    wire N__64266;
    wire N__64263;
    wire N__64260;
    wire N__64255;
    wire N__64252;
    wire N__64251;
    wire N__64246;
    wire N__64245;
    wire N__64242;
    wire N__64239;
    wire N__64234;
    wire N__64231;
    wire N__64230;
    wire N__64225;
    wire N__64222;
    wire N__64219;
    wire N__64216;
    wire N__64213;
    wire N__64210;
    wire N__64207;
    wire N__64204;
    wire N__64201;
    wire N__64198;
    wire N__64195;
    wire N__64192;
    wire N__64189;
    wire N__64188;
    wire N__64183;
    wire N__64180;
    wire N__64177;
    wire N__64174;
    wire N__64173;
    wire N__64170;
    wire N__64167;
    wire N__64164;
    wire N__64161;
    wire N__64158;
    wire N__64155;
    wire N__64150;
    wire N__64147;
    wire N__64144;
    wire N__64141;
    wire N__64138;
    wire N__64135;
    wire N__64132;
    wire N__64129;
    wire N__64126;
    wire N__64123;
    wire N__64120;
    wire N__64117;
    wire N__64114;
    wire N__64111;
    wire N__64108;
    wire N__64105;
    wire N__64104;
    wire N__64099;
    wire N__64096;
    wire N__64095;
    wire N__64090;
    wire N__64087;
    wire N__64086;
    wire N__64085;
    wire N__64082;
    wire N__64079;
    wire N__64076;
    wire N__64069;
    wire N__64066;
    wire N__64063;
    wire N__64062;
    wire N__64057;
    wire N__64054;
    wire N__64053;
    wire N__64052;
    wire N__64049;
    wire N__64046;
    wire N__64043;
    wire N__64036;
    wire N__64033;
    wire N__64030;
    wire N__64029;
    wire N__64026;
    wire N__64023;
    wire N__64018;
    wire N__64015;
    wire N__64014;
    wire N__64011;
    wire N__64008;
    wire N__64005;
    wire N__64002;
    wire N__63999;
    wire N__63994;
    wire N__63993;
    wire N__63990;
    wire N__63987;
    wire N__63984;
    wire N__63981;
    wire N__63976;
    wire N__63975;
    wire N__63972;
    wire N__63969;
    wire N__63964;
    wire N__63961;
    wire N__63960;
    wire N__63959;
    wire N__63956;
    wire N__63951;
    wire N__63946;
    wire N__63943;
    wire N__63942;
    wire N__63941;
    wire N__63934;
    wire N__63931;
    wire N__63928;
    wire N__63925;
    wire N__63922;
    wire N__63919;
    wire N__63916;
    wire N__63913;
    wire N__63910;
    wire N__63907;
    wire N__63904;
    wire N__63901;
    wire N__63898;
    wire N__63895;
    wire N__63892;
    wire N__63889;
    wire N__63886;
    wire N__63883;
    wire N__63882;
    wire N__63879;
    wire N__63876;
    wire N__63871;
    wire N__63870;
    wire N__63867;
    wire N__63864;
    wire N__63859;
    wire N__63858;
    wire N__63853;
    wire N__63850;
    wire N__63849;
    wire N__63846;
    wire N__63843;
    wire N__63838;
    wire N__63837;
    wire N__63836;
    wire N__63833;
    wire N__63830;
    wire N__63827;
    wire N__63820;
    wire N__63817;
    wire N__63814;
    wire N__63811;
    wire N__63808;
    wire N__63807;
    wire N__63802;
    wire N__63799;
    wire N__63796;
    wire N__63793;
    wire N__63790;
    wire N__63789;
    wire N__63784;
    wire N__63781;
    wire N__63778;
    wire N__63777;
    wire N__63772;
    wire N__63769;
    wire N__63766;
    wire N__63763;
    wire N__63762;
    wire N__63761;
    wire N__63758;
    wire N__63753;
    wire N__63748;
    wire N__63745;
    wire N__63742;
    wire N__63739;
    wire N__63736;
    wire N__63735;
    wire N__63734;
    wire N__63727;
    wire N__63724;
    wire N__63721;
    wire N__63718;
    wire N__63715;
    wire N__63712;
    wire N__63709;
    wire N__63708;
    wire N__63707;
    wire N__63706;
    wire N__63705;
    wire N__63704;
    wire N__63703;
    wire N__63702;
    wire N__63699;
    wire N__63698;
    wire N__63695;
    wire N__63694;
    wire N__63691;
    wire N__63690;
    wire N__63687;
    wire N__63686;
    wire N__63683;
    wire N__63682;
    wire N__63679;
    wire N__63678;
    wire N__63677;
    wire N__63674;
    wire N__63673;
    wire N__63662;
    wire N__63645;
    wire N__63638;
    wire N__63635;
    wire N__63632;
    wire N__63629;
    wire N__63622;
    wire N__63619;
    wire N__63616;
    wire N__63615;
    wire N__63612;
    wire N__63609;
    wire N__63606;
    wire N__63603;
    wire N__63600;
    wire N__63595;
    wire N__63594;
    wire N__63589;
    wire N__63586;
    wire N__63583;
    wire N__63582;
    wire N__63577;
    wire N__63574;
    wire N__63573;
    wire N__63568;
    wire N__63565;
    wire N__63564;
    wire N__63559;
    wire N__63556;
    wire N__63553;
    wire N__63550;
    wire N__63547;
    wire N__63544;
    wire N__63543;
    wire N__63538;
    wire N__63535;
    wire N__63532;
    wire N__63529;
    wire N__63526;
    wire N__63523;
    wire N__63520;
    wire N__63517;
    wire N__63514;
    wire N__63511;
    wire N__63508;
    wire N__63505;
    wire N__63502;
    wire N__63499;
    wire N__63496;
    wire N__63493;
    wire N__63490;
    wire N__63487;
    wire N__63484;
    wire N__63481;
    wire N__63478;
    wire N__63475;
    wire N__63472;
    wire N__63469;
    wire N__63466;
    wire N__63463;
    wire N__63460;
    wire N__63457;
    wire N__63454;
    wire N__63451;
    wire N__63448;
    wire N__63445;
    wire N__63442;
    wire N__63439;
    wire N__63436;
    wire N__63433;
    wire N__63430;
    wire N__63427;
    wire N__63424;
    wire N__63421;
    wire N__63418;
    wire N__63415;
    wire N__63412;
    wire N__63409;
    wire N__63406;
    wire N__63403;
    wire N__63400;
    wire N__63397;
    wire N__63394;
    wire N__63391;
    wire N__63388;
    wire N__63385;
    wire N__63382;
    wire N__63379;
    wire N__63376;
    wire N__63373;
    wire N__63370;
    wire N__63367;
    wire N__63364;
    wire N__63361;
    wire N__63358;
    wire N__63355;
    wire N__63352;
    wire N__63349;
    wire N__63346;
    wire N__63343;
    wire N__63340;
    wire N__63339;
    wire N__63336;
    wire N__63333;
    wire N__63330;
    wire N__63325;
    wire N__63322;
    wire N__63319;
    wire N__63316;
    wire N__63313;
    wire N__63310;
    wire N__63307;
    wire N__63306;
    wire N__63303;
    wire N__63300;
    wire N__63297;
    wire N__63292;
    wire N__63289;
    wire N__63286;
    wire N__63283;
    wire N__63280;
    wire N__63277;
    wire N__63274;
    wire N__63271;
    wire N__63268;
    wire N__63267;
    wire N__63264;
    wire N__63261;
    wire N__63256;
    wire N__63253;
    wire N__63250;
    wire N__63247;
    wire N__63244;
    wire N__63241;
    wire N__63238;
    wire N__63237;
    wire N__63234;
    wire N__63231;
    wire N__63226;
    wire N__63223;
    wire N__63220;
    wire N__63217;
    wire N__63214;
    wire N__63213;
    wire N__63210;
    wire N__63207;
    wire N__63204;
    wire N__63201;
    wire N__63196;
    wire N__63193;
    wire N__63190;
    wire N__63187;
    wire N__63184;
    wire N__63181;
    wire N__63178;
    wire N__63177;
    wire N__63174;
    wire N__63171;
    wire N__63166;
    wire N__63163;
    wire N__63160;
    wire N__63157;
    wire N__63156;
    wire N__63155;
    wire N__63154;
    wire N__63151;
    wire N__63146;
    wire N__63143;
    wire N__63138;
    wire N__63133;
    wire N__63130;
    wire N__63127;
    wire N__63126;
    wire N__63121;
    wire N__63118;
    wire N__63115;
    wire N__63112;
    wire N__63109;
    wire N__63106;
    wire N__63103;
    wire N__63100;
    wire N__63097;
    wire N__63094;
    wire N__63091;
    wire N__63088;
    wire N__63085;
    wire N__63082;
    wire N__63079;
    wire N__63076;
    wire N__63073;
    wire N__63070;
    wire N__63067;
    wire N__63064;
    wire N__63061;
    wire N__63058;
    wire N__63055;
    wire N__63052;
    wire N__63049;
    wire N__63046;
    wire N__63043;
    wire N__63040;
    wire N__63037;
    wire N__63034;
    wire N__63031;
    wire N__63028;
    wire N__63025;
    wire N__63022;
    wire N__63019;
    wire N__63016;
    wire N__63015;
    wire N__63012;
    wire N__63009;
    wire N__63006;
    wire N__63005;
    wire N__63002;
    wire N__62999;
    wire N__62996;
    wire N__62993;
    wire N__62986;
    wire N__62983;
    wire N__62980;
    wire N__62977;
    wire N__62974;
    wire N__62971;
    wire N__62968;
    wire N__62965;
    wire N__62964;
    wire N__62959;
    wire N__62956;
    wire N__62953;
    wire N__62950;
    wire N__62947;
    wire N__62944;
    wire N__62941;
    wire N__62938;
    wire N__62935;
    wire N__62932;
    wire N__62929;
    wire N__62926;
    wire N__62923;
    wire N__62920;
    wire N__62917;
    wire N__62916;
    wire N__62915;
    wire N__62912;
    wire N__62907;
    wire N__62902;
    wire N__62899;
    wire N__62896;
    wire N__62895;
    wire N__62894;
    wire N__62893;
    wire N__62890;
    wire N__62889;
    wire N__62886;
    wire N__62885;
    wire N__62884;
    wire N__62883;
    wire N__62882;
    wire N__62881;
    wire N__62880;
    wire N__62877;
    wire N__62876;
    wire N__62865;
    wire N__62862;
    wire N__62861;
    wire N__62858;
    wire N__62857;
    wire N__62854;
    wire N__62853;
    wire N__62850;
    wire N__62849;
    wire N__62842;
    wire N__62839;
    wire N__62822;
    wire N__62819;
    wire N__62812;
    wire N__62809;
    wire N__62806;
    wire N__62803;
    wire N__62800;
    wire N__62797;
    wire N__62794;
    wire N__62793;
    wire N__62792;
    wire N__62791;
    wire N__62790;
    wire N__62789;
    wire N__62788;
    wire N__62787;
    wire N__62784;
    wire N__62783;
    wire N__62780;
    wire N__62777;
    wire N__62776;
    wire N__62773;
    wire N__62772;
    wire N__62771;
    wire N__62770;
    wire N__62769;
    wire N__62768;
    wire N__62759;
    wire N__62756;
    wire N__62751;
    wire N__62748;
    wire N__62743;
    wire N__62742;
    wire N__62739;
    wire N__62736;
    wire N__62733;
    wire N__62730;
    wire N__62727;
    wire N__62724;
    wire N__62721;
    wire N__62714;
    wire N__62707;
    wire N__62704;
    wire N__62699;
    wire N__62696;
    wire N__62691;
    wire N__62684;
    wire N__62677;
    wire N__62676;
    wire N__62673;
    wire N__62670;
    wire N__62667;
    wire N__62664;
    wire N__62659;
    wire N__62656;
    wire N__62653;
    wire N__62650;
    wire N__62647;
    wire N__62644;
    wire N__62641;
    wire N__62638;
    wire N__62635;
    wire N__62632;
    wire N__62631;
    wire N__62630;
    wire N__62627;
    wire N__62622;
    wire N__62617;
    wire N__62614;
    wire N__62611;
    wire N__62608;
    wire N__62607;
    wire N__62606;
    wire N__62603;
    wire N__62600;
    wire N__62597;
    wire N__62592;
    wire N__62589;
    wire N__62584;
    wire N__62581;
    wire N__62578;
    wire N__62575;
    wire N__62572;
    wire N__62569;
    wire N__62566;
    wire N__62563;
    wire N__62560;
    wire N__62557;
    wire N__62554;
    wire N__62551;
    wire N__62548;
    wire N__62545;
    wire N__62542;
    wire N__62539;
    wire N__62536;
    wire N__62533;
    wire N__62530;
    wire N__62527;
    wire N__62524;
    wire N__62521;
    wire N__62518;
    wire N__62515;
    wire N__62512;
    wire N__62509;
    wire N__62506;
    wire N__62503;
    wire N__62500;
    wire N__62497;
    wire N__62494;
    wire N__62491;
    wire N__62488;
    wire N__62487;
    wire N__62484;
    wire N__62481;
    wire N__62480;
    wire N__62475;
    wire N__62472;
    wire N__62467;
    wire N__62464;
    wire N__62461;
    wire N__62458;
    wire N__62455;
    wire N__62452;
    wire N__62451;
    wire N__62448;
    wire N__62445;
    wire N__62440;
    wire N__62437;
    wire N__62434;
    wire N__62431;
    wire N__62428;
    wire N__62425;
    wire N__62422;
    wire N__62421;
    wire N__62418;
    wire N__62415;
    wire N__62412;
    wire N__62409;
    wire N__62404;
    wire N__62401;
    wire N__62398;
    wire N__62395;
    wire N__62392;
    wire N__62389;
    wire N__62386;
    wire N__62383;
    wire N__62380;
    wire N__62377;
    wire N__62374;
    wire N__62371;
    wire N__62368;
    wire N__62365;
    wire N__62362;
    wire N__62359;
    wire N__62356;
    wire N__62353;
    wire N__62350;
    wire N__62347;
    wire N__62344;
    wire N__62343;
    wire N__62340;
    wire N__62337;
    wire N__62332;
    wire N__62329;
    wire N__62328;
    wire N__62323;
    wire N__62320;
    wire N__62317;
    wire N__62314;
    wire N__62311;
    wire N__62308;
    wire N__62307;
    wire N__62304;
    wire N__62301;
    wire N__62296;
    wire N__62295;
    wire N__62292;
    wire N__62289;
    wire N__62284;
    wire N__62281;
    wire N__62280;
    wire N__62275;
    wire N__62272;
    wire N__62271;
    wire N__62266;
    wire N__62263;
    wire N__62260;
    wire N__62259;
    wire N__62256;
    wire N__62253;
    wire N__62248;
    wire N__62245;
    wire N__62244;
    wire N__62241;
    wire N__62238;
    wire N__62233;
    wire N__62232;
    wire N__62229;
    wire N__62226;
    wire N__62223;
    wire N__62218;
    wire N__62217;
    wire N__62214;
    wire N__62211;
    wire N__62208;
    wire N__62203;
    wire N__62200;
    wire N__62197;
    wire N__62194;
    wire N__62193;
    wire N__62190;
    wire N__62187;
    wire N__62182;
    wire N__62181;
    wire N__62178;
    wire N__62175;
    wire N__62170;
    wire N__62169;
    wire N__62166;
    wire N__62163;
    wire N__62160;
    wire N__62157;
    wire N__62152;
    wire N__62151;
    wire N__62148;
    wire N__62145;
    wire N__62142;
    wire N__62139;
    wire N__62136;
    wire N__62131;
    wire N__62128;
    wire N__62125;
    wire N__62122;
    wire N__62119;
    wire N__62118;
    wire N__62115;
    wire N__62112;
    wire N__62107;
    wire N__62106;
    wire N__62103;
    wire N__62100;
    wire N__62095;
    wire N__62092;
    wire N__62089;
    wire N__62086;
    wire N__62083;
    wire N__62080;
    wire N__62079;
    wire N__62076;
    wire N__62073;
    wire N__62068;
    wire N__62065;
    wire N__62064;
    wire N__62061;
    wire N__62058;
    wire N__62057;
    wire N__62056;
    wire N__62051;
    wire N__62046;
    wire N__62041;
    wire N__62040;
    wire N__62039;
    wire N__62036;
    wire N__62031;
    wire N__62028;
    wire N__62025;
    wire N__62022;
    wire N__62017;
    wire N__62014;
    wire N__62013;
    wire N__62010;
    wire N__62007;
    wire N__62002;
    wire N__61999;
    wire N__61996;
    wire N__61993;
    wire N__61990;
    wire N__61987;
    wire N__61984;
    wire N__61981;
    wire N__61978;
    wire N__61975;
    wire N__61972;
    wire N__61969;
    wire N__61968;
    wire N__61967;
    wire N__61966;
    wire N__61963;
    wire N__61958;
    wire N__61955;
    wire N__61952;
    wire N__61949;
    wire N__61944;
    wire N__61941;
    wire N__61936;
    wire N__61933;
    wire N__61932;
    wire N__61929;
    wire N__61926;
    wire N__61921;
    wire N__61918;
    wire N__61917;
    wire N__61914;
    wire N__61911;
    wire N__61906;
    wire N__61903;
    wire N__61900;
    wire N__61897;
    wire N__61894;
    wire N__61893;
    wire N__61890;
    wire N__61887;
    wire N__61882;
    wire N__61879;
    wire N__61876;
    wire N__61873;
    wire N__61870;
    wire N__61867;
    wire N__61864;
    wire N__61861;
    wire N__61858;
    wire N__61855;
    wire N__61854;
    wire N__61851;
    wire N__61848;
    wire N__61843;
    wire N__61840;
    wire N__61837;
    wire N__61836;
    wire N__61833;
    wire N__61830;
    wire N__61825;
    wire N__61824;
    wire N__61821;
    wire N__61818;
    wire N__61813;
    wire N__61810;
    wire N__61807;
    wire N__61804;
    wire N__61801;
    wire N__61798;
    wire N__61795;
    wire N__61794;
    wire N__61793;
    wire N__61786;
    wire N__61783;
    wire N__61782;
    wire N__61779;
    wire N__61778;
    wire N__61775;
    wire N__61772;
    wire N__61767;
    wire N__61764;
    wire N__61759;
    wire N__61756;
    wire N__61753;
    wire N__61750;
    wire N__61747;
    wire N__61744;
    wire N__61741;
    wire N__61738;
    wire N__61737;
    wire N__61732;
    wire N__61729;
    wire N__61726;
    wire N__61723;
    wire N__61720;
    wire N__61717;
    wire N__61716;
    wire N__61711;
    wire N__61708;
    wire N__61707;
    wire N__61706;
    wire N__61705;
    wire N__61704;
    wire N__61701;
    wire N__61698;
    wire N__61691;
    wire N__61684;
    wire N__61681;
    wire N__61680;
    wire N__61675;
    wire N__61672;
    wire N__61669;
    wire N__61668;
    wire N__61665;
    wire N__61660;
    wire N__61657;
    wire N__61654;
    wire N__61651;
    wire N__61650;
    wire N__61647;
    wire N__61644;
    wire N__61641;
    wire N__61636;
    wire N__61633;
    wire N__61632;
    wire N__61629;
    wire N__61626;
    wire N__61623;
    wire N__61620;
    wire N__61617;
    wire N__61612;
    wire N__61609;
    wire N__61606;
    wire N__61603;
    wire N__61600;
    wire N__61597;
    wire N__61594;
    wire N__61591;
    wire N__61588;
    wire N__61585;
    wire N__61582;
    wire N__61579;
    wire N__61578;
    wire N__61575;
    wire N__61572;
    wire N__61567;
    wire N__61564;
    wire N__61561;
    wire N__61558;
    wire N__61557;
    wire N__61554;
    wire N__61551;
    wire N__61546;
    wire N__61545;
    wire N__61542;
    wire N__61539;
    wire N__61534;
    wire N__61531;
    wire N__61528;
    wire N__61525;
    wire N__61522;
    wire N__61519;
    wire N__61516;
    wire N__61513;
    wire N__61510;
    wire N__61507;
    wire N__61504;
    wire N__61501;
    wire N__61498;
    wire N__61495;
    wire N__61492;
    wire N__61489;
    wire N__61486;
    wire N__61483;
    wire N__61480;
    wire N__61477;
    wire N__61476;
    wire N__61471;
    wire N__61468;
    wire N__61467;
    wire N__61462;
    wire N__61459;
    wire N__61456;
    wire N__61453;
    wire N__61450;
    wire N__61447;
    wire N__61444;
    wire N__61443;
    wire N__61440;
    wire N__61437;
    wire N__61434;
    wire N__61429;
    wire N__61428;
    wire N__61423;
    wire N__61420;
    wire N__61417;
    wire N__61414;
    wire N__61411;
    wire N__61408;
    wire N__61405;
    wire N__61404;
    wire N__61399;
    wire N__61396;
    wire N__61393;
    wire N__61390;
    wire N__61387;
    wire N__61384;
    wire N__61381;
    wire N__61378;
    wire N__61375;
    wire N__61372;
    wire N__61371;
    wire N__61368;
    wire N__61365;
    wire N__61364;
    wire N__61363;
    wire N__61360;
    wire N__61357;
    wire N__61352;
    wire N__61345;
    wire N__61342;
    wire N__61339;
    wire N__61338;
    wire N__61337;
    wire N__61336;
    wire N__61335;
    wire N__61334;
    wire N__61331;
    wire N__61328;
    wire N__61319;
    wire N__61312;
    wire N__61309;
    wire N__61306;
    wire N__61303;
    wire N__61302;
    wire N__61299;
    wire N__61296;
    wire N__61291;
    wire N__61290;
    wire N__61287;
    wire N__61284;
    wire N__61279;
    wire N__61276;
    wire N__61273;
    wire N__61270;
    wire N__61267;
    wire N__61264;
    wire N__61261;
    wire N__61258;
    wire N__61255;
    wire N__61254;
    wire N__61249;
    wire N__61246;
    wire N__61243;
    wire N__61242;
    wire N__61237;
    wire N__61234;
    wire N__61231;
    wire N__61228;
    wire N__61225;
    wire N__61222;
    wire N__61219;
    wire N__61216;
    wire N__61215;
    wire N__61214;
    wire N__61207;
    wire N__61204;
    wire N__61201;
    wire N__61198;
    wire N__61195;
    wire N__61192;
    wire N__61189;
    wire N__61186;
    wire N__61183;
    wire N__61180;
    wire N__61177;
    wire N__61174;
    wire N__61171;
    wire N__61168;
    wire N__61165;
    wire N__61162;
    wire N__61159;
    wire N__61156;
    wire N__61153;
    wire N__61152;
    wire N__61149;
    wire N__61146;
    wire N__61141;
    wire N__61140;
    wire N__61135;
    wire N__61132;
    wire N__61129;
    wire N__61126;
    wire N__61123;
    wire N__61120;
    wire N__61117;
    wire N__61114;
    wire N__61111;
    wire N__61108;
    wire N__61105;
    wire N__61102;
    wire N__61099;
    wire N__61096;
    wire N__61093;
    wire N__61092;
    wire N__61091;
    wire N__61088;
    wire N__61083;
    wire N__61078;
    wire N__61075;
    wire N__61072;
    wire N__61069;
    wire N__61066;
    wire N__61065;
    wire N__61062;
    wire N__61059;
    wire N__61054;
    wire N__61051;
    wire N__61048;
    wire N__61045;
    wire N__61042;
    wire N__61039;
    wire N__61036;
    wire N__61033;
    wire N__61030;
    wire N__61027;
    wire N__61024;
    wire N__61021;
    wire N__61018;
    wire N__61015;
    wire N__61014;
    wire N__61011;
    wire N__61008;
    wire N__61003;
    wire N__61000;
    wire N__60997;
    wire N__60994;
    wire N__60991;
    wire N__60988;
    wire N__60985;
    wire N__60982;
    wire N__60979;
    wire N__60976;
    wire N__60975;
    wire N__60970;
    wire N__60967;
    wire N__60964;
    wire N__60961;
    wire N__60958;
    wire N__60955;
    wire N__60952;
    wire N__60949;
    wire N__60946;
    wire N__60943;
    wire N__60940;
    wire N__60937;
    wire N__60934;
    wire N__60931;
    wire N__60928;
    wire N__60925;
    wire N__60922;
    wire N__60919;
    wire N__60916;
    wire N__60913;
    wire N__60910;
    wire N__60907;
    wire N__60904;
    wire N__60901;
    wire N__60898;
    wire N__60895;
    wire N__60892;
    wire N__60889;
    wire N__60886;
    wire N__60883;
    wire N__60880;
    wire N__60877;
    wire N__60874;
    wire N__60871;
    wire N__60868;
    wire N__60865;
    wire N__60862;
    wire N__60861;
    wire N__60856;
    wire N__60853;
    wire N__60850;
    wire N__60847;
    wire N__60844;
    wire N__60841;
    wire N__60838;
    wire N__60835;
    wire N__60832;
    wire N__60829;
    wire N__60826;
    wire N__60823;
    wire N__60820;
    wire N__60817;
    wire N__60814;
    wire N__60811;
    wire N__60808;
    wire N__60805;
    wire N__60804;
    wire N__60799;
    wire N__60798;
    wire N__60795;
    wire N__60792;
    wire N__60791;
    wire N__60790;
    wire N__60789;
    wire N__60786;
    wire N__60785;
    wire N__60784;
    wire N__60783;
    wire N__60780;
    wire N__60773;
    wire N__60770;
    wire N__60763;
    wire N__60754;
    wire N__60753;
    wire N__60752;
    wire N__60749;
    wire N__60748;
    wire N__60747;
    wire N__60746;
    wire N__60745;
    wire N__60744;
    wire N__60743;
    wire N__60740;
    wire N__60737;
    wire N__60724;
    wire N__60719;
    wire N__60716;
    wire N__60715;
    wire N__60712;
    wire N__60711;
    wire N__60706;
    wire N__60703;
    wire N__60700;
    wire N__60699;
    wire N__60698;
    wire N__60695;
    wire N__60692;
    wire N__60691;
    wire N__60688;
    wire N__60685;
    wire N__60680;
    wire N__60677;
    wire N__60674;
    wire N__60671;
    wire N__60668;
    wire N__60655;
    wire N__60652;
    wire N__60649;
    wire N__60646;
    wire N__60643;
    wire N__60640;
    wire N__60637;
    wire N__60634;
    wire N__60631;
    wire N__60628;
    wire N__60625;
    wire N__60622;
    wire N__60619;
    wire N__60618;
    wire N__60613;
    wire N__60610;
    wire N__60607;
    wire N__60604;
    wire N__60601;
    wire N__60598;
    wire N__60595;
    wire N__60594;
    wire N__60589;
    wire N__60586;
    wire N__60585;
    wire N__60580;
    wire N__60577;
    wire N__60576;
    wire N__60573;
    wire N__60570;
    wire N__60565;
    wire N__60562;
    wire N__60559;
    wire N__60556;
    wire N__60553;
    wire N__60550;
    wire N__60549;
    wire N__60548;
    wire N__60545;
    wire N__60542;
    wire N__60541;
    wire N__60538;
    wire N__60537;
    wire N__60536;
    wire N__60533;
    wire N__60530;
    wire N__60527;
    wire N__60524;
    wire N__60521;
    wire N__60518;
    wire N__60511;
    wire N__60508;
    wire N__60503;
    wire N__60500;
    wire N__60497;
    wire N__60494;
    wire N__60491;
    wire N__60484;
    wire N__60481;
    wire N__60478;
    wire N__60477;
    wire N__60472;
    wire N__60469;
    wire N__60468;
    wire N__60467;
    wire N__60464;
    wire N__60459;
    wire N__60454;
    wire N__60453;
    wire N__60452;
    wire N__60451;
    wire N__60450;
    wire N__60449;
    wire N__60446;
    wire N__60445;
    wire N__60444;
    wire N__60443;
    wire N__60442;
    wire N__60439;
    wire N__60434;
    wire N__60431;
    wire N__60430;
    wire N__60427;
    wire N__60424;
    wire N__60421;
    wire N__60416;
    wire N__60413;
    wire N__60406;
    wire N__60403;
    wire N__60400;
    wire N__60397;
    wire N__60394;
    wire N__60391;
    wire N__60388;
    wire N__60385;
    wire N__60380;
    wire N__60377;
    wire N__60374;
    wire N__60367;
    wire N__60364;
    wire N__60355;
    wire N__60354;
    wire N__60353;
    wire N__60346;
    wire N__60343;
    wire N__60340;
    wire N__60337;
    wire N__60334;
    wire N__60333;
    wire N__60332;
    wire N__60327;
    wire N__60326;
    wire N__60323;
    wire N__60322;
    wire N__60321;
    wire N__60318;
    wire N__60315;
    wire N__60310;
    wire N__60307;
    wire N__60298;
    wire N__60295;
    wire N__60292;
    wire N__60289;
    wire N__60286;
    wire N__60285;
    wire N__60284;
    wire N__60281;
    wire N__60276;
    wire N__60271;
    wire N__60268;
    wire N__60267;
    wire N__60264;
    wire N__60261;
    wire N__60256;
    wire N__60253;
    wire N__60250;
    wire N__60247;
    wire N__60244;
    wire N__60241;
    wire N__60240;
    wire N__60239;
    wire N__60236;
    wire N__60231;
    wire N__60226;
    wire N__60223;
    wire N__60220;
    wire N__60219;
    wire N__60216;
    wire N__60213;
    wire N__60210;
    wire N__60207;
    wire N__60204;
    wire N__60201;
    wire N__60196;
    wire N__60195;
    wire N__60194;
    wire N__60187;
    wire N__60186;
    wire N__60185;
    wire N__60184;
    wire N__60183;
    wire N__60182;
    wire N__60181;
    wire N__60180;
    wire N__60179;
    wire N__60176;
    wire N__60163;
    wire N__60158;
    wire N__60155;
    wire N__60150;
    wire N__60149;
    wire N__60146;
    wire N__60143;
    wire N__60140;
    wire N__60133;
    wire N__60132;
    wire N__60131;
    wire N__60124;
    wire N__60123;
    wire N__60122;
    wire N__60119;
    wire N__60114;
    wire N__60109;
    wire N__60108;
    wire N__60105;
    wire N__60102;
    wire N__60099;
    wire N__60096;
    wire N__60091;
    wire N__60088;
    wire N__60085;
    wire N__60082;
    wire N__60081;
    wire N__60078;
    wire N__60077;
    wire N__60074;
    wire N__60071;
    wire N__60066;
    wire N__60061;
    wire N__60058;
    wire N__60057;
    wire N__60054;
    wire N__60051;
    wire N__60046;
    wire N__60043;
    wire N__60040;
    wire N__60037;
    wire N__60036;
    wire N__60033;
    wire N__60030;
    wire N__60029;
    wire N__60024;
    wire N__60021;
    wire N__60020;
    wire N__60017;
    wire N__60014;
    wire N__60011;
    wire N__60008;
    wire N__60005;
    wire N__60002;
    wire N__59995;
    wire N__59992;
    wire N__59991;
    wire N__59990;
    wire N__59987;
    wire N__59984;
    wire N__59981;
    wire N__59978;
    wire N__59975;
    wire N__59972;
    wire N__59971;
    wire N__59968;
    wire N__59963;
    wire N__59960;
    wire N__59957;
    wire N__59954;
    wire N__59951;
    wire N__59950;
    wire N__59947;
    wire N__59942;
    wire N__59939;
    wire N__59932;
    wire N__59929;
    wire N__59926;
    wire N__59923;
    wire N__59922;
    wire N__59917;
    wire N__59916;
    wire N__59915;
    wire N__59912;
    wire N__59907;
    wire N__59902;
    wire N__59899;
    wire N__59896;
    wire N__59893;
    wire N__59890;
    wire N__59887;
    wire N__59884;
    wire N__59881;
    wire N__59878;
    wire N__59877;
    wire N__59872;
    wire N__59869;
    wire N__59866;
    wire N__59863;
    wire N__59860;
    wire N__59857;
    wire N__59856;
    wire N__59855;
    wire N__59848;
    wire N__59845;
    wire N__59844;
    wire N__59843;
    wire N__59838;
    wire N__59835;
    wire N__59830;
    wire N__59827;
    wire N__59824;
    wire N__59823;
    wire N__59818;
    wire N__59817;
    wire N__59816;
    wire N__59815;
    wire N__59814;
    wire N__59811;
    wire N__59808;
    wire N__59803;
    wire N__59800;
    wire N__59791;
    wire N__59788;
    wire N__59785;
    wire N__59784;
    wire N__59783;
    wire N__59782;
    wire N__59781;
    wire N__59778;
    wire N__59773;
    wire N__59770;
    wire N__59769;
    wire N__59768;
    wire N__59767;
    wire N__59764;
    wire N__59759;
    wire N__59756;
    wire N__59753;
    wire N__59752;
    wire N__59749;
    wire N__59746;
    wire N__59743;
    wire N__59736;
    wire N__59733;
    wire N__59730;
    wire N__59719;
    wire N__59718;
    wire N__59717;
    wire N__59716;
    wire N__59715;
    wire N__59708;
    wire N__59705;
    wire N__59702;
    wire N__59701;
    wire N__59700;
    wire N__59699;
    wire N__59694;
    wire N__59691;
    wire N__59688;
    wire N__59683;
    wire N__59680;
    wire N__59673;
    wire N__59668;
    wire N__59667;
    wire N__59666;
    wire N__59661;
    wire N__59658;
    wire N__59655;
    wire N__59652;
    wire N__59651;
    wire N__59646;
    wire N__59643;
    wire N__59638;
    wire N__59637;
    wire N__59636;
    wire N__59633;
    wire N__59630;
    wire N__59627;
    wire N__59620;
    wire N__59619;
    wire N__59618;
    wire N__59615;
    wire N__59612;
    wire N__59607;
    wire N__59602;
    wire N__59601;
    wire N__59600;
    wire N__59597;
    wire N__59596;
    wire N__59591;
    wire N__59588;
    wire N__59585;
    wire N__59582;
    wire N__59579;
    wire N__59576;
    wire N__59569;
    wire N__59566;
    wire N__59563;
    wire N__59562;
    wire N__59561;
    wire N__59556;
    wire N__59553;
    wire N__59550;
    wire N__59545;
    wire N__59544;
    wire N__59539;
    wire N__59538;
    wire N__59535;
    wire N__59532;
    wire N__59527;
    wire N__59524;
    wire N__59521;
    wire N__59518;
    wire N__59515;
    wire N__59512;
    wire N__59509;
    wire N__59506;
    wire N__59503;
    wire N__59500;
    wire N__59499;
    wire N__59496;
    wire N__59493;
    wire N__59492;
    wire N__59487;
    wire N__59484;
    wire N__59479;
    wire N__59476;
    wire N__59475;
    wire N__59472;
    wire N__59469;
    wire N__59468;
    wire N__59465;
    wire N__59462;
    wire N__59459;
    wire N__59452;
    wire N__59451;
    wire N__59450;
    wire N__59447;
    wire N__59444;
    wire N__59441;
    wire N__59438;
    wire N__59431;
    wire N__59430;
    wire N__59427;
    wire N__59426;
    wire N__59423;
    wire N__59420;
    wire N__59417;
    wire N__59410;
    wire N__59409;
    wire N__59406;
    wire N__59403;
    wire N__59400;
    wire N__59399;
    wire N__59396;
    wire N__59395;
    wire N__59392;
    wire N__59389;
    wire N__59386;
    wire N__59383;
    wire N__59378;
    wire N__59373;
    wire N__59370;
    wire N__59367;
    wire N__59362;
    wire N__59361;
    wire N__59356;
    wire N__59353;
    wire N__59350;
    wire N__59347;
    wire N__59344;
    wire N__59341;
    wire N__59338;
    wire N__59335;
    wire N__59332;
    wire N__59331;
    wire N__59328;
    wire N__59325;
    wire N__59320;
    wire N__59317;
    wire N__59314;
    wire N__59311;
    wire N__59308;
    wire N__59307;
    wire N__59304;
    wire N__59301;
    wire N__59298;
    wire N__59293;
    wire N__59290;
    wire N__59287;
    wire N__59284;
    wire N__59283;
    wire N__59280;
    wire N__59277;
    wire N__59272;
    wire N__59269;
    wire N__59266;
    wire N__59263;
    wire N__59260;
    wire N__59257;
    wire N__59256;
    wire N__59255;
    wire N__59254;
    wire N__59253;
    wire N__59252;
    wire N__59251;
    wire N__59250;
    wire N__59249;
    wire N__59246;
    wire N__59243;
    wire N__59242;
    wire N__59241;
    wire N__59238;
    wire N__59237;
    wire N__59230;
    wire N__59217;
    wire N__59210;
    wire N__59207;
    wire N__59200;
    wire N__59199;
    wire N__59198;
    wire N__59195;
    wire N__59194;
    wire N__59193;
    wire N__59190;
    wire N__59181;
    wire N__59176;
    wire N__59175;
    wire N__59172;
    wire N__59169;
    wire N__59166;
    wire N__59163;
    wire N__59160;
    wire N__59157;
    wire N__59154;
    wire N__59149;
    wire N__59148;
    wire N__59145;
    wire N__59142;
    wire N__59141;
    wire N__59138;
    wire N__59135;
    wire N__59132;
    wire N__59129;
    wire N__59126;
    wire N__59123;
    wire N__59120;
    wire N__59115;
    wire N__59110;
    wire N__59107;
    wire N__59104;
    wire N__59101;
    wire N__59098;
    wire N__59095;
    wire N__59092;
    wire N__59089;
    wire N__59086;
    wire N__59083;
    wire N__59080;
    wire N__59079;
    wire N__59078;
    wire N__59077;
    wire N__59074;
    wire N__59071;
    wire N__59066;
    wire N__59059;
    wire N__59056;
    wire N__59053;
    wire N__59050;
    wire N__59047;
    wire N__59044;
    wire N__59041;
    wire N__59040;
    wire N__59039;
    wire N__59036;
    wire N__59033;
    wire N__59030;
    wire N__59025;
    wire N__59020;
    wire N__59017;
    wire N__59014;
    wire N__59011;
    wire N__59008;
    wire N__59005;
    wire N__59002;
    wire N__58999;
    wire N__58996;
    wire N__58993;
    wire N__58990;
    wire N__58989;
    wire N__58988;
    wire N__58987;
    wire N__58982;
    wire N__58977;
    wire N__58972;
    wire N__58969;
    wire N__58966;
    wire N__58963;
    wire N__58960;
    wire N__58957;
    wire N__58954;
    wire N__58951;
    wire N__58948;
    wire N__58945;
    wire N__58944;
    wire N__58941;
    wire N__58938;
    wire N__58933;
    wire N__58930;
    wire N__58927;
    wire N__58924;
    wire N__58921;
    wire N__58918;
    wire N__58915;
    wire N__58914;
    wire N__58913;
    wire N__58912;
    wire N__58911;
    wire N__58906;
    wire N__58899;
    wire N__58894;
    wire N__58891;
    wire N__58888;
    wire N__58885;
    wire N__58882;
    wire N__58879;
    wire N__58876;
    wire N__58873;
    wire N__58872;
    wire N__58871;
    wire N__58868;
    wire N__58867;
    wire N__58866;
    wire N__58863;
    wire N__58862;
    wire N__58855;
    wire N__58852;
    wire N__58849;
    wire N__58846;
    wire N__58843;
    wire N__58840;
    wire N__58839;
    wire N__58836;
    wire N__58829;
    wire N__58826;
    wire N__58819;
    wire N__58816;
    wire N__58813;
    wire N__58810;
    wire N__58807;
    wire N__58804;
    wire N__58801;
    wire N__58798;
    wire N__58795;
    wire N__58792;
    wire N__58789;
    wire N__58786;
    wire N__58783;
    wire N__58780;
    wire N__58777;
    wire N__58774;
    wire N__58771;
    wire N__58768;
    wire N__58765;
    wire N__58762;
    wire N__58759;
    wire N__58756;
    wire N__58753;
    wire N__58750;
    wire N__58747;
    wire N__58744;
    wire N__58741;
    wire N__58738;
    wire N__58735;
    wire N__58732;
    wire N__58729;
    wire N__58726;
    wire N__58723;
    wire N__58720;
    wire N__58717;
    wire N__58714;
    wire N__58711;
    wire N__58708;
    wire N__58705;
    wire N__58702;
    wire N__58699;
    wire N__58696;
    wire N__58693;
    wire N__58690;
    wire N__58687;
    wire N__58684;
    wire N__58681;
    wire N__58678;
    wire N__58675;
    wire N__58672;
    wire N__58669;
    wire N__58666;
    wire N__58663;
    wire N__58660;
    wire N__58657;
    wire N__58654;
    wire N__58653;
    wire N__58650;
    wire N__58649;
    wire N__58646;
    wire N__58643;
    wire N__58638;
    wire N__58635;
    wire N__58632;
    wire N__58629;
    wire N__58626;
    wire N__58621;
    wire N__58618;
    wire N__58617;
    wire N__58614;
    wire N__58611;
    wire N__58608;
    wire N__58607;
    wire N__58606;
    wire N__58601;
    wire N__58596;
    wire N__58591;
    wire N__58588;
    wire N__58585;
    wire N__58584;
    wire N__58579;
    wire N__58578;
    wire N__58575;
    wire N__58572;
    wire N__58571;
    wire N__58570;
    wire N__58567;
    wire N__58564;
    wire N__58559;
    wire N__58552;
    wire N__58549;
    wire N__58546;
    wire N__58543;
    wire N__58540;
    wire N__58539;
    wire N__58538;
    wire N__58535;
    wire N__58532;
    wire N__58529;
    wire N__58526;
    wire N__58521;
    wire N__58516;
    wire N__58513;
    wire N__58510;
    wire N__58507;
    wire N__58504;
    wire N__58501;
    wire N__58498;
    wire N__58495;
    wire N__58492;
    wire N__58489;
    wire N__58486;
    wire N__58483;
    wire N__58480;
    wire N__58477;
    wire N__58474;
    wire N__58471;
    wire N__58468;
    wire N__58465;
    wire N__58464;
    wire N__58463;
    wire N__58460;
    wire N__58459;
    wire N__58454;
    wire N__58451;
    wire N__58448;
    wire N__58445;
    wire N__58438;
    wire N__58435;
    wire N__58432;
    wire N__58431;
    wire N__58430;
    wire N__58429;
    wire N__58426;
    wire N__58421;
    wire N__58418;
    wire N__58413;
    wire N__58408;
    wire N__58405;
    wire N__58402;
    wire N__58401;
    wire N__58398;
    wire N__58395;
    wire N__58394;
    wire N__58391;
    wire N__58388;
    wire N__58385;
    wire N__58382;
    wire N__58377;
    wire N__58372;
    wire N__58369;
    wire N__58368;
    wire N__58365;
    wire N__58364;
    wire N__58361;
    wire N__58358;
    wire N__58355;
    wire N__58352;
    wire N__58349;
    wire N__58346;
    wire N__58343;
    wire N__58340;
    wire N__58335;
    wire N__58330;
    wire N__58327;
    wire N__58326;
    wire N__58323;
    wire N__58320;
    wire N__58317;
    wire N__58314;
    wire N__58311;
    wire N__58306;
    wire N__58303;
    wire N__58300;
    wire N__58297;
    wire N__58294;
    wire N__58291;
    wire N__58288;
    wire N__58285;
    wire N__58284;
    wire N__58283;
    wire N__58280;
    wire N__58275;
    wire N__58272;
    wire N__58269;
    wire N__58264;
    wire N__58261;
    wire N__58258;
    wire N__58255;
    wire N__58254;
    wire N__58251;
    wire N__58248;
    wire N__58245;
    wire N__58240;
    wire N__58237;
    wire N__58234;
    wire N__58231;
    wire N__58230;
    wire N__58229;
    wire N__58226;
    wire N__58221;
    wire N__58218;
    wire N__58215;
    wire N__58210;
    wire N__58207;
    wire N__58204;
    wire N__58201;
    wire N__58200;
    wire N__58199;
    wire N__58196;
    wire N__58191;
    wire N__58188;
    wire N__58185;
    wire N__58180;
    wire N__58177;
    wire N__58174;
    wire N__58171;
    wire N__58168;
    wire N__58165;
    wire N__58162;
    wire N__58159;
    wire N__58156;
    wire N__58155;
    wire N__58154;
    wire N__58151;
    wire N__58146;
    wire N__58141;
    wire N__58138;
    wire N__58135;
    wire N__58132;
    wire N__58129;
    wire N__58126;
    wire N__58123;
    wire N__58122;
    wire N__58117;
    wire N__58114;
    wire N__58111;
    wire N__58110;
    wire N__58105;
    wire N__58102;
    wire N__58099;
    wire N__58096;
    wire N__58093;
    wire N__58090;
    wire N__58087;
    wire N__58086;
    wire N__58085;
    wire N__58082;
    wire N__58077;
    wire N__58072;
    wire N__58069;
    wire N__58066;
    wire N__58063;
    wire N__58060;
    wire N__58057;
    wire N__58054;
    wire N__58051;
    wire N__58048;
    wire N__58045;
    wire N__58042;
    wire N__58039;
    wire N__58036;
    wire N__58035;
    wire N__58034;
    wire N__58033;
    wire N__58030;
    wire N__58029;
    wire N__58028;
    wire N__58025;
    wire N__58020;
    wire N__58017;
    wire N__58016;
    wire N__58013;
    wire N__58012;
    wire N__58011;
    wire N__58008;
    wire N__58003;
    wire N__58000;
    wire N__57997;
    wire N__57994;
    wire N__57991;
    wire N__57988;
    wire N__57983;
    wire N__57980;
    wire N__57977;
    wire N__57968;
    wire N__57965;
    wire N__57962;
    wire N__57959;
    wire N__57952;
    wire N__57949;
    wire N__57948;
    wire N__57947;
    wire N__57946;
    wire N__57943;
    wire N__57942;
    wire N__57941;
    wire N__57940;
    wire N__57939;
    wire N__57938;
    wire N__57935;
    wire N__57932;
    wire N__57929;
    wire N__57926;
    wire N__57921;
    wire N__57918;
    wire N__57915;
    wire N__57912;
    wire N__57907;
    wire N__57902;
    wire N__57899;
    wire N__57896;
    wire N__57885;
    wire N__57882;
    wire N__57879;
    wire N__57874;
    wire N__57873;
    wire N__57872;
    wire N__57871;
    wire N__57870;
    wire N__57869;
    wire N__57868;
    wire N__57865;
    wire N__57862;
    wire N__57859;
    wire N__57856;
    wire N__57853;
    wire N__57850;
    wire N__57847;
    wire N__57844;
    wire N__57837;
    wire N__57834;
    wire N__57825;
    wire N__57822;
    wire N__57819;
    wire N__57814;
    wire N__57813;
    wire N__57810;
    wire N__57807;
    wire N__57804;
    wire N__57801;
    wire N__57798;
    wire N__57793;
    wire N__57792;
    wire N__57791;
    wire N__57790;
    wire N__57789;
    wire N__57786;
    wire N__57785;
    wire N__57782;
    wire N__57781;
    wire N__57778;
    wire N__57775;
    wire N__57772;
    wire N__57769;
    wire N__57766;
    wire N__57763;
    wire N__57760;
    wire N__57751;
    wire N__57748;
    wire N__57743;
    wire N__57740;
    wire N__57733;
    wire N__57730;
    wire N__57727;
    wire N__57724;
    wire N__57723;
    wire N__57722;
    wire N__57721;
    wire N__57718;
    wire N__57715;
    wire N__57712;
    wire N__57711;
    wire N__57710;
    wire N__57709;
    wire N__57708;
    wire N__57707;
    wire N__57704;
    wire N__57697;
    wire N__57694;
    wire N__57689;
    wire N__57684;
    wire N__57681;
    wire N__57678;
    wire N__57669;
    wire N__57664;
    wire N__57661;
    wire N__57658;
    wire N__57655;
    wire N__57652;
    wire N__57649;
    wire N__57648;
    wire N__57645;
    wire N__57642;
    wire N__57641;
    wire N__57636;
    wire N__57633;
    wire N__57630;
    wire N__57627;
    wire N__57624;
    wire N__57621;
    wire N__57616;
    wire N__57613;
    wire N__57612;
    wire N__57611;
    wire N__57610;
    wire N__57607;
    wire N__57604;
    wire N__57599;
    wire N__57596;
    wire N__57591;
    wire N__57588;
    wire N__57585;
    wire N__57580;
    wire N__57577;
    wire N__57574;
    wire N__57571;
    wire N__57568;
    wire N__57565;
    wire N__57562;
    wire N__57559;
    wire N__57558;
    wire N__57557;
    wire N__57554;
    wire N__57549;
    wire N__57544;
    wire N__57541;
    wire N__57538;
    wire N__57535;
    wire N__57532;
    wire N__57529;
    wire N__57526;
    wire N__57523;
    wire N__57520;
    wire N__57517;
    wire N__57516;
    wire N__57513;
    wire N__57510;
    wire N__57509;
    wire N__57504;
    wire N__57501;
    wire N__57498;
    wire N__57495;
    wire N__57490;
    wire N__57489;
    wire N__57486;
    wire N__57485;
    wire N__57482;
    wire N__57479;
    wire N__57478;
    wire N__57475;
    wire N__57472;
    wire N__57469;
    wire N__57466;
    wire N__57463;
    wire N__57460;
    wire N__57457;
    wire N__57454;
    wire N__57451;
    wire N__57448;
    wire N__57443;
    wire N__57436;
    wire N__57433;
    wire N__57430;
    wire N__57427;
    wire N__57424;
    wire N__57421;
    wire N__57418;
    wire N__57415;
    wire N__57414;
    wire N__57413;
    wire N__57412;
    wire N__57409;
    wire N__57406;
    wire N__57403;
    wire N__57400;
    wire N__57399;
    wire N__57396;
    wire N__57393;
    wire N__57390;
    wire N__57387;
    wire N__57384;
    wire N__57379;
    wire N__57374;
    wire N__57371;
    wire N__57368;
    wire N__57365;
    wire N__57362;
    wire N__57359;
    wire N__57356;
    wire N__57349;
    wire N__57346;
    wire N__57343;
    wire N__57340;
    wire N__57337;
    wire N__57334;
    wire N__57331;
    wire N__57328;
    wire N__57327;
    wire N__57326;
    wire N__57325;
    wire N__57322;
    wire N__57321;
    wire N__57320;
    wire N__57319;
    wire N__57318;
    wire N__57317;
    wire N__57314;
    wire N__57311;
    wire N__57308;
    wire N__57305;
    wire N__57300;
    wire N__57297;
    wire N__57294;
    wire N__57291;
    wire N__57288;
    wire N__57279;
    wire N__57276;
    wire N__57267;
    wire N__57264;
    wire N__57261;
    wire N__57256;
    wire N__57253;
    wire N__57250;
    wire N__57249;
    wire N__57248;
    wire N__57245;
    wire N__57244;
    wire N__57243;
    wire N__57242;
    wire N__57239;
    wire N__57236;
    wire N__57233;
    wire N__57230;
    wire N__57227;
    wire N__57226;
    wire N__57223;
    wire N__57218;
    wire N__57213;
    wire N__57210;
    wire N__57207;
    wire N__57202;
    wire N__57199;
    wire N__57194;
    wire N__57191;
    wire N__57184;
    wire N__57181;
    wire N__57178;
    wire N__57175;
    wire N__57172;
    wire N__57169;
    wire N__57166;
    wire N__57163;
    wire N__57160;
    wire N__57159;
    wire N__57156;
    wire N__57155;
    wire N__57152;
    wire N__57151;
    wire N__57150;
    wire N__57149;
    wire N__57148;
    wire N__57147;
    wire N__57144;
    wire N__57141;
    wire N__57138;
    wire N__57137;
    wire N__57134;
    wire N__57131;
    wire N__57128;
    wire N__57125;
    wire N__57122;
    wire N__57115;
    wire N__57112;
    wire N__57109;
    wire N__57106;
    wire N__57097;
    wire N__57088;
    wire N__57085;
    wire N__57082;
    wire N__57079;
    wire N__57076;
    wire N__57073;
    wire N__57072;
    wire N__57069;
    wire N__57066;
    wire N__57063;
    wire N__57060;
    wire N__57057;
    wire N__57052;
    wire N__57049;
    wire N__57046;
    wire N__57043;
    wire N__57040;
    wire N__57037;
    wire N__57034;
    wire N__57031;
    wire N__57028;
    wire N__57025;
    wire N__57022;
    wire N__57019;
    wire N__57016;
    wire N__57013;
    wire N__57010;
    wire N__57007;
    wire N__57004;
    wire N__57003;
    wire N__57000;
    wire N__56997;
    wire N__56992;
    wire N__56991;
    wire N__56988;
    wire N__56985;
    wire N__56982;
    wire N__56979;
    wire N__56974;
    wire N__56971;
    wire N__56968;
    wire N__56965;
    wire N__56962;
    wire N__56959;
    wire N__56956;
    wire N__56953;
    wire N__56950;
    wire N__56949;
    wire N__56946;
    wire N__56943;
    wire N__56938;
    wire N__56935;
    wire N__56932;
    wire N__56929;
    wire N__56926;
    wire N__56923;
    wire N__56920;
    wire N__56917;
    wire N__56914;
    wire N__56911;
    wire N__56908;
    wire N__56907;
    wire N__56906;
    wire N__56905;
    wire N__56904;
    wire N__56903;
    wire N__56902;
    wire N__56901;
    wire N__56884;
    wire N__56881;
    wire N__56878;
    wire N__56877;
    wire N__56876;
    wire N__56873;
    wire N__56870;
    wire N__56869;
    wire N__56868;
    wire N__56867;
    wire N__56866;
    wire N__56863;
    wire N__56862;
    wire N__56859;
    wire N__56856;
    wire N__56855;
    wire N__56854;
    wire N__56853;
    wire N__56852;
    wire N__56849;
    wire N__56846;
    wire N__56843;
    wire N__56840;
    wire N__56837;
    wire N__56834;
    wire N__56831;
    wire N__56828;
    wire N__56827;
    wire N__56810;
    wire N__56805;
    wire N__56802;
    wire N__56799;
    wire N__56798;
    wire N__56795;
    wire N__56792;
    wire N__56789;
    wire N__56784;
    wire N__56781;
    wire N__56770;
    wire N__56769;
    wire N__56766;
    wire N__56763;
    wire N__56760;
    wire N__56757;
    wire N__56756;
    wire N__56751;
    wire N__56748;
    wire N__56743;
    wire N__56740;
    wire N__56737;
    wire N__56734;
    wire N__56731;
    wire N__56728;
    wire N__56727;
    wire N__56724;
    wire N__56721;
    wire N__56716;
    wire N__56715;
    wire N__56712;
    wire N__56709;
    wire N__56706;
    wire N__56703;
    wire N__56698;
    wire N__56695;
    wire N__56694;
    wire N__56691;
    wire N__56688;
    wire N__56683;
    wire N__56682;
    wire N__56679;
    wire N__56676;
    wire N__56673;
    wire N__56670;
    wire N__56665;
    wire N__56662;
    wire N__56661;
    wire N__56658;
    wire N__56655;
    wire N__56650;
    wire N__56649;
    wire N__56646;
    wire N__56643;
    wire N__56640;
    wire N__56637;
    wire N__56632;
    wire N__56631;
    wire N__56630;
    wire N__56623;
    wire N__56622;
    wire N__56621;
    wire N__56620;
    wire N__56617;
    wire N__56612;
    wire N__56611;
    wire N__56610;
    wire N__56607;
    wire N__56606;
    wire N__56601;
    wire N__56596;
    wire N__56595;
    wire N__56594;
    wire N__56589;
    wire N__56586;
    wire N__56583;
    wire N__56578;
    wire N__56569;
    wire N__56566;
    wire N__56565;
    wire N__56564;
    wire N__56557;
    wire N__56556;
    wire N__56555;
    wire N__56554;
    wire N__56551;
    wire N__56546;
    wire N__56545;
    wire N__56544;
    wire N__56543;
    wire N__56540;
    wire N__56539;
    wire N__56534;
    wire N__56529;
    wire N__56526;
    wire N__56521;
    wire N__56518;
    wire N__56515;
    wire N__56512;
    wire N__56503;
    wire N__56502;
    wire N__56501;
    wire N__56494;
    wire N__56493;
    wire N__56492;
    wire N__56491;
    wire N__56488;
    wire N__56483;
    wire N__56480;
    wire N__56479;
    wire N__56478;
    wire N__56473;
    wire N__56468;
    wire N__56467;
    wire N__56464;
    wire N__56461;
    wire N__56458;
    wire N__56455;
    wire N__56446;
    wire N__56443;
    wire N__56440;
    wire N__56437;
    wire N__56434;
    wire N__56431;
    wire N__56428;
    wire N__56425;
    wire N__56422;
    wire N__56419;
    wire N__56416;
    wire N__56413;
    wire N__56410;
    wire N__56407;
    wire N__56404;
    wire N__56401;
    wire N__56398;
    wire N__56395;
    wire N__56394;
    wire N__56391;
    wire N__56388;
    wire N__56383;
    wire N__56380;
    wire N__56377;
    wire N__56374;
    wire N__56373;
    wire N__56368;
    wire N__56365;
    wire N__56362;
    wire N__56359;
    wire N__56356;
    wire N__56353;
    wire N__56350;
    wire N__56347;
    wire N__56344;
    wire N__56341;
    wire N__56338;
    wire N__56335;
    wire N__56332;
    wire N__56329;
    wire N__56326;
    wire N__56325;
    wire N__56324;
    wire N__56323;
    wire N__56320;
    wire N__56317;
    wire N__56316;
    wire N__56313;
    wire N__56310;
    wire N__56309;
    wire N__56308;
    wire N__56307;
    wire N__56306;
    wire N__56305;
    wire N__56304;
    wire N__56303;
    wire N__56302;
    wire N__56301;
    wire N__56300;
    wire N__56299;
    wire N__56298;
    wire N__56297;
    wire N__56284;
    wire N__56275;
    wire N__56274;
    wire N__56271;
    wire N__56270;
    wire N__56269;
    wire N__56262;
    wire N__56255;
    wire N__56252;
    wire N__56251;
    wire N__56246;
    wire N__56243;
    wire N__56242;
    wire N__56241;
    wire N__56240;
    wire N__56239;
    wire N__56238;
    wire N__56237;
    wire N__56236;
    wire N__56233;
    wire N__56228;
    wire N__56225;
    wire N__56220;
    wire N__56217;
    wire N__56216;
    wire N__56215;
    wire N__56212;
    wire N__56209;
    wire N__56206;
    wire N__56193;
    wire N__56190;
    wire N__56185;
    wire N__56182;
    wire N__56175;
    wire N__56172;
    wire N__56169;
    wire N__56152;
    wire N__56149;
    wire N__56146;
    wire N__56143;
    wire N__56140;
    wire N__56137;
    wire N__56134;
    wire N__56131;
    wire N__56128;
    wire N__56125;
    wire N__56122;
    wire N__56119;
    wire N__56116;
    wire N__56113;
    wire N__56110;
    wire N__56107;
    wire N__56104;
    wire N__56101;
    wire N__56100;
    wire N__56097;
    wire N__56094;
    wire N__56089;
    wire N__56086;
    wire N__56083;
    wire N__56080;
    wire N__56077;
    wire N__56074;
    wire N__56071;
    wire N__56068;
    wire N__56065;
    wire N__56062;
    wire N__56059;
    wire N__56056;
    wire N__56055;
    wire N__56052;
    wire N__56049;
    wire N__56044;
    wire N__56041;
    wire N__56038;
    wire N__56035;
    wire N__56032;
    wire N__56031;
    wire N__56028;
    wire N__56025;
    wire N__56022;
    wire N__56019;
    wire N__56016;
    wire N__56013;
    wire N__56008;
    wire N__56005;
    wire N__56004;
    wire N__56001;
    wire N__55998;
    wire N__55995;
    wire N__55992;
    wire N__55989;
    wire N__55986;
    wire N__55981;
    wire N__55978;
    wire N__55975;
    wire N__55972;
    wire N__55969;
    wire N__55966;
    wire N__55963;
    wire N__55960;
    wire N__55957;
    wire N__55954;
    wire N__55951;
    wire N__55950;
    wire N__55947;
    wire N__55944;
    wire N__55939;
    wire N__55936;
    wire N__55935;
    wire N__55930;
    wire N__55927;
    wire N__55926;
    wire N__55923;
    wire N__55920;
    wire N__55917;
    wire N__55914;
    wire N__55909;
    wire N__55906;
    wire N__55903;
    wire N__55900;
    wire N__55897;
    wire N__55894;
    wire N__55893;
    wire N__55890;
    wire N__55887;
    wire N__55884;
    wire N__55881;
    wire N__55878;
    wire N__55875;
    wire N__55872;
    wire N__55869;
    wire N__55866;
    wire N__55863;
    wire N__55860;
    wire N__55855;
    wire N__55852;
    wire N__55851;
    wire N__55848;
    wire N__55845;
    wire N__55842;
    wire N__55839;
    wire N__55834;
    wire N__55831;
    wire N__55828;
    wire N__55827;
    wire N__55824;
    wire N__55821;
    wire N__55818;
    wire N__55815;
    wire N__55812;
    wire N__55807;
    wire N__55804;
    wire N__55801;
    wire N__55798;
    wire N__55795;
    wire N__55794;
    wire N__55793;
    wire N__55792;
    wire N__55789;
    wire N__55782;
    wire N__55777;
    wire N__55774;
    wire N__55771;
    wire N__55768;
    wire N__55765;
    wire N__55764;
    wire N__55761;
    wire N__55758;
    wire N__55753;
    wire N__55750;
    wire N__55747;
    wire N__55744;
    wire N__55743;
    wire N__55740;
    wire N__55737;
    wire N__55734;
    wire N__55731;
    wire N__55728;
    wire N__55725;
    wire N__55722;
    wire N__55719;
    wire N__55714;
    wire N__55713;
    wire N__55708;
    wire N__55705;
    wire N__55702;
    wire N__55701;
    wire N__55698;
    wire N__55695;
    wire N__55692;
    wire N__55689;
    wire N__55686;
    wire N__55683;
    wire N__55680;
    wire N__55677;
    wire N__55674;
    wire N__55671;
    wire N__55668;
    wire N__55665;
    wire N__55660;
    wire N__55657;
    wire N__55654;
    wire N__55651;
    wire N__55650;
    wire N__55645;
    wire N__55642;
    wire N__55639;
    wire N__55638;
    wire N__55635;
    wire N__55634;
    wire N__55627;
    wire N__55624;
    wire N__55621;
    wire N__55620;
    wire N__55615;
    wire N__55612;
    wire N__55609;
    wire N__55606;
    wire N__55603;
    wire N__55600;
    wire N__55597;
    wire N__55594;
    wire N__55591;
    wire N__55588;
    wire N__55585;
    wire N__55582;
    wire N__55581;
    wire N__55576;
    wire N__55573;
    wire N__55570;
    wire N__55567;
    wire N__55564;
    wire N__55561;
    wire N__55558;
    wire N__55557;
    wire N__55554;
    wire N__55551;
    wire N__55548;
    wire N__55545;
    wire N__55540;
    wire N__55537;
    wire N__55534;
    wire N__55533;
    wire N__55530;
    wire N__55527;
    wire N__55522;
    wire N__55519;
    wire N__55516;
    wire N__55513;
    wire N__55510;
    wire N__55507;
    wire N__55504;
    wire N__55501;
    wire N__55498;
    wire N__55495;
    wire N__55492;
    wire N__55489;
    wire N__55486;
    wire N__55483;
    wire N__55480;
    wire N__55477;
    wire N__55474;
    wire N__55471;
    wire N__55468;
    wire N__55465;
    wire N__55462;
    wire N__55459;
    wire N__55456;
    wire N__55453;
    wire N__55450;
    wire N__55447;
    wire N__55444;
    wire N__55441;
    wire N__55438;
    wire N__55435;
    wire N__55432;
    wire N__55429;
    wire N__55426;
    wire N__55423;
    wire N__55420;
    wire N__55417;
    wire N__55414;
    wire N__55411;
    wire N__55408;
    wire N__55405;
    wire N__55402;
    wire N__55399;
    wire N__55396;
    wire N__55393;
    wire N__55390;
    wire N__55387;
    wire N__55384;
    wire N__55381;
    wire N__55378;
    wire N__55375;
    wire N__55372;
    wire N__55369;
    wire N__55366;
    wire N__55363;
    wire N__55360;
    wire N__55357;
    wire N__55354;
    wire N__55351;
    wire N__55348;
    wire N__55345;
    wire N__55342;
    wire N__55339;
    wire N__55336;
    wire N__55333;
    wire N__55330;
    wire N__55327;
    wire N__55324;
    wire N__55321;
    wire N__55318;
    wire N__55315;
    wire N__55312;
    wire N__55309;
    wire N__55306;
    wire N__55303;
    wire N__55300;
    wire N__55297;
    wire N__55294;
    wire N__55291;
    wire N__55288;
    wire N__55285;
    wire N__55282;
    wire N__55281;
    wire N__55280;
    wire N__55279;
    wire N__55278;
    wire N__55273;
    wire N__55270;
    wire N__55269;
    wire N__55268;
    wire N__55267;
    wire N__55264;
    wire N__55263;
    wire N__55262;
    wire N__55259;
    wire N__55258;
    wire N__55257;
    wire N__55256;
    wire N__55255;
    wire N__55254;
    wire N__55253;
    wire N__55248;
    wire N__55247;
    wire N__55244;
    wire N__55243;
    wire N__55242;
    wire N__55241;
    wire N__55240;
    wire N__55235;
    wire N__55234;
    wire N__55231;
    wire N__55228;
    wire N__55225;
    wire N__55222;
    wire N__55219;
    wire N__55212;
    wire N__55209;
    wire N__55208;
    wire N__55207;
    wire N__55206;
    wire N__55205;
    wire N__55202;
    wire N__55199;
    wire N__55186;
    wire N__55183;
    wire N__55180;
    wire N__55175;
    wire N__55168;
    wire N__55165;
    wire N__55162;
    wire N__55159;
    wire N__55158;
    wire N__55157;
    wire N__55150;
    wire N__55147;
    wire N__55144;
    wire N__55135;
    wire N__55128;
    wire N__55121;
    wire N__55118;
    wire N__55105;
    wire N__55102;
    wire N__55101;
    wire N__55098;
    wire N__55095;
    wire N__55092;
    wire N__55089;
    wire N__55084;
    wire N__55081;
    wire N__55080;
    wire N__55077;
    wire N__55074;
    wire N__55069;
    wire N__55068;
    wire N__55065;
    wire N__55062;
    wire N__55057;
    wire N__55056;
    wire N__55053;
    wire N__55050;
    wire N__55047;
    wire N__55042;
    wire N__55041;
    wire N__55038;
    wire N__55035;
    wire N__55030;
    wire N__55029;
    wire N__55028;
    wire N__55027;
    wire N__55026;
    wire N__55019;
    wire N__55014;
    wire N__55011;
    wire N__55008;
    wire N__55005;
    wire N__55000;
    wire N__54997;
    wire N__54996;
    wire N__54993;
    wire N__54990;
    wire N__54985;
    wire N__54982;
    wire N__54979;
    wire N__54976;
    wire N__54975;
    wire N__54972;
    wire N__54969;
    wire N__54966;
    wire N__54963;
    wire N__54960;
    wire N__54957;
    wire N__54952;
    wire N__54949;
    wire N__54946;
    wire N__54945;
    wire N__54942;
    wire N__54941;
    wire N__54940;
    wire N__54937;
    wire N__54936;
    wire N__54931;
    wire N__54924;
    wire N__54919;
    wire N__54918;
    wire N__54917;
    wire N__54916;
    wire N__54913;
    wire N__54908;
    wire N__54905;
    wire N__54898;
    wire N__54897;
    wire N__54894;
    wire N__54891;
    wire N__54888;
    wire N__54883;
    wire N__54882;
    wire N__54879;
    wire N__54876;
    wire N__54871;
    wire N__54868;
    wire N__54865;
    wire N__54864;
    wire N__54861;
    wire N__54858;
    wire N__54855;
    wire N__54850;
    wire N__54849;
    wire N__54846;
    wire N__54843;
    wire N__54840;
    wire N__54835;
    wire N__54832;
    wire N__54829;
    wire N__54826;
    wire N__54823;
    wire N__54822;
    wire N__54819;
    wire N__54816;
    wire N__54815;
    wire N__54814;
    wire N__54813;
    wire N__54812;
    wire N__54807;
    wire N__54802;
    wire N__54799;
    wire N__54796;
    wire N__54793;
    wire N__54784;
    wire N__54783;
    wire N__54782;
    wire N__54779;
    wire N__54776;
    wire N__54775;
    wire N__54774;
    wire N__54773;
    wire N__54772;
    wire N__54769;
    wire N__54764;
    wire N__54757;
    wire N__54756;
    wire N__54755;
    wire N__54752;
    wire N__54749;
    wire N__54744;
    wire N__54739;
    wire N__54730;
    wire N__54727;
    wire N__54724;
    wire N__54723;
    wire N__54720;
    wire N__54717;
    wire N__54712;
    wire N__54709;
    wire N__54706;
    wire N__54703;
    wire N__54700;
    wire N__54699;
    wire N__54696;
    wire N__54693;
    wire N__54688;
    wire N__54685;
    wire N__54682;
    wire N__54679;
    wire N__54676;
    wire N__54673;
    wire N__54672;
    wire N__54671;
    wire N__54668;
    wire N__54665;
    wire N__54662;
    wire N__54657;
    wire N__54654;
    wire N__54651;
    wire N__54646;
    wire N__54643;
    wire N__54642;
    wire N__54641;
    wire N__54638;
    wire N__54635;
    wire N__54632;
    wire N__54629;
    wire N__54626;
    wire N__54623;
    wire N__54618;
    wire N__54613;
    wire N__54610;
    wire N__54607;
    wire N__54604;
    wire N__54603;
    wire N__54602;
    wire N__54599;
    wire N__54596;
    wire N__54593;
    wire N__54590;
    wire N__54587;
    wire N__54584;
    wire N__54581;
    wire N__54578;
    wire N__54571;
    wire N__54570;
    wire N__54569;
    wire N__54566;
    wire N__54563;
    wire N__54560;
    wire N__54555;
    wire N__54552;
    wire N__54549;
    wire N__54544;
    wire N__54543;
    wire N__54540;
    wire N__54537;
    wire N__54536;
    wire N__54533;
    wire N__54530;
    wire N__54527;
    wire N__54524;
    wire N__54521;
    wire N__54514;
    wire N__54511;
    wire N__54510;
    wire N__54509;
    wire N__54506;
    wire N__54503;
    wire N__54500;
    wire N__54495;
    wire N__54492;
    wire N__54489;
    wire N__54484;
    wire N__54483;
    wire N__54480;
    wire N__54477;
    wire N__54474;
    wire N__54473;
    wire N__54470;
    wire N__54467;
    wire N__54464;
    wire N__54461;
    wire N__54458;
    wire N__54451;
    wire N__54448;
    wire N__54447;
    wire N__54444;
    wire N__54441;
    wire N__54438;
    wire N__54437;
    wire N__54434;
    wire N__54431;
    wire N__54428;
    wire N__54425;
    wire N__54422;
    wire N__54415;
    wire N__54414;
    wire N__54411;
    wire N__54410;
    wire N__54407;
    wire N__54404;
    wire N__54401;
    wire N__54398;
    wire N__54395;
    wire N__54390;
    wire N__54385;
    wire N__54384;
    wire N__54381;
    wire N__54378;
    wire N__54375;
    wire N__54374;
    wire N__54371;
    wire N__54368;
    wire N__54365;
    wire N__54362;
    wire N__54359;
    wire N__54354;
    wire N__54349;
    wire N__54348;
    wire N__54345;
    wire N__54342;
    wire N__54341;
    wire N__54338;
    wire N__54335;
    wire N__54332;
    wire N__54329;
    wire N__54326;
    wire N__54319;
    wire N__54316;
    wire N__54315;
    wire N__54312;
    wire N__54311;
    wire N__54308;
    wire N__54305;
    wire N__54302;
    wire N__54299;
    wire N__54296;
    wire N__54289;
    wire N__54288;
    wire N__54287;
    wire N__54284;
    wire N__54281;
    wire N__54278;
    wire N__54275;
    wire N__54272;
    wire N__54269;
    wire N__54262;
    wire N__54261;
    wire N__54260;
    wire N__54259;
    wire N__54256;
    wire N__54255;
    wire N__54252;
    wire N__54251;
    wire N__54250;
    wire N__54249;
    wire N__54246;
    wire N__54245;
    wire N__54242;
    wire N__54239;
    wire N__54238;
    wire N__54235;
    wire N__54232;
    wire N__54231;
    wire N__54228;
    wire N__54227;
    wire N__54222;
    wire N__54219;
    wire N__54216;
    wire N__54213;
    wire N__54210;
    wire N__54207;
    wire N__54204;
    wire N__54201;
    wire N__54196;
    wire N__54195;
    wire N__54194;
    wire N__54193;
    wire N__54190;
    wire N__54187;
    wire N__54182;
    wire N__54179;
    wire N__54176;
    wire N__54173;
    wire N__54166;
    wire N__54165;
    wire N__54164;
    wire N__54163;
    wire N__54162;
    wire N__54159;
    wire N__54156;
    wire N__54151;
    wire N__54144;
    wire N__54137;
    wire N__54128;
    wire N__54115;
    wire N__54114;
    wire N__54111;
    wire N__54110;
    wire N__54109;
    wire N__54108;
    wire N__54107;
    wire N__54106;
    wire N__54103;
    wire N__54102;
    wire N__54099;
    wire N__54096;
    wire N__54093;
    wire N__54090;
    wire N__54085;
    wire N__54082;
    wire N__54079;
    wire N__54078;
    wire N__54077;
    wire N__54076;
    wire N__54075;
    wire N__54074;
    wire N__54071;
    wire N__54068;
    wire N__54065;
    wire N__54060;
    wire N__54057;
    wire N__54054;
    wire N__54051;
    wire N__54050;
    wire N__54049;
    wire N__54048;
    wire N__54047;
    wire N__54042;
    wire N__54037;
    wire N__54034;
    wire N__54031;
    wire N__54026;
    wire N__54019;
    wire N__54010;
    wire N__53995;
    wire N__53992;
    wire N__53989;
    wire N__53986;
    wire N__53985;
    wire N__53984;
    wire N__53983;
    wire N__53980;
    wire N__53979;
    wire N__53976;
    wire N__53975;
    wire N__53974;
    wire N__53973;
    wire N__53970;
    wire N__53967;
    wire N__53964;
    wire N__53961;
    wire N__53958;
    wire N__53955;
    wire N__53952;
    wire N__53945;
    wire N__53932;
    wire N__53931;
    wire N__53928;
    wire N__53925;
    wire N__53922;
    wire N__53917;
    wire N__53914;
    wire N__53911;
    wire N__53908;
    wire N__53907;
    wire N__53904;
    wire N__53901;
    wire N__53896;
    wire N__53893;
    wire N__53890;
    wire N__53887;
    wire N__53886;
    wire N__53883;
    wire N__53880;
    wire N__53877;
    wire N__53874;
    wire N__53871;
    wire N__53868;
    wire N__53865;
    wire N__53862;
    wire N__53859;
    wire N__53856;
    wire N__53851;
    wire N__53848;
    wire N__53845;
    wire N__53842;
    wire N__53839;
    wire N__53836;
    wire N__53833;
    wire N__53830;
    wire N__53827;
    wire N__53824;
    wire N__53821;
    wire N__53818;
    wire N__53815;
    wire N__53812;
    wire N__53809;
    wire N__53808;
    wire N__53807;
    wire N__53806;
    wire N__53805;
    wire N__53802;
    wire N__53799;
    wire N__53798;
    wire N__53797;
    wire N__53796;
    wire N__53795;
    wire N__53794;
    wire N__53793;
    wire N__53790;
    wire N__53789;
    wire N__53788;
    wire N__53787;
    wire N__53782;
    wire N__53781;
    wire N__53780;
    wire N__53779;
    wire N__53776;
    wire N__53773;
    wire N__53772;
    wire N__53771;
    wire N__53768;
    wire N__53761;
    wire N__53754;
    wire N__53747;
    wire N__53744;
    wire N__53741;
    wire N__53736;
    wire N__53731;
    wire N__53726;
    wire N__53721;
    wire N__53716;
    wire N__53709;
    wire N__53698;
    wire N__53697;
    wire N__53696;
    wire N__53695;
    wire N__53694;
    wire N__53693;
    wire N__53692;
    wire N__53691;
    wire N__53690;
    wire N__53687;
    wire N__53686;
    wire N__53683;
    wire N__53682;
    wire N__53681;
    wire N__53680;
    wire N__53679;
    wire N__53676;
    wire N__53673;
    wire N__53666;
    wire N__53661;
    wire N__53660;
    wire N__53657;
    wire N__53656;
    wire N__53653;
    wire N__53648;
    wire N__53645;
    wire N__53644;
    wire N__53643;
    wire N__53640;
    wire N__53639;
    wire N__53638;
    wire N__53635;
    wire N__53630;
    wire N__53627;
    wire N__53626;
    wire N__53625;
    wire N__53622;
    wire N__53619;
    wire N__53616;
    wire N__53613;
    wire N__53610;
    wire N__53607;
    wire N__53600;
    wire N__53593;
    wire N__53586;
    wire N__53581;
    wire N__53576;
    wire N__53557;
    wire N__53554;
    wire N__53551;
    wire N__53550;
    wire N__53547;
    wire N__53544;
    wire N__53541;
    wire N__53538;
    wire N__53533;
    wire N__53530;
    wire N__53527;
    wire N__53524;
    wire N__53521;
    wire N__53520;
    wire N__53519;
    wire N__53518;
    wire N__53517;
    wire N__53508;
    wire N__53507;
    wire N__53504;
    wire N__53503;
    wire N__53502;
    wire N__53501;
    wire N__53498;
    wire N__53495;
    wire N__53492;
    wire N__53485;
    wire N__53482;
    wire N__53473;
    wire N__53470;
    wire N__53467;
    wire N__53464;
    wire N__53461;
    wire N__53458;
    wire N__53455;
    wire N__53454;
    wire N__53451;
    wire N__53448;
    wire N__53445;
    wire N__53442;
    wire N__53441;
    wire N__53436;
    wire N__53433;
    wire N__53430;
    wire N__53425;
    wire N__53422;
    wire N__53421;
    wire N__53418;
    wire N__53417;
    wire N__53414;
    wire N__53411;
    wire N__53408;
    wire N__53401;
    wire N__53398;
    wire N__53397;
    wire N__53394;
    wire N__53391;
    wire N__53390;
    wire N__53387;
    wire N__53384;
    wire N__53381;
    wire N__53378;
    wire N__53375;
    wire N__53368;
    wire N__53365;
    wire N__53364;
    wire N__53361;
    wire N__53360;
    wire N__53357;
    wire N__53354;
    wire N__53351;
    wire N__53348;
    wire N__53345;
    wire N__53338;
    wire N__53335;
    wire N__53334;
    wire N__53333;
    wire N__53328;
    wire N__53325;
    wire N__53322;
    wire N__53317;
    wire N__53314;
    wire N__53313;
    wire N__53312;
    wire N__53307;
    wire N__53304;
    wire N__53301;
    wire N__53296;
    wire N__53293;
    wire N__53292;
    wire N__53289;
    wire N__53286;
    wire N__53285;
    wire N__53282;
    wire N__53279;
    wire N__53276;
    wire N__53271;
    wire N__53266;
    wire N__53263;
    wire N__53262;
    wire N__53259;
    wire N__53256;
    wire N__53255;
    wire N__53252;
    wire N__53249;
    wire N__53246;
    wire N__53243;
    wire N__53240;
    wire N__53233;
    wire N__53230;
    wire N__53227;
    wire N__53226;
    wire N__53225;
    wire N__53224;
    wire N__53221;
    wire N__53218;
    wire N__53213;
    wire N__53210;
    wire N__53203;
    wire N__53202;
    wire N__53201;
    wire N__53198;
    wire N__53195;
    wire N__53192;
    wire N__53185;
    wire N__53184;
    wire N__53181;
    wire N__53178;
    wire N__53175;
    wire N__53172;
    wire N__53169;
    wire N__53166;
    wire N__53163;
    wire N__53158;
    wire N__53155;
    wire N__53154;
    wire N__53153;
    wire N__53150;
    wire N__53147;
    wire N__53144;
    wire N__53141;
    wire N__53134;
    wire N__53131;
    wire N__53130;
    wire N__53129;
    wire N__53126;
    wire N__53123;
    wire N__53120;
    wire N__53113;
    wire N__53110;
    wire N__53109;
    wire N__53108;
    wire N__53105;
    wire N__53102;
    wire N__53099;
    wire N__53092;
    wire N__53089;
    wire N__53088;
    wire N__53087;
    wire N__53084;
    wire N__53081;
    wire N__53078;
    wire N__53071;
    wire N__53068;
    wire N__53067;
    wire N__53066;
    wire N__53063;
    wire N__53060;
    wire N__53057;
    wire N__53054;
    wire N__53051;
    wire N__53044;
    wire N__53041;
    wire N__53040;
    wire N__53037;
    wire N__53036;
    wire N__53033;
    wire N__53030;
    wire N__53027;
    wire N__53020;
    wire N__53017;
    wire N__53016;
    wire N__53013;
    wire N__53012;
    wire N__53009;
    wire N__53006;
    wire N__53003;
    wire N__52996;
    wire N__52993;
    wire N__52992;
    wire N__52989;
    wire N__52988;
    wire N__52985;
    wire N__52982;
    wire N__52979;
    wire N__52972;
    wire N__52969;
    wire N__52966;
    wire N__52963;
    wire N__52960;
    wire N__52957;
    wire N__52954;
    wire N__52951;
    wire N__52948;
    wire N__52945;
    wire N__52942;
    wire N__52939;
    wire N__52938;
    wire N__52933;
    wire N__52930;
    wire N__52927;
    wire N__52924;
    wire N__52921;
    wire N__52918;
    wire N__52915;
    wire N__52912;
    wire N__52909;
    wire N__52906;
    wire N__52905;
    wire N__52902;
    wire N__52901;
    wire N__52900;
    wire N__52899;
    wire N__52896;
    wire N__52895;
    wire N__52894;
    wire N__52893;
    wire N__52892;
    wire N__52891;
    wire N__52890;
    wire N__52889;
    wire N__52888;
    wire N__52887;
    wire N__52886;
    wire N__52885;
    wire N__52884;
    wire N__52883;
    wire N__52882;
    wire N__52881;
    wire N__52880;
    wire N__52879;
    wire N__52878;
    wire N__52877;
    wire N__52874;
    wire N__52869;
    wire N__52868;
    wire N__52867;
    wire N__52866;
    wire N__52865;
    wire N__52864;
    wire N__52863;
    wire N__52862;
    wire N__52861;
    wire N__52860;
    wire N__52859;
    wire N__52856;
    wire N__52853;
    wire N__52848;
    wire N__52841;
    wire N__52838;
    wire N__52833;
    wire N__52830;
    wire N__52825;
    wire N__52818;
    wire N__52813;
    wire N__52806;
    wire N__52805;
    wire N__52804;
    wire N__52803;
    wire N__52802;
    wire N__52801;
    wire N__52800;
    wire N__52799;
    wire N__52794;
    wire N__52791;
    wire N__52782;
    wire N__52771;
    wire N__52770;
    wire N__52769;
    wire N__52768;
    wire N__52767;
    wire N__52766;
    wire N__52765;
    wire N__52764;
    wire N__52759;
    wire N__52756;
    wire N__52743;
    wire N__52742;
    wire N__52741;
    wire N__52738;
    wire N__52735;
    wire N__52720;
    wire N__52713;
    wire N__52712;
    wire N__52711;
    wire N__52708;
    wire N__52701;
    wire N__52692;
    wire N__52685;
    wire N__52682;
    wire N__52681;
    wire N__52680;
    wire N__52679;
    wire N__52678;
    wire N__52677;
    wire N__52674;
    wire N__52671;
    wire N__52664;
    wire N__52659;
    wire N__52648;
    wire N__52637;
    wire N__52624;
    wire N__52623;
    wire N__52622;
    wire N__52619;
    wire N__52616;
    wire N__52613;
    wire N__52610;
    wire N__52603;
    wire N__52600;
    wire N__52599;
    wire N__52598;
    wire N__52595;
    wire N__52592;
    wire N__52589;
    wire N__52586;
    wire N__52579;
    wire N__52576;
    wire N__52575;
    wire N__52572;
    wire N__52571;
    wire N__52568;
    wire N__52565;
    wire N__52562;
    wire N__52557;
    wire N__52552;
    wire N__52549;
    wire N__52546;
    wire N__52543;
    wire N__52540;
    wire N__52537;
    wire N__52534;
    wire N__52533;
    wire N__52530;
    wire N__52527;
    wire N__52522;
    wire N__52519;
    wire N__52516;
    wire N__52513;
    wire N__52510;
    wire N__52507;
    wire N__52504;
    wire N__52501;
    wire N__52498;
    wire N__52495;
    wire N__52492;
    wire N__52489;
    wire N__52486;
    wire N__52483;
    wire N__52480;
    wire N__52477;
    wire N__52474;
    wire N__52471;
    wire N__52468;
    wire N__52465;
    wire N__52464;
    wire N__52463;
    wire N__52462;
    wire N__52461;
    wire N__52458;
    wire N__52457;
    wire N__52454;
    wire N__52445;
    wire N__52442;
    wire N__52439;
    wire N__52436;
    wire N__52433;
    wire N__52430;
    wire N__52423;
    wire N__52420;
    wire N__52419;
    wire N__52416;
    wire N__52413;
    wire N__52410;
    wire N__52405;
    wire N__52402;
    wire N__52401;
    wire N__52398;
    wire N__52395;
    wire N__52390;
    wire N__52387;
    wire N__52384;
    wire N__52381;
    wire N__52380;
    wire N__52375;
    wire N__52372;
    wire N__52369;
    wire N__52366;
    wire N__52363;
    wire N__52360;
    wire N__52357;
    wire N__52354;
    wire N__52351;
    wire N__52348;
    wire N__52345;
    wire N__52342;
    wire N__52339;
    wire N__52336;
    wire N__52333;
    wire N__52330;
    wire N__52329;
    wire N__52326;
    wire N__52323;
    wire N__52320;
    wire N__52317;
    wire N__52314;
    wire N__52311;
    wire N__52306;
    wire N__52303;
    wire N__52300;
    wire N__52297;
    wire N__52294;
    wire N__52291;
    wire N__52288;
    wire N__52285;
    wire N__52282;
    wire N__52279;
    wire N__52276;
    wire N__52273;
    wire N__52270;
    wire N__52267;
    wire N__52264;
    wire N__52261;
    wire N__52258;
    wire N__52255;
    wire N__52252;
    wire N__52249;
    wire N__52246;
    wire N__52243;
    wire N__52242;
    wire N__52241;
    wire N__52238;
    wire N__52237;
    wire N__52236;
    wire N__52235;
    wire N__52234;
    wire N__52231;
    wire N__52230;
    wire N__52229;
    wire N__52226;
    wire N__52225;
    wire N__52222;
    wire N__52219;
    wire N__52216;
    wire N__52213;
    wire N__52210;
    wire N__52209;
    wire N__52208;
    wire N__52207;
    wire N__52206;
    wire N__52203;
    wire N__52200;
    wire N__52197;
    wire N__52194;
    wire N__52191;
    wire N__52188;
    wire N__52185;
    wire N__52170;
    wire N__52167;
    wire N__52164;
    wire N__52157;
    wire N__52154;
    wire N__52151;
    wire N__52146;
    wire N__52141;
    wire N__52132;
    wire N__52129;
    wire N__52126;
    wire N__52125;
    wire N__52124;
    wire N__52123;
    wire N__52120;
    wire N__52113;
    wire N__52108;
    wire N__52107;
    wire N__52106;
    wire N__52105;
    wire N__52102;
    wire N__52099;
    wire N__52094;
    wire N__52091;
    wire N__52088;
    wire N__52081;
    wire N__52078;
    wire N__52075;
    wire N__52072;
    wire N__52071;
    wire N__52068;
    wire N__52065;
    wire N__52062;
    wire N__52057;
    wire N__52056;
    wire N__52053;
    wire N__52050;
    wire N__52049;
    wire N__52046;
    wire N__52045;
    wire N__52040;
    wire N__52037;
    wire N__52034;
    wire N__52027;
    wire N__52024;
    wire N__52021;
    wire N__52018;
    wire N__52017;
    wire N__52014;
    wire N__52011;
    wire N__52010;
    wire N__52007;
    wire N__52004;
    wire N__52001;
    wire N__51996;
    wire N__51991;
    wire N__51990;
    wire N__51987;
    wire N__51984;
    wire N__51981;
    wire N__51976;
    wire N__51973;
    wire N__51972;
    wire N__51969;
    wire N__51966;
    wire N__51963;
    wire N__51958;
    wire N__51955;
    wire N__51952;
    wire N__51949;
    wire N__51946;
    wire N__51943;
    wire N__51940;
    wire N__51939;
    wire N__51936;
    wire N__51933;
    wire N__51930;
    wire N__51925;
    wire N__51922;
    wire N__51919;
    wire N__51916;
    wire N__51913;
    wire N__51912;
    wire N__51909;
    wire N__51906;
    wire N__51903;
    wire N__51898;
    wire N__51895;
    wire N__51894;
    wire N__51891;
    wire N__51888;
    wire N__51885;
    wire N__51880;
    wire N__51877;
    wire N__51876;
    wire N__51873;
    wire N__51870;
    wire N__51867;
    wire N__51862;
    wire N__51859;
    wire N__51856;
    wire N__51853;
    wire N__51852;
    wire N__51849;
    wire N__51846;
    wire N__51841;
    wire N__51838;
    wire N__51835;
    wire N__51834;
    wire N__51831;
    wire N__51828;
    wire N__51825;
    wire N__51820;
    wire N__51817;
    wire N__51814;
    wire N__51811;
    wire N__51808;
    wire N__51807;
    wire N__51804;
    wire N__51801;
    wire N__51796;
    wire N__51793;
    wire N__51790;
    wire N__51787;
    wire N__51784;
    wire N__51781;
    wire N__51778;
    wire N__51777;
    wire N__51774;
    wire N__51773;
    wire N__51772;
    wire N__51765;
    wire N__51762;
    wire N__51757;
    wire N__51754;
    wire N__51753;
    wire N__51752;
    wire N__51749;
    wire N__51744;
    wire N__51741;
    wire N__51736;
    wire N__51733;
    wire N__51730;
    wire N__51729;
    wire N__51726;
    wire N__51723;
    wire N__51718;
    wire N__51715;
    wire N__51714;
    wire N__51711;
    wire N__51708;
    wire N__51703;
    wire N__51700;
    wire N__51697;
    wire N__51696;
    wire N__51693;
    wire N__51690;
    wire N__51685;
    wire N__51682;
    wire N__51681;
    wire N__51678;
    wire N__51675;
    wire N__51670;
    wire N__51667;
    wire N__51664;
    wire N__51661;
    wire N__51658;
    wire N__51655;
    wire N__51652;
    wire N__51649;
    wire N__51646;
    wire N__51643;
    wire N__51640;
    wire N__51637;
    wire N__51634;
    wire N__51631;
    wire N__51630;
    wire N__51627;
    wire N__51626;
    wire N__51623;
    wire N__51620;
    wire N__51615;
    wire N__51612;
    wire N__51607;
    wire N__51604;
    wire N__51601;
    wire N__51598;
    wire N__51595;
    wire N__51592;
    wire N__51591;
    wire N__51590;
    wire N__51589;
    wire N__51586;
    wire N__51583;
    wire N__51578;
    wire N__51575;
    wire N__51568;
    wire N__51567;
    wire N__51564;
    wire N__51563;
    wire N__51562;
    wire N__51561;
    wire N__51558;
    wire N__51555;
    wire N__51552;
    wire N__51549;
    wire N__51544;
    wire N__51539;
    wire N__51536;
    wire N__51533;
    wire N__51530;
    wire N__51527;
    wire N__51520;
    wire N__51519;
    wire N__51518;
    wire N__51515;
    wire N__51514;
    wire N__51513;
    wire N__51510;
    wire N__51509;
    wire N__51506;
    wire N__51503;
    wire N__51498;
    wire N__51497;
    wire N__51496;
    wire N__51493;
    wire N__51490;
    wire N__51483;
    wire N__51478;
    wire N__51469;
    wire N__51468;
    wire N__51463;
    wire N__51460;
    wire N__51459;
    wire N__51458;
    wire N__51455;
    wire N__51450;
    wire N__51445;
    wire N__51442;
    wire N__51441;
    wire N__51440;
    wire N__51437;
    wire N__51432;
    wire N__51427;
    wire N__51424;
    wire N__51421;
    wire N__51418;
    wire N__51415;
    wire N__51412;
    wire N__51409;
    wire N__51406;
    wire N__51403;
    wire N__51402;
    wire N__51399;
    wire N__51396;
    wire N__51393;
    wire N__51390;
    wire N__51385;
    wire N__51382;
    wire N__51379;
    wire N__51378;
    wire N__51375;
    wire N__51374;
    wire N__51373;
    wire N__51372;
    wire N__51371;
    wire N__51370;
    wire N__51369;
    wire N__51368;
    wire N__51367;
    wire N__51366;
    wire N__51365;
    wire N__51360;
    wire N__51359;
    wire N__51358;
    wire N__51357;
    wire N__51356;
    wire N__51355;
    wire N__51354;
    wire N__51353;
    wire N__51352;
    wire N__51351;
    wire N__51350;
    wire N__51347;
    wire N__51346;
    wire N__51345;
    wire N__51344;
    wire N__51341;
    wire N__51338;
    wire N__51335;
    wire N__51332;
    wire N__51329;
    wire N__51328;
    wire N__51327;
    wire N__51324;
    wire N__51323;
    wire N__51322;
    wire N__51321;
    wire N__51320;
    wire N__51319;
    wire N__51318;
    wire N__51317;
    wire N__51314;
    wire N__51311;
    wire N__51308;
    wire N__51305;
    wire N__51298;
    wire N__51297;
    wire N__51296;
    wire N__51295;
    wire N__51292;
    wire N__51289;
    wire N__51288;
    wire N__51287;
    wire N__51286;
    wire N__51285;
    wire N__51282;
    wire N__51279;
    wire N__51278;
    wire N__51275;
    wire N__51272;
    wire N__51271;
    wire N__51268;
    wire N__51267;
    wire N__51262;
    wire N__51261;
    wire N__51260;
    wire N__51259;
    wire N__51246;
    wire N__51243;
    wire N__51238;
    wire N__51235;
    wire N__51234;
    wire N__51231;
    wire N__51228;
    wire N__51225;
    wire N__51224;
    wire N__51223;
    wire N__51222;
    wire N__51219;
    wire N__51206;
    wire N__51201;
    wire N__51190;
    wire N__51177;
    wire N__51170;
    wire N__51163;
    wire N__51160;
    wire N__51155;
    wire N__51152;
    wire N__51149;
    wire N__51144;
    wire N__51141;
    wire N__51126;
    wire N__51119;
    wire N__51116;
    wire N__51113;
    wire N__51104;
    wire N__51097;
    wire N__51090;
    wire N__51087;
    wire N__51082;
    wire N__51079;
    wire N__51076;
    wire N__51067;
    wire N__51064;
    wire N__51063;
    wire N__51060;
    wire N__51057;
    wire N__51054;
    wire N__51051;
    wire N__51048;
    wire N__51043;
    wire N__51040;
    wire N__51037;
    wire N__51034;
    wire N__51031;
    wire N__51028;
    wire N__51025;
    wire N__51022;
    wire N__51019;
    wire N__51018;
    wire N__51015;
    wire N__51012;
    wire N__51007;
    wire N__51004;
    wire N__51001;
    wire N__50998;
    wire N__50995;
    wire N__50992;
    wire N__50989;
    wire N__50986;
    wire N__50985;
    wire N__50984;
    wire N__50983;
    wire N__50982;
    wire N__50981;
    wire N__50980;
    wire N__50979;
    wire N__50970;
    wire N__50961;
    wire N__50960;
    wire N__50959;
    wire N__50958;
    wire N__50957;
    wire N__50956;
    wire N__50951;
    wire N__50950;
    wire N__50949;
    wire N__50944;
    wire N__50941;
    wire N__50938;
    wire N__50935;
    wire N__50934;
    wire N__50931;
    wire N__50928;
    wire N__50925;
    wire N__50922;
    wire N__50921;
    wire N__50920;
    wire N__50915;
    wire N__50912;
    wire N__50909;
    wire N__50904;
    wire N__50899;
    wire N__50896;
    wire N__50893;
    wire N__50886;
    wire N__50881;
    wire N__50878;
    wire N__50869;
    wire N__50866;
    wire N__50863;
    wire N__50860;
    wire N__50857;
    wire N__50854;
    wire N__50851;
    wire N__50850;
    wire N__50849;
    wire N__50848;
    wire N__50845;
    wire N__50842;
    wire N__50839;
    wire N__50836;
    wire N__50833;
    wire N__50830;
    wire N__50825;
    wire N__50818;
    wire N__50815;
    wire N__50812;
    wire N__50809;
    wire N__50806;
    wire N__50803;
    wire N__50800;
    wire N__50797;
    wire N__50796;
    wire N__50793;
    wire N__50790;
    wire N__50787;
    wire N__50784;
    wire N__50783;
    wire N__50782;
    wire N__50779;
    wire N__50778;
    wire N__50775;
    wire N__50770;
    wire N__50767;
    wire N__50764;
    wire N__50755;
    wire N__50752;
    wire N__50749;
    wire N__50746;
    wire N__50743;
    wire N__50740;
    wire N__50739;
    wire N__50736;
    wire N__50733;
    wire N__50730;
    wire N__50727;
    wire N__50724;
    wire N__50721;
    wire N__50716;
    wire N__50713;
    wire N__50710;
    wire N__50707;
    wire N__50704;
    wire N__50701;
    wire N__50700;
    wire N__50697;
    wire N__50696;
    wire N__50693;
    wire N__50690;
    wire N__50687;
    wire N__50684;
    wire N__50681;
    wire N__50678;
    wire N__50671;
    wire N__50668;
    wire N__50665;
    wire N__50662;
    wire N__50659;
    wire N__50656;
    wire N__50653;
    wire N__50650;
    wire N__50647;
    wire N__50644;
    wire N__50641;
    wire N__50638;
    wire N__50637;
    wire N__50634;
    wire N__50631;
    wire N__50630;
    wire N__50627;
    wire N__50624;
    wire N__50621;
    wire N__50616;
    wire N__50611;
    wire N__50608;
    wire N__50605;
    wire N__50602;
    wire N__50599;
    wire N__50598;
    wire N__50595;
    wire N__50594;
    wire N__50591;
    wire N__50588;
    wire N__50585;
    wire N__50584;
    wire N__50583;
    wire N__50580;
    wire N__50577;
    wire N__50574;
    wire N__50571;
    wire N__50568;
    wire N__50565;
    wire N__50560;
    wire N__50559;
    wire N__50556;
    wire N__50553;
    wire N__50550;
    wire N__50547;
    wire N__50544;
    wire N__50539;
    wire N__50530;
    wire N__50529;
    wire N__50528;
    wire N__50525;
    wire N__50522;
    wire N__50519;
    wire N__50516;
    wire N__50513;
    wire N__50510;
    wire N__50507;
    wire N__50504;
    wire N__50497;
    wire N__50496;
    wire N__50495;
    wire N__50492;
    wire N__50491;
    wire N__50486;
    wire N__50483;
    wire N__50482;
    wire N__50479;
    wire N__50474;
    wire N__50469;
    wire N__50466;
    wire N__50463;
    wire N__50460;
    wire N__50457;
    wire N__50452;
    wire N__50451;
    wire N__50448;
    wire N__50445;
    wire N__50440;
    wire N__50439;
    wire N__50438;
    wire N__50437;
    wire N__50434;
    wire N__50427;
    wire N__50422;
    wire N__50419;
    wire N__50418;
    wire N__50415;
    wire N__50414;
    wire N__50411;
    wire N__50408;
    wire N__50405;
    wire N__50402;
    wire N__50399;
    wire N__50396;
    wire N__50391;
    wire N__50386;
    wire N__50385;
    wire N__50384;
    wire N__50383;
    wire N__50380;
    wire N__50379;
    wire N__50376;
    wire N__50373;
    wire N__50370;
    wire N__50367;
    wire N__50364;
    wire N__50361;
    wire N__50358;
    wire N__50355;
    wire N__50350;
    wire N__50349;
    wire N__50344;
    wire N__50341;
    wire N__50338;
    wire N__50335;
    wire N__50332;
    wire N__50327;
    wire N__50324;
    wire N__50317;
    wire N__50314;
    wire N__50311;
    wire N__50308;
    wire N__50305;
    wire N__50302;
    wire N__50299;
    wire N__50296;
    wire N__50293;
    wire N__50290;
    wire N__50287;
    wire N__50284;
    wire N__50281;
    wire N__50280;
    wire N__50277;
    wire N__50274;
    wire N__50271;
    wire N__50266;
    wire N__50263;
    wire N__50260;
    wire N__50257;
    wire N__50254;
    wire N__50251;
    wire N__50248;
    wire N__50245;
    wire N__50242;
    wire N__50241;
    wire N__50238;
    wire N__50235;
    wire N__50234;
    wire N__50231;
    wire N__50228;
    wire N__50225;
    wire N__50222;
    wire N__50219;
    wire N__50216;
    wire N__50213;
    wire N__50210;
    wire N__50203;
    wire N__50200;
    wire N__50197;
    wire N__50194;
    wire N__50191;
    wire N__50188;
    wire N__50185;
    wire N__50184;
    wire N__50181;
    wire N__50178;
    wire N__50175;
    wire N__50174;
    wire N__50171;
    wire N__50168;
    wire N__50165;
    wire N__50160;
    wire N__50157;
    wire N__50152;
    wire N__50149;
    wire N__50146;
    wire N__50143;
    wire N__50140;
    wire N__50137;
    wire N__50134;
    wire N__50131;
    wire N__50128;
    wire N__50125;
    wire N__50122;
    wire N__50119;
    wire N__50118;
    wire N__50117;
    wire N__50114;
    wire N__50111;
    wire N__50110;
    wire N__50107;
    wire N__50104;
    wire N__50101;
    wire N__50098;
    wire N__50095;
    wire N__50092;
    wire N__50089;
    wire N__50084;
    wire N__50077;
    wire N__50074;
    wire N__50071;
    wire N__50068;
    wire N__50065;
    wire N__50062;
    wire N__50059;
    wire N__50056;
    wire N__50053;
    wire N__50050;
    wire N__50047;
    wire N__50044;
    wire N__50041;
    wire N__50038;
    wire N__50035;
    wire N__50032;
    wire N__50029;
    wire N__50026;
    wire N__50023;
    wire N__50020;
    wire N__50017;
    wire N__50014;
    wire N__50013;
    wire N__50010;
    wire N__50009;
    wire N__50008;
    wire N__50005;
    wire N__50002;
    wire N__49999;
    wire N__49994;
    wire N__49989;
    wire N__49986;
    wire N__49981;
    wire N__49978;
    wire N__49975;
    wire N__49972;
    wire N__49969;
    wire N__49968;
    wire N__49967;
    wire N__49964;
    wire N__49961;
    wire N__49960;
    wire N__49957;
    wire N__49954;
    wire N__49951;
    wire N__49948;
    wire N__49945;
    wire N__49942;
    wire N__49939;
    wire N__49936;
    wire N__49933;
    wire N__49928;
    wire N__49921;
    wire N__49918;
    wire N__49915;
    wire N__49912;
    wire N__49911;
    wire N__49908;
    wire N__49905;
    wire N__49900;
    wire N__49897;
    wire N__49894;
    wire N__49891;
    wire N__49888;
    wire N__49885;
    wire N__49882;
    wire N__49879;
    wire N__49876;
    wire N__49873;
    wire N__49870;
    wire N__49867;
    wire N__49864;
    wire N__49861;
    wire N__49858;
    wire N__49855;
    wire N__49854;
    wire N__49851;
    wire N__49848;
    wire N__49845;
    wire N__49842;
    wire N__49839;
    wire N__49836;
    wire N__49831;
    wire N__49828;
    wire N__49825;
    wire N__49822;
    wire N__49819;
    wire N__49816;
    wire N__49813;
    wire N__49810;
    wire N__49809;
    wire N__49806;
    wire N__49803;
    wire N__49798;
    wire N__49797;
    wire N__49794;
    wire N__49791;
    wire N__49786;
    wire N__49783;
    wire N__49782;
    wire N__49781;
    wire N__49780;
    wire N__49779;
    wire N__49776;
    wire N__49771;
    wire N__49766;
    wire N__49765;
    wire N__49764;
    wire N__49761;
    wire N__49758;
    wire N__49755;
    wire N__49750;
    wire N__49741;
    wire N__49740;
    wire N__49737;
    wire N__49734;
    wire N__49733;
    wire N__49730;
    wire N__49727;
    wire N__49724;
    wire N__49721;
    wire N__49716;
    wire N__49713;
    wire N__49710;
    wire N__49705;
    wire N__49702;
    wire N__49701;
    wire N__49700;
    wire N__49699;
    wire N__49698;
    wire N__49697;
    wire N__49696;
    wire N__49693;
    wire N__49692;
    wire N__49691;
    wire N__49690;
    wire N__49687;
    wire N__49680;
    wire N__49677;
    wire N__49676;
    wire N__49673;
    wire N__49672;
    wire N__49669;
    wire N__49664;
    wire N__49659;
    wire N__49658;
    wire N__49657;
    wire N__49652;
    wire N__49649;
    wire N__49648;
    wire N__49647;
    wire N__49646;
    wire N__49645;
    wire N__49644;
    wire N__49643;
    wire N__49642;
    wire N__49641;
    wire N__49636;
    wire N__49629;
    wire N__49624;
    wire N__49623;
    wire N__49620;
    wire N__49615;
    wire N__49608;
    wire N__49599;
    wire N__49592;
    wire N__49589;
    wire N__49586;
    wire N__49583;
    wire N__49580;
    wire N__49575;
    wire N__49564;
    wire N__49563;
    wire N__49562;
    wire N__49555;
    wire N__49552;
    wire N__49551;
    wire N__49550;
    wire N__49549;
    wire N__49546;
    wire N__49539;
    wire N__49534;
    wire N__49533;
    wire N__49532;
    wire N__49531;
    wire N__49528;
    wire N__49523;
    wire N__49520;
    wire N__49517;
    wire N__49514;
    wire N__49511;
    wire N__49504;
    wire N__49503;
    wire N__49502;
    wire N__49501;
    wire N__49500;
    wire N__49499;
    wire N__49496;
    wire N__49495;
    wire N__49492;
    wire N__49489;
    wire N__49486;
    wire N__49483;
    wire N__49482;
    wire N__49481;
    wire N__49480;
    wire N__49477;
    wire N__49472;
    wire N__49465;
    wire N__49456;
    wire N__49455;
    wire N__49454;
    wire N__49453;
    wire N__49452;
    wire N__49451;
    wire N__49448;
    wire N__49445;
    wire N__49444;
    wire N__49443;
    wire N__49442;
    wire N__49437;
    wire N__49426;
    wire N__49421;
    wire N__49416;
    wire N__49413;
    wire N__49410;
    wire N__49405;
    wire N__49396;
    wire N__49395;
    wire N__49394;
    wire N__49391;
    wire N__49390;
    wire N__49387;
    wire N__49386;
    wire N__49385;
    wire N__49384;
    wire N__49383;
    wire N__49382;
    wire N__49381;
    wire N__49378;
    wire N__49371;
    wire N__49370;
    wire N__49369;
    wire N__49366;
    wire N__49363;
    wire N__49360;
    wire N__49357;
    wire N__49354;
    wire N__49351;
    wire N__49348;
    wire N__49345;
    wire N__49340;
    wire N__49333;
    wire N__49328;
    wire N__49325;
    wire N__49322;
    wire N__49319;
    wire N__49314;
    wire N__49309;
    wire N__49308;
    wire N__49307;
    wire N__49306;
    wire N__49305;
    wire N__49304;
    wire N__49303;
    wire N__49300;
    wire N__49293;
    wire N__49280;
    wire N__49273;
    wire N__49270;
    wire N__49267;
    wire N__49264;
    wire N__49261;
    wire N__49258;
    wire N__49255;
    wire N__49252;
    wire N__49249;
    wire N__49246;
    wire N__49245;
    wire N__49242;
    wire N__49239;
    wire N__49236;
    wire N__49233;
    wire N__49230;
    wire N__49227;
    wire N__49224;
    wire N__49219;
    wire N__49218;
    wire N__49217;
    wire N__49214;
    wire N__49211;
    wire N__49206;
    wire N__49203;
    wire N__49200;
    wire N__49197;
    wire N__49194;
    wire N__49189;
    wire N__49186;
    wire N__49183;
    wire N__49180;
    wire N__49179;
    wire N__49176;
    wire N__49173;
    wire N__49172;
    wire N__49169;
    wire N__49166;
    wire N__49163;
    wire N__49156;
    wire N__49153;
    wire N__49150;
    wire N__49147;
    wire N__49144;
    wire N__49141;
    wire N__49138;
    wire N__49137;
    wire N__49136;
    wire N__49133;
    wire N__49130;
    wire N__49127;
    wire N__49126;
    wire N__49123;
    wire N__49118;
    wire N__49115;
    wire N__49112;
    wire N__49109;
    wire N__49106;
    wire N__49099;
    wire N__49096;
    wire N__49093;
    wire N__49092;
    wire N__49089;
    wire N__49086;
    wire N__49081;
    wire N__49078;
    wire N__49075;
    wire N__49072;
    wire N__49071;
    wire N__49068;
    wire N__49065;
    wire N__49064;
    wire N__49063;
    wire N__49060;
    wire N__49055;
    wire N__49052;
    wire N__49047;
    wire N__49042;
    wire N__49039;
    wire N__49036;
    wire N__49035;
    wire N__49032;
    wire N__49029;
    wire N__49024;
    wire N__49021;
    wire N__49018;
    wire N__49015;
    wire N__49012;
    wire N__49009;
    wire N__49006;
    wire N__49005;
    wire N__49004;
    wire N__49001;
    wire N__48998;
    wire N__48995;
    wire N__48988;
    wire N__48985;
    wire N__48982;
    wire N__48979;
    wire N__48976;
    wire N__48973;
    wire N__48970;
    wire N__48967;
    wire N__48964;
    wire N__48963;
    wire N__48962;
    wire N__48961;
    wire N__48958;
    wire N__48955;
    wire N__48952;
    wire N__48949;
    wire N__48946;
    wire N__48943;
    wire N__48940;
    wire N__48937;
    wire N__48934;
    wire N__48929;
    wire N__48926;
    wire N__48921;
    wire N__48916;
    wire N__48913;
    wire N__48910;
    wire N__48907;
    wire N__48904;
    wire N__48901;
    wire N__48898;
    wire N__48895;
    wire N__48892;
    wire N__48889;
    wire N__48886;
    wire N__48883;
    wire N__48880;
    wire N__48877;
    wire N__48874;
    wire N__48871;
    wire N__48870;
    wire N__48869;
    wire N__48866;
    wire N__48861;
    wire N__48856;
    wire N__48853;
    wire N__48850;
    wire N__48847;
    wire N__48844;
    wire N__48841;
    wire N__48838;
    wire N__48837;
    wire N__48836;
    wire N__48835;
    wire N__48830;
    wire N__48825;
    wire N__48820;
    wire N__48817;
    wire N__48814;
    wire N__48811;
    wire N__48808;
    wire N__48805;
    wire N__48804;
    wire N__48801;
    wire N__48800;
    wire N__48799;
    wire N__48796;
    wire N__48793;
    wire N__48790;
    wire N__48785;
    wire N__48780;
    wire N__48777;
    wire N__48772;
    wire N__48771;
    wire N__48770;
    wire N__48767;
    wire N__48764;
    wire N__48763;
    wire N__48760;
    wire N__48757;
    wire N__48754;
    wire N__48749;
    wire N__48744;
    wire N__48741;
    wire N__48736;
    wire N__48733;
    wire N__48730;
    wire N__48727;
    wire N__48726;
    wire N__48723;
    wire N__48720;
    wire N__48715;
    wire N__48712;
    wire N__48709;
    wire N__48708;
    wire N__48705;
    wire N__48702;
    wire N__48701;
    wire N__48696;
    wire N__48693;
    wire N__48692;
    wire N__48691;
    wire N__48686;
    wire N__48683;
    wire N__48680;
    wire N__48677;
    wire N__48674;
    wire N__48671;
    wire N__48666;
    wire N__48663;
    wire N__48660;
    wire N__48657;
    wire N__48652;
    wire N__48649;
    wire N__48646;
    wire N__48643;
    wire N__48640;
    wire N__48637;
    wire N__48634;
    wire N__48631;
    wire N__48628;
    wire N__48625;
    wire N__48624;
    wire N__48621;
    wire N__48618;
    wire N__48617;
    wire N__48614;
    wire N__48611;
    wire N__48608;
    wire N__48603;
    wire N__48598;
    wire N__48597;
    wire N__48594;
    wire N__48591;
    wire N__48588;
    wire N__48583;
    wire N__48580;
    wire N__48577;
    wire N__48574;
    wire N__48571;
    wire N__48568;
    wire N__48565;
    wire N__48562;
    wire N__48559;
    wire N__48558;
    wire N__48557;
    wire N__48556;
    wire N__48555;
    wire N__48554;
    wire N__48553;
    wire N__48552;
    wire N__48551;
    wire N__48550;
    wire N__48549;
    wire N__48548;
    wire N__48545;
    wire N__48544;
    wire N__48543;
    wire N__48540;
    wire N__48535;
    wire N__48526;
    wire N__48523;
    wire N__48518;
    wire N__48515;
    wire N__48508;
    wire N__48503;
    wire N__48490;
    wire N__48487;
    wire N__48484;
    wire N__48481;
    wire N__48478;
    wire N__48475;
    wire N__48472;
    wire N__48469;
    wire N__48466;
    wire N__48463;
    wire N__48460;
    wire N__48457;
    wire N__48454;
    wire N__48451;
    wire N__48448;
    wire N__48445;
    wire N__48442;
    wire N__48439;
    wire N__48436;
    wire N__48433;
    wire N__48430;
    wire N__48427;
    wire N__48424;
    wire N__48421;
    wire N__48418;
    wire N__48415;
    wire N__48412;
    wire N__48409;
    wire N__48406;
    wire N__48403;
    wire N__48400;
    wire N__48397;
    wire N__48396;
    wire N__48393;
    wire N__48390;
    wire N__48385;
    wire N__48384;
    wire N__48381;
    wire N__48378;
    wire N__48375;
    wire N__48372;
    wire N__48371;
    wire N__48366;
    wire N__48363;
    wire N__48358;
    wire N__48355;
    wire N__48352;
    wire N__48349;
    wire N__48346;
    wire N__48343;
    wire N__48340;
    wire N__48337;
    wire N__48334;
    wire N__48331;
    wire N__48328;
    wire N__48327;
    wire N__48326;
    wire N__48325;
    wire N__48322;
    wire N__48321;
    wire N__48318;
    wire N__48315;
    wire N__48312;
    wire N__48309;
    wire N__48304;
    wire N__48295;
    wire N__48292;
    wire N__48291;
    wire N__48288;
    wire N__48287;
    wire N__48286;
    wire N__48283;
    wire N__48280;
    wire N__48277;
    wire N__48274;
    wire N__48265;
    wire N__48262;
    wire N__48261;
    wire N__48258;
    wire N__48255;
    wire N__48254;
    wire N__48251;
    wire N__48248;
    wire N__48245;
    wire N__48242;
    wire N__48239;
    wire N__48232;
    wire N__48229;
    wire N__48226;
    wire N__48225;
    wire N__48220;
    wire N__48217;
    wire N__48216;
    wire N__48213;
    wire N__48210;
    wire N__48205;
    wire N__48202;
    wire N__48199;
    wire N__48196;
    wire N__48195;
    wire N__48194;
    wire N__48191;
    wire N__48186;
    wire N__48181;
    wire N__48178;
    wire N__48175;
    wire N__48172;
    wire N__48169;
    wire N__48166;
    wire N__48163;
    wire N__48160;
    wire N__48157;
    wire N__48154;
    wire N__48151;
    wire N__48148;
    wire N__48145;
    wire N__48142;
    wire N__48139;
    wire N__48136;
    wire N__48133;
    wire N__48130;
    wire N__48127;
    wire N__48124;
    wire N__48121;
    wire N__48118;
    wire N__48115;
    wire N__48112;
    wire N__48109;
    wire N__48108;
    wire N__48107;
    wire N__48104;
    wire N__48103;
    wire N__48100;
    wire N__48097;
    wire N__48094;
    wire N__48091;
    wire N__48088;
    wire N__48085;
    wire N__48082;
    wire N__48079;
    wire N__48074;
    wire N__48067;
    wire N__48064;
    wire N__48063;
    wire N__48062;
    wire N__48059;
    wire N__48056;
    wire N__48053;
    wire N__48050;
    wire N__48047;
    wire N__48044;
    wire N__48039;
    wire N__48036;
    wire N__48031;
    wire N__48028;
    wire N__48025;
    wire N__48022;
    wire N__48019;
    wire N__48016;
    wire N__48013;
    wire N__48010;
    wire N__48007;
    wire N__48004;
    wire N__48001;
    wire N__47998;
    wire N__47995;
    wire N__47992;
    wire N__47989;
    wire N__47986;
    wire N__47985;
    wire N__47984;
    wire N__47981;
    wire N__47980;
    wire N__47977;
    wire N__47974;
    wire N__47973;
    wire N__47970;
    wire N__47967;
    wire N__47964;
    wire N__47961;
    wire N__47958;
    wire N__47955;
    wire N__47954;
    wire N__47951;
    wire N__47948;
    wire N__47945;
    wire N__47942;
    wire N__47939;
    wire N__47936;
    wire N__47933;
    wire N__47928;
    wire N__47923;
    wire N__47914;
    wire N__47913;
    wire N__47912;
    wire N__47909;
    wire N__47908;
    wire N__47905;
    wire N__47902;
    wire N__47899;
    wire N__47894;
    wire N__47887;
    wire N__47886;
    wire N__47885;
    wire N__47882;
    wire N__47879;
    wire N__47874;
    wire N__47869;
    wire N__47866;
    wire N__47863;
    wire N__47860;
    wire N__47857;
    wire N__47854;
    wire N__47851;
    wire N__47848;
    wire N__47845;
    wire N__47842;
    wire N__47839;
    wire N__47836;
    wire N__47833;
    wire N__47830;
    wire N__47827;
    wire N__47824;
    wire N__47821;
    wire N__47818;
    wire N__47815;
    wire N__47812;
    wire N__47809;
    wire N__47806;
    wire N__47803;
    wire N__47800;
    wire N__47797;
    wire N__47794;
    wire N__47791;
    wire N__47788;
    wire N__47785;
    wire N__47782;
    wire N__47779;
    wire N__47776;
    wire N__47773;
    wire N__47770;
    wire N__47767;
    wire N__47764;
    wire N__47761;
    wire N__47758;
    wire N__47755;
    wire N__47752;
    wire N__47749;
    wire N__47746;
    wire N__47743;
    wire N__47740;
    wire N__47739;
    wire N__47734;
    wire N__47731;
    wire N__47728;
    wire N__47725;
    wire N__47722;
    wire N__47721;
    wire N__47720;
    wire N__47717;
    wire N__47714;
    wire N__47711;
    wire N__47706;
    wire N__47701;
    wire N__47698;
    wire N__47695;
    wire N__47692;
    wire N__47689;
    wire N__47686;
    wire N__47683;
    wire N__47680;
    wire N__47677;
    wire N__47674;
    wire N__47671;
    wire N__47668;
    wire N__47665;
    wire N__47662;
    wire N__47659;
    wire N__47656;
    wire N__47653;
    wire N__47650;
    wire N__47647;
    wire N__47644;
    wire N__47641;
    wire N__47638;
    wire N__47635;
    wire N__47632;
    wire N__47629;
    wire N__47626;
    wire N__47623;
    wire N__47620;
    wire N__47617;
    wire N__47614;
    wire N__47611;
    wire N__47608;
    wire N__47605;
    wire N__47602;
    wire N__47599;
    wire N__47596;
    wire N__47593;
    wire N__47590;
    wire N__47587;
    wire N__47584;
    wire N__47581;
    wire N__47578;
    wire N__47575;
    wire N__47572;
    wire N__47569;
    wire N__47566;
    wire N__47563;
    wire N__47560;
    wire N__47557;
    wire N__47554;
    wire N__47553;
    wire N__47550;
    wire N__47549;
    wire N__47546;
    wire N__47543;
    wire N__47540;
    wire N__47537;
    wire N__47534;
    wire N__47529;
    wire N__47526;
    wire N__47521;
    wire N__47520;
    wire N__47517;
    wire N__47516;
    wire N__47513;
    wire N__47512;
    wire N__47509;
    wire N__47508;
    wire N__47505;
    wire N__47502;
    wire N__47499;
    wire N__47496;
    wire N__47493;
    wire N__47490;
    wire N__47487;
    wire N__47484;
    wire N__47483;
    wire N__47482;
    wire N__47481;
    wire N__47480;
    wire N__47475;
    wire N__47468;
    wire N__47459;
    wire N__47452;
    wire N__47451;
    wire N__47448;
    wire N__47447;
    wire N__47446;
    wire N__47445;
    wire N__47442;
    wire N__47439;
    wire N__47438;
    wire N__47437;
    wire N__47436;
    wire N__47435;
    wire N__47434;
    wire N__47433;
    wire N__47432;
    wire N__47431;
    wire N__47424;
    wire N__47421;
    wire N__47418;
    wire N__47415;
    wire N__47412;
    wire N__47411;
    wire N__47410;
    wire N__47409;
    wire N__47404;
    wire N__47399;
    wire N__47398;
    wire N__47397;
    wire N__47394;
    wire N__47391;
    wire N__47388;
    wire N__47379;
    wire N__47372;
    wire N__47369;
    wire N__47366;
    wire N__47361;
    wire N__47358;
    wire N__47357;
    wire N__47356;
    wire N__47355;
    wire N__47354;
    wire N__47351;
    wire N__47344;
    wire N__47343;
    wire N__47342;
    wire N__47339;
    wire N__47332;
    wire N__47327;
    wire N__47324;
    wire N__47321;
    wire N__47316;
    wire N__47311;
    wire N__47296;
    wire N__47293;
    wire N__47290;
    wire N__47287;
    wire N__47284;
    wire N__47281;
    wire N__47278;
    wire N__47275;
    wire N__47272;
    wire N__47269;
    wire N__47266;
    wire N__47263;
    wire N__47260;
    wire N__47257;
    wire N__47254;
    wire N__47251;
    wire N__47248;
    wire N__47245;
    wire N__47242;
    wire N__47239;
    wire N__47236;
    wire N__47233;
    wire N__47230;
    wire N__47229;
    wire N__47228;
    wire N__47225;
    wire N__47220;
    wire N__47217;
    wire N__47212;
    wire N__47209;
    wire N__47206;
    wire N__47203;
    wire N__47200;
    wire N__47197;
    wire N__47194;
    wire N__47193;
    wire N__47190;
    wire N__47187;
    wire N__47186;
    wire N__47183;
    wire N__47180;
    wire N__47177;
    wire N__47174;
    wire N__47171;
    wire N__47168;
    wire N__47165;
    wire N__47160;
    wire N__47157;
    wire N__47154;
    wire N__47149;
    wire N__47146;
    wire N__47143;
    wire N__47142;
    wire N__47139;
    wire N__47136;
    wire N__47135;
    wire N__47130;
    wire N__47129;
    wire N__47126;
    wire N__47123;
    wire N__47120;
    wire N__47117;
    wire N__47112;
    wire N__47109;
    wire N__47106;
    wire N__47101;
    wire N__47098;
    wire N__47095;
    wire N__47092;
    wire N__47089;
    wire N__47086;
    wire N__47085;
    wire N__47084;
    wire N__47081;
    wire N__47078;
    wire N__47075;
    wire N__47072;
    wire N__47069;
    wire N__47062;
    wire N__47059;
    wire N__47056;
    wire N__47053;
    wire N__47050;
    wire N__47047;
    wire N__47046;
    wire N__47043;
    wire N__47040;
    wire N__47037;
    wire N__47034;
    wire N__47029;
    wire N__47026;
    wire N__47025;
    wire N__47022;
    wire N__47019;
    wire N__47016;
    wire N__47011;
    wire N__47008;
    wire N__47005;
    wire N__47002;
    wire N__46999;
    wire N__46996;
    wire N__46995;
    wire N__46994;
    wire N__46991;
    wire N__46988;
    wire N__46985;
    wire N__46982;
    wire N__46979;
    wire N__46976;
    wire N__46971;
    wire N__46966;
    wire N__46963;
    wire N__46962;
    wire N__46959;
    wire N__46956;
    wire N__46955;
    wire N__46952;
    wire N__46949;
    wire N__46946;
    wire N__46943;
    wire N__46940;
    wire N__46933;
    wire N__46930;
    wire N__46927;
    wire N__46924;
    wire N__46921;
    wire N__46918;
    wire N__46915;
    wire N__46912;
    wire N__46909;
    wire N__46908;
    wire N__46907;
    wire N__46904;
    wire N__46901;
    wire N__46898;
    wire N__46895;
    wire N__46894;
    wire N__46889;
    wire N__46886;
    wire N__46883;
    wire N__46880;
    wire N__46877;
    wire N__46874;
    wire N__46871;
    wire N__46864;
    wire N__46861;
    wire N__46858;
    wire N__46855;
    wire N__46852;
    wire N__46849;
    wire N__46846;
    wire N__46843;
    wire N__46840;
    wire N__46837;
    wire N__46834;
    wire N__46831;
    wire N__46828;
    wire N__46825;
    wire N__46822;
    wire N__46819;
    wire N__46816;
    wire N__46813;
    wire N__46810;
    wire N__46807;
    wire N__46804;
    wire N__46803;
    wire N__46800;
    wire N__46797;
    wire N__46796;
    wire N__46793;
    wire N__46792;
    wire N__46789;
    wire N__46786;
    wire N__46783;
    wire N__46780;
    wire N__46777;
    wire N__46772;
    wire N__46769;
    wire N__46766;
    wire N__46759;
    wire N__46756;
    wire N__46753;
    wire N__46750;
    wire N__46747;
    wire N__46744;
    wire N__46741;
    wire N__46740;
    wire N__46739;
    wire N__46736;
    wire N__46733;
    wire N__46730;
    wire N__46727;
    wire N__46724;
    wire N__46721;
    wire N__46718;
    wire N__46715;
    wire N__46710;
    wire N__46705;
    wire N__46704;
    wire N__46701;
    wire N__46700;
    wire N__46697;
    wire N__46694;
    wire N__46691;
    wire N__46688;
    wire N__46685;
    wire N__46678;
    wire N__46675;
    wire N__46672;
    wire N__46669;
    wire N__46666;
    wire N__46663;
    wire N__46660;
    wire N__46657;
    wire N__46654;
    wire N__46651;
    wire N__46648;
    wire N__46645;
    wire N__46644;
    wire N__46643;
    wire N__46642;
    wire N__46639;
    wire N__46634;
    wire N__46629;
    wire N__46626;
    wire N__46623;
    wire N__46620;
    wire N__46617;
    wire N__46612;
    wire N__46609;
    wire N__46606;
    wire N__46603;
    wire N__46600;
    wire N__46597;
    wire N__46594;
    wire N__46591;
    wire N__46588;
    wire N__46585;
    wire N__46582;
    wire N__46579;
    wire N__46576;
    wire N__46573;
    wire N__46570;
    wire N__46567;
    wire N__46564;
    wire N__46561;
    wire N__46558;
    wire N__46555;
    wire N__46552;
    wire N__46549;
    wire N__46546;
    wire N__46543;
    wire N__46540;
    wire N__46537;
    wire N__46534;
    wire N__46531;
    wire N__46528;
    wire N__46527;
    wire N__46524;
    wire N__46521;
    wire N__46520;
    wire N__46517;
    wire N__46514;
    wire N__46513;
    wire N__46510;
    wire N__46507;
    wire N__46504;
    wire N__46499;
    wire N__46496;
    wire N__46493;
    wire N__46490;
    wire N__46483;
    wire N__46480;
    wire N__46479;
    wire N__46476;
    wire N__46473;
    wire N__46472;
    wire N__46469;
    wire N__46466;
    wire N__46463;
    wire N__46458;
    wire N__46453;
    wire N__46450;
    wire N__46447;
    wire N__46444;
    wire N__46443;
    wire N__46442;
    wire N__46441;
    wire N__46440;
    wire N__46439;
    wire N__46432;
    wire N__46427;
    wire N__46424;
    wire N__46417;
    wire N__46414;
    wire N__46411;
    wire N__46408;
    wire N__46405;
    wire N__46402;
    wire N__46399;
    wire N__46396;
    wire N__46393;
    wire N__46390;
    wire N__46387;
    wire N__46384;
    wire N__46381;
    wire N__46378;
    wire N__46375;
    wire N__46372;
    wire N__46369;
    wire N__46366;
    wire N__46365;
    wire N__46362;
    wire N__46359;
    wire N__46356;
    wire N__46353;
    wire N__46348;
    wire N__46345;
    wire N__46342;
    wire N__46339;
    wire N__46338;
    wire N__46335;
    wire N__46334;
    wire N__46331;
    wire N__46330;
    wire N__46329;
    wire N__46326;
    wire N__46321;
    wire N__46316;
    wire N__46313;
    wire N__46306;
    wire N__46305;
    wire N__46304;
    wire N__46303;
    wire N__46294;
    wire N__46291;
    wire N__46288;
    wire N__46287;
    wire N__46286;
    wire N__46283;
    wire N__46280;
    wire N__46275;
    wire N__46270;
    wire N__46269;
    wire N__46268;
    wire N__46267;
    wire N__46266;
    wire N__46265;
    wire N__46256;
    wire N__46251;
    wire N__46246;
    wire N__46243;
    wire N__46242;
    wire N__46239;
    wire N__46236;
    wire N__46231;
    wire N__46228;
    wire N__46225;
    wire N__46224;
    wire N__46221;
    wire N__46218;
    wire N__46215;
    wire N__46210;
    wire N__46207;
    wire N__46206;
    wire N__46203;
    wire N__46200;
    wire N__46195;
    wire N__46192;
    wire N__46191;
    wire N__46188;
    wire N__46185;
    wire N__46182;
    wire N__46179;
    wire N__46174;
    wire N__46171;
    wire N__46168;
    wire N__46165;
    wire N__46162;
    wire N__46159;
    wire N__46156;
    wire N__46153;
    wire N__46150;
    wire N__46147;
    wire N__46144;
    wire N__46141;
    wire N__46138;
    wire N__46135;
    wire N__46132;
    wire N__46129;
    wire N__46126;
    wire N__46123;
    wire N__46120;
    wire N__46117;
    wire N__46114;
    wire N__46113;
    wire N__46110;
    wire N__46107;
    wire N__46104;
    wire N__46101;
    wire N__46096;
    wire N__46093;
    wire N__46090;
    wire N__46087;
    wire N__46084;
    wire N__46081;
    wire N__46078;
    wire N__46077;
    wire N__46076;
    wire N__46075;
    wire N__46074;
    wire N__46073;
    wire N__46070;
    wire N__46069;
    wire N__46066;
    wire N__46057;
    wire N__46052;
    wire N__46045;
    wire N__46042;
    wire N__46039;
    wire N__46036;
    wire N__46033;
    wire N__46032;
    wire N__46029;
    wire N__46026;
    wire N__46021;
    wire N__46018;
    wire N__46017;
    wire N__46014;
    wire N__46011;
    wire N__46008;
    wire N__46003;
    wire N__46000;
    wire N__45999;
    wire N__45996;
    wire N__45993;
    wire N__45988;
    wire N__45985;
    wire N__45984;
    wire N__45981;
    wire N__45980;
    wire N__45979;
    wire N__45976;
    wire N__45973;
    wire N__45968;
    wire N__45961;
    wire N__45960;
    wire N__45957;
    wire N__45954;
    wire N__45949;
    wire N__45946;
    wire N__45945;
    wire N__45942;
    wire N__45939;
    wire N__45934;
    wire N__45933;
    wire N__45930;
    wire N__45927;
    wire N__45924;
    wire N__45919;
    wire N__45918;
    wire N__45915;
    wire N__45914;
    wire N__45913;
    wire N__45912;
    wire N__45909;
    wire N__45908;
    wire N__45907;
    wire N__45898;
    wire N__45891;
    wire N__45886;
    wire N__45883;
    wire N__45880;
    wire N__45877;
    wire N__45874;
    wire N__45871;
    wire N__45870;
    wire N__45867;
    wire N__45864;
    wire N__45861;
    wire N__45856;
    wire N__45855;
    wire N__45852;
    wire N__45849;
    wire N__45844;
    wire N__45843;
    wire N__45842;
    wire N__45841;
    wire N__45840;
    wire N__45837;
    wire N__45834;
    wire N__45831;
    wire N__45826;
    wire N__45821;
    wire N__45816;
    wire N__45811;
    wire N__45808;
    wire N__45805;
    wire N__45802;
    wire N__45799;
    wire N__45796;
    wire N__45795;
    wire N__45794;
    wire N__45791;
    wire N__45790;
    wire N__45789;
    wire N__45786;
    wire N__45785;
    wire N__45782;
    wire N__45781;
    wire N__45780;
    wire N__45777;
    wire N__45772;
    wire N__45769;
    wire N__45766;
    wire N__45759;
    wire N__45748;
    wire N__45745;
    wire N__45742;
    wire N__45739;
    wire N__45736;
    wire N__45733;
    wire N__45730;
    wire N__45727;
    wire N__45724;
    wire N__45721;
    wire N__45718;
    wire N__45715;
    wire N__45714;
    wire N__45711;
    wire N__45708;
    wire N__45703;
    wire N__45700;
    wire N__45697;
    wire N__45696;
    wire N__45693;
    wire N__45690;
    wire N__45685;
    wire N__45682;
    wire N__45681;
    wire N__45678;
    wire N__45675;
    wire N__45672;
    wire N__45669;
    wire N__45666;
    wire N__45663;
    wire N__45660;
    wire N__45657;
    wire N__45654;
    wire N__45651;
    wire N__45646;
    wire N__45645;
    wire N__45642;
    wire N__45639;
    wire N__45636;
    wire N__45633;
    wire N__45630;
    wire N__45627;
    wire N__45624;
    wire N__45621;
    wire N__45618;
    wire N__45613;
    wire N__45610;
    wire N__45607;
    wire N__45606;
    wire N__45603;
    wire N__45600;
    wire N__45597;
    wire N__45594;
    wire N__45591;
    wire N__45588;
    wire N__45585;
    wire N__45582;
    wire N__45577;
    wire N__45574;
    wire N__45571;
    wire N__45570;
    wire N__45567;
    wire N__45564;
    wire N__45561;
    wire N__45558;
    wire N__45555;
    wire N__45552;
    wire N__45549;
    wire N__45546;
    wire N__45541;
    wire N__45538;
    wire N__45537;
    wire N__45536;
    wire N__45533;
    wire N__45530;
    wire N__45527;
    wire N__45520;
    wire N__45517;
    wire N__45516;
    wire N__45513;
    wire N__45510;
    wire N__45507;
    wire N__45504;
    wire N__45499;
    wire N__45496;
    wire N__45495;
    wire N__45492;
    wire N__45489;
    wire N__45484;
    wire N__45481;
    wire N__45478;
    wire N__45475;
    wire N__45472;
    wire N__45469;
    wire N__45466;
    wire N__45463;
    wire N__45460;
    wire N__45457;
    wire N__45454;
    wire N__45451;
    wire N__45448;
    wire N__45445;
    wire N__45442;
    wire N__45439;
    wire N__45436;
    wire N__45433;
    wire N__45430;
    wire N__45427;
    wire N__45424;
    wire N__45421;
    wire N__45418;
    wire N__45415;
    wire N__45412;
    wire N__45409;
    wire N__45406;
    wire N__45403;
    wire N__45400;
    wire N__45397;
    wire N__45394;
    wire N__45391;
    wire N__45388;
    wire N__45385;
    wire N__45382;
    wire N__45379;
    wire N__45376;
    wire N__45375;
    wire N__45372;
    wire N__45369;
    wire N__45366;
    wire N__45363;
    wire N__45360;
    wire N__45357;
    wire N__45354;
    wire N__45351;
    wire N__45348;
    wire N__45345;
    wire N__45340;
    wire N__45339;
    wire N__45336;
    wire N__45333;
    wire N__45330;
    wire N__45327;
    wire N__45324;
    wire N__45321;
    wire N__45318;
    wire N__45315;
    wire N__45312;
    wire N__45307;
    wire N__45304;
    wire N__45301;
    wire N__45298;
    wire N__45297;
    wire N__45294;
    wire N__45291;
    wire N__45288;
    wire N__45285;
    wire N__45282;
    wire N__45279;
    wire N__45274;
    wire N__45271;
    wire N__45268;
    wire N__45267;
    wire N__45266;
    wire N__45263;
    wire N__45260;
    wire N__45259;
    wire N__45256;
    wire N__45253;
    wire N__45248;
    wire N__45241;
    wire N__45238;
    wire N__45237;
    wire N__45236;
    wire N__45235;
    wire N__45232;
    wire N__45229;
    wire N__45226;
    wire N__45223;
    wire N__45214;
    wire N__45211;
    wire N__45208;
    wire N__45205;
    wire N__45202;
    wire N__45199;
    wire N__45196;
    wire N__45193;
    wire N__45190;
    wire N__45187;
    wire N__45184;
    wire N__45183;
    wire N__45182;
    wire N__45181;
    wire N__45178;
    wire N__45175;
    wire N__45172;
    wire N__45169;
    wire N__45166;
    wire N__45163;
    wire N__45156;
    wire N__45151;
    wire N__45148;
    wire N__45145;
    wire N__45142;
    wire N__45139;
    wire N__45136;
    wire N__45133;
    wire N__45132;
    wire N__45129;
    wire N__45128;
    wire N__45125;
    wire N__45122;
    wire N__45119;
    wire N__45116;
    wire N__45111;
    wire N__45106;
    wire N__45103;
    wire N__45102;
    wire N__45099;
    wire N__45096;
    wire N__45093;
    wire N__45092;
    wire N__45089;
    wire N__45086;
    wire N__45083;
    wire N__45076;
    wire N__45073;
    wire N__45070;
    wire N__45067;
    wire N__45064;
    wire N__45061;
    wire N__45060;
    wire N__45059;
    wire N__45056;
    wire N__45053;
    wire N__45050;
    wire N__45047;
    wire N__45044;
    wire N__45041;
    wire N__45038;
    wire N__45035;
    wire N__45028;
    wire N__45025;
    wire N__45022;
    wire N__45021;
    wire N__45018;
    wire N__45017;
    wire N__45014;
    wire N__45011;
    wire N__45008;
    wire N__45001;
    wire N__44998;
    wire N__44995;
    wire N__44992;
    wire N__44989;
    wire N__44986;
    wire N__44983;
    wire N__44982;
    wire N__44979;
    wire N__44978;
    wire N__44975;
    wire N__44972;
    wire N__44969;
    wire N__44966;
    wire N__44963;
    wire N__44956;
    wire N__44955;
    wire N__44952;
    wire N__44949;
    wire N__44946;
    wire N__44941;
    wire N__44938;
    wire N__44937;
    wire N__44934;
    wire N__44931;
    wire N__44928;
    wire N__44923;
    wire N__44922;
    wire N__44921;
    wire N__44916;
    wire N__44913;
    wire N__44908;
    wire N__44907;
    wire N__44906;
    wire N__44905;
    wire N__44902;
    wire N__44899;
    wire N__44898;
    wire N__44897;
    wire N__44892;
    wire N__44891;
    wire N__44886;
    wire N__44881;
    wire N__44878;
    wire N__44875;
    wire N__44866;
    wire N__44865;
    wire N__44862;
    wire N__44859;
    wire N__44856;
    wire N__44853;
    wire N__44852;
    wire N__44851;
    wire N__44848;
    wire N__44845;
    wire N__44842;
    wire N__44839;
    wire N__44836;
    wire N__44833;
    wire N__44830;
    wire N__44827;
    wire N__44818;
    wire N__44815;
    wire N__44814;
    wire N__44811;
    wire N__44808;
    wire N__44805;
    wire N__44804;
    wire N__44801;
    wire N__44798;
    wire N__44795;
    wire N__44788;
    wire N__44785;
    wire N__44782;
    wire N__44779;
    wire N__44778;
    wire N__44775;
    wire N__44774;
    wire N__44771;
    wire N__44768;
    wire N__44765;
    wire N__44758;
    wire N__44755;
    wire N__44754;
    wire N__44753;
    wire N__44750;
    wire N__44747;
    wire N__44744;
    wire N__44741;
    wire N__44734;
    wire N__44731;
    wire N__44728;
    wire N__44725;
    wire N__44722;
    wire N__44719;
    wire N__44716;
    wire N__44713;
    wire N__44710;
    wire N__44709;
    wire N__44708;
    wire N__44705;
    wire N__44700;
    wire N__44697;
    wire N__44692;
    wire N__44689;
    wire N__44686;
    wire N__44683;
    wire N__44682;
    wire N__44681;
    wire N__44680;
    wire N__44679;
    wire N__44678;
    wire N__44675;
    wire N__44672;
    wire N__44669;
    wire N__44668;
    wire N__44665;
    wire N__44662;
    wire N__44659;
    wire N__44656;
    wire N__44651;
    wire N__44650;
    wire N__44649;
    wire N__44648;
    wire N__44645;
    wire N__44638;
    wire N__44635;
    wire N__44632;
    wire N__44627;
    wire N__44622;
    wire N__44619;
    wire N__44608;
    wire N__44607;
    wire N__44604;
    wire N__44601;
    wire N__44598;
    wire N__44597;
    wire N__44596;
    wire N__44595;
    wire N__44594;
    wire N__44593;
    wire N__44590;
    wire N__44587;
    wire N__44584;
    wire N__44581;
    wire N__44578;
    wire N__44575;
    wire N__44574;
    wire N__44573;
    wire N__44572;
    wire N__44571;
    wire N__44570;
    wire N__44567;
    wire N__44564;
    wire N__44559;
    wire N__44552;
    wire N__44547;
    wire N__44544;
    wire N__44539;
    wire N__44536;
    wire N__44521;
    wire N__44518;
    wire N__44515;
    wire N__44514;
    wire N__44513;
    wire N__44512;
    wire N__44511;
    wire N__44510;
    wire N__44509;
    wire N__44506;
    wire N__44503;
    wire N__44502;
    wire N__44499;
    wire N__44496;
    wire N__44493;
    wire N__44490;
    wire N__44487;
    wire N__44482;
    wire N__44479;
    wire N__44478;
    wire N__44475;
    wire N__44468;
    wire N__44467;
    wire N__44466;
    wire N__44459;
    wire N__44458;
    wire N__44457;
    wire N__44456;
    wire N__44453;
    wire N__44448;
    wire N__44445;
    wire N__44442;
    wire N__44439;
    wire N__44434;
    wire N__44431;
    wire N__44422;
    wire N__44413;
    wire N__44410;
    wire N__44407;
    wire N__44404;
    wire N__44401;
    wire N__44398;
    wire N__44395;
    wire N__44392;
    wire N__44389;
    wire N__44386;
    wire N__44383;
    wire N__44382;
    wire N__44379;
    wire N__44376;
    wire N__44371;
    wire N__44368;
    wire N__44365;
    wire N__44362;
    wire N__44359;
    wire N__44356;
    wire N__44353;
    wire N__44350;
    wire N__44347;
    wire N__44344;
    wire N__44343;
    wire N__44340;
    wire N__44337;
    wire N__44334;
    wire N__44331;
    wire N__44330;
    wire N__44329;
    wire N__44328;
    wire N__44325;
    wire N__44322;
    wire N__44319;
    wire N__44314;
    wire N__44305;
    wire N__44304;
    wire N__44301;
    wire N__44298;
    wire N__44293;
    wire N__44292;
    wire N__44289;
    wire N__44286;
    wire N__44281;
    wire N__44280;
    wire N__44279;
    wire N__44278;
    wire N__44275;
    wire N__44272;
    wire N__44269;
    wire N__44266;
    wire N__44263;
    wire N__44260;
    wire N__44257;
    wire N__44256;
    wire N__44251;
    wire N__44246;
    wire N__44243;
    wire N__44240;
    wire N__44233;
    wire N__44230;
    wire N__44227;
    wire N__44224;
    wire N__44221;
    wire N__44220;
    wire N__44217;
    wire N__44214;
    wire N__44209;
    wire N__44206;
    wire N__44203;
    wire N__44200;
    wire N__44197;
    wire N__44194;
    wire N__44191;
    wire N__44188;
    wire N__44185;
    wire N__44182;
    wire N__44179;
    wire N__44176;
    wire N__44173;
    wire N__44170;
    wire N__44167;
    wire N__44164;
    wire N__44163;
    wire N__44160;
    wire N__44157;
    wire N__44154;
    wire N__44149;
    wire N__44146;
    wire N__44143;
    wire N__44142;
    wire N__44139;
    wire N__44136;
    wire N__44131;
    wire N__44128;
    wire N__44125;
    wire N__44122;
    wire N__44119;
    wire N__44118;
    wire N__44115;
    wire N__44114;
    wire N__44113;
    wire N__44110;
    wire N__44107;
    wire N__44104;
    wire N__44101;
    wire N__44092;
    wire N__44089;
    wire N__44086;
    wire N__44083;
    wire N__44080;
    wire N__44077;
    wire N__44074;
    wire N__44071;
    wire N__44068;
    wire N__44065;
    wire N__44062;
    wire N__44059;
    wire N__44056;
    wire N__44053;
    wire N__44050;
    wire N__44047;
    wire N__44044;
    wire N__44041;
    wire N__44038;
    wire N__44035;
    wire N__44032;
    wire N__44029;
    wire N__44026;
    wire N__44023;
    wire N__44020;
    wire N__44017;
    wire N__44014;
    wire N__44011;
    wire N__44008;
    wire N__44005;
    wire N__44002;
    wire N__43999;
    wire N__43996;
    wire N__43993;
    wire N__43990;
    wire N__43987;
    wire N__43986;
    wire N__43983;
    wire N__43980;
    wire N__43975;
    wire N__43972;
    wire N__43969;
    wire N__43966;
    wire N__43963;
    wire N__43960;
    wire N__43957;
    wire N__43954;
    wire N__43951;
    wire N__43948;
    wire N__43945;
    wire N__43944;
    wire N__43941;
    wire N__43938;
    wire N__43933;
    wire N__43930;
    wire N__43927;
    wire N__43924;
    wire N__43923;
    wire N__43920;
    wire N__43917;
    wire N__43916;
    wire N__43913;
    wire N__43910;
    wire N__43907;
    wire N__43900;
    wire N__43897;
    wire N__43894;
    wire N__43891;
    wire N__43888;
    wire N__43885;
    wire N__43882;
    wire N__43879;
    wire N__43876;
    wire N__43873;
    wire N__43870;
    wire N__43867;
    wire N__43864;
    wire N__43861;
    wire N__43858;
    wire N__43855;
    wire N__43852;
    wire N__43849;
    wire N__43846;
    wire N__43845;
    wire N__43842;
    wire N__43839;
    wire N__43836;
    wire N__43833;
    wire N__43828;
    wire N__43825;
    wire N__43822;
    wire N__43819;
    wire N__43816;
    wire N__43813;
    wire N__43810;
    wire N__43807;
    wire N__43804;
    wire N__43803;
    wire N__43800;
    wire N__43797;
    wire N__43792;
    wire N__43789;
    wire N__43786;
    wire N__43783;
    wire N__43780;
    wire N__43779;
    wire N__43774;
    wire N__43771;
    wire N__43768;
    wire N__43765;
    wire N__43764;
    wire N__43761;
    wire N__43758;
    wire N__43755;
    wire N__43752;
    wire N__43747;
    wire N__43746;
    wire N__43741;
    wire N__43738;
    wire N__43737;
    wire N__43736;
    wire N__43731;
    wire N__43728;
    wire N__43727;
    wire N__43726;
    wire N__43723;
    wire N__43718;
    wire N__43717;
    wire N__43714;
    wire N__43713;
    wire N__43712;
    wire N__43711;
    wire N__43708;
    wire N__43705;
    wire N__43702;
    wire N__43701;
    wire N__43698;
    wire N__43691;
    wire N__43686;
    wire N__43681;
    wire N__43672;
    wire N__43669;
    wire N__43666;
    wire N__43663;
    wire N__43660;
    wire N__43657;
    wire N__43654;
    wire N__43651;
    wire N__43648;
    wire N__43645;
    wire N__43642;
    wire N__43639;
    wire N__43636;
    wire N__43633;
    wire N__43630;
    wire N__43627;
    wire N__43626;
    wire N__43623;
    wire N__43620;
    wire N__43617;
    wire N__43614;
    wire N__43609;
    wire N__43606;
    wire N__43603;
    wire N__43600;
    wire N__43597;
    wire N__43594;
    wire N__43591;
    wire N__43588;
    wire N__43585;
    wire N__43584;
    wire N__43581;
    wire N__43578;
    wire N__43575;
    wire N__43570;
    wire N__43569;
    wire N__43566;
    wire N__43563;
    wire N__43562;
    wire N__43559;
    wire N__43556;
    wire N__43553;
    wire N__43546;
    wire N__43543;
    wire N__43540;
    wire N__43537;
    wire N__43534;
    wire N__43531;
    wire N__43528;
    wire N__43525;
    wire N__43524;
    wire N__43521;
    wire N__43518;
    wire N__43515;
    wire N__43512;
    wire N__43507;
    wire N__43504;
    wire N__43501;
    wire N__43498;
    wire N__43495;
    wire N__43494;
    wire N__43493;
    wire N__43490;
    wire N__43485;
    wire N__43480;
    wire N__43479;
    wire N__43476;
    wire N__43475;
    wire N__43474;
    wire N__43471;
    wire N__43468;
    wire N__43463;
    wire N__43456;
    wire N__43453;
    wire N__43450;
    wire N__43449;
    wire N__43448;
    wire N__43445;
    wire N__43442;
    wire N__43437;
    wire N__43432;
    wire N__43429;
    wire N__43428;
    wire N__43427;
    wire N__43424;
    wire N__43419;
    wire N__43414;
    wire N__43411;
    wire N__43410;
    wire N__43409;
    wire N__43406;
    wire N__43403;
    wire N__43400;
    wire N__43393;
    wire N__43390;
    wire N__43387;
    wire N__43384;
    wire N__43381;
    wire N__43378;
    wire N__43375;
    wire N__43372;
    wire N__43371;
    wire N__43368;
    wire N__43365;
    wire N__43362;
    wire N__43359;
    wire N__43356;
    wire N__43353;
    wire N__43348;
    wire N__43347;
    wire N__43344;
    wire N__43341;
    wire N__43338;
    wire N__43333;
    wire N__43332;
    wire N__43329;
    wire N__43326;
    wire N__43323;
    wire N__43318;
    wire N__43317;
    wire N__43314;
    wire N__43311;
    wire N__43308;
    wire N__43303;
    wire N__43300;
    wire N__43299;
    wire N__43296;
    wire N__43293;
    wire N__43290;
    wire N__43285;
    wire N__43282;
    wire N__43279;
    wire N__43276;
    wire N__43275;
    wire N__43272;
    wire N__43269;
    wire N__43264;
    wire N__43263;
    wire N__43260;
    wire N__43257;
    wire N__43254;
    wire N__43249;
    wire N__43248;
    wire N__43245;
    wire N__43242;
    wire N__43239;
    wire N__43234;
    wire N__43233;
    wire N__43230;
    wire N__43227;
    wire N__43224;
    wire N__43219;
    wire N__43216;
    wire N__43213;
    wire N__43212;
    wire N__43211;
    wire N__43208;
    wire N__43203;
    wire N__43198;
    wire N__43195;
    wire N__43192;
    wire N__43189;
    wire N__43186;
    wire N__43183;
    wire N__43180;
    wire N__43177;
    wire N__43174;
    wire N__43171;
    wire N__43168;
    wire N__43165;
    wire N__43162;
    wire N__43159;
    wire N__43158;
    wire N__43157;
    wire N__43154;
    wire N__43149;
    wire N__43146;
    wire N__43141;
    wire N__43138;
    wire N__43135;
    wire N__43132;
    wire N__43129;
    wire N__43126;
    wire N__43123;
    wire N__43120;
    wire N__43117;
    wire N__43114;
    wire N__43111;
    wire N__43110;
    wire N__43105;
    wire N__43102;
    wire N__43101;
    wire N__43100;
    wire N__43099;
    wire N__43092;
    wire N__43089;
    wire N__43084;
    wire N__43083;
    wire N__43082;
    wire N__43081;
    wire N__43080;
    wire N__43079;
    wire N__43078;
    wire N__43077;
    wire N__43076;
    wire N__43075;
    wire N__43074;
    wire N__43063;
    wire N__43050;
    wire N__43045;
    wire N__43044;
    wire N__43043;
    wire N__43042;
    wire N__43041;
    wire N__43038;
    wire N__43035;
    wire N__43034;
    wire N__43033;
    wire N__43030;
    wire N__43029;
    wire N__43026;
    wire N__43025;
    wire N__43024;
    wire N__43015;
    wire N__43002;
    wire N__42997;
    wire N__42996;
    wire N__42995;
    wire N__42994;
    wire N__42993;
    wire N__42992;
    wire N__42991;
    wire N__42990;
    wire N__42989;
    wire N__42986;
    wire N__42981;
    wire N__42968;
    wire N__42961;
    wire N__42958;
    wire N__42955;
    wire N__42952;
    wire N__42949;
    wire N__42946;
    wire N__42943;
    wire N__42940;
    wire N__42937;
    wire N__42934;
    wire N__42931;
    wire N__42930;
    wire N__42929;
    wire N__42926;
    wire N__42923;
    wire N__42920;
    wire N__42913;
    wire N__42910;
    wire N__42909;
    wire N__42908;
    wire N__42905;
    wire N__42902;
    wire N__42899;
    wire N__42896;
    wire N__42893;
    wire N__42886;
    wire N__42883;
    wire N__42882;
    wire N__42881;
    wire N__42878;
    wire N__42873;
    wire N__42868;
    wire N__42865;
    wire N__42864;
    wire N__42861;
    wire N__42860;
    wire N__42857;
    wire N__42852;
    wire N__42847;
    wire N__42844;
    wire N__42843;
    wire N__42842;
    wire N__42839;
    wire N__42836;
    wire N__42833;
    wire N__42826;
    wire N__42823;
    wire N__42822;
    wire N__42821;
    wire N__42820;
    wire N__42817;
    wire N__42812;
    wire N__42809;
    wire N__42802;
    wire N__42799;
    wire N__42798;
    wire N__42795;
    wire N__42794;
    wire N__42793;
    wire N__42790;
    wire N__42785;
    wire N__42782;
    wire N__42775;
    wire N__42772;
    wire N__42771;
    wire N__42770;
    wire N__42767;
    wire N__42764;
    wire N__42761;
    wire N__42754;
    wire N__42751;
    wire N__42748;
    wire N__42745;
    wire N__42742;
    wire N__42739;
    wire N__42736;
    wire N__42735;
    wire N__42732;
    wire N__42729;
    wire N__42726;
    wire N__42723;
    wire N__42718;
    wire N__42715;
    wire N__42712;
    wire N__42709;
    wire N__42708;
    wire N__42705;
    wire N__42702;
    wire N__42699;
    wire N__42696;
    wire N__42691;
    wire N__42688;
    wire N__42685;
    wire N__42682;
    wire N__42679;
    wire N__42676;
    wire N__42673;
    wire N__42670;
    wire N__42667;
    wire N__42664;
    wire N__42661;
    wire N__42658;
    wire N__42657;
    wire N__42656;
    wire N__42653;
    wire N__42650;
    wire N__42647;
    wire N__42640;
    wire N__42637;
    wire N__42636;
    wire N__42635;
    wire N__42632;
    wire N__42629;
    wire N__42626;
    wire N__42619;
    wire N__42616;
    wire N__42613;
    wire N__42610;
    wire N__42607;
    wire N__42604;
    wire N__42601;
    wire N__42600;
    wire N__42595;
    wire N__42592;
    wire N__42589;
    wire N__42586;
    wire N__42583;
    wire N__42580;
    wire N__42579;
    wire N__42574;
    wire N__42571;
    wire N__42568;
    wire N__42565;
    wire N__42562;
    wire N__42559;
    wire N__42558;
    wire N__42553;
    wire N__42550;
    wire N__42547;
    wire N__42544;
    wire N__42541;
    wire N__42538;
    wire N__42537;
    wire N__42532;
    wire N__42529;
    wire N__42526;
    wire N__42523;
    wire N__42520;
    wire N__42517;
    wire N__42516;
    wire N__42511;
    wire N__42508;
    wire N__42505;
    wire N__42502;
    wire N__42501;
    wire N__42496;
    wire N__42493;
    wire N__42490;
    wire N__42489;
    wire N__42486;
    wire N__42483;
    wire N__42478;
    wire N__42475;
    wire N__42474;
    wire N__42471;
    wire N__42468;
    wire N__42463;
    wire N__42460;
    wire N__42457;
    wire N__42454;
    wire N__42453;
    wire N__42452;
    wire N__42449;
    wire N__42444;
    wire N__42441;
    wire N__42438;
    wire N__42433;
    wire N__42430;
    wire N__42429;
    wire N__42426;
    wire N__42423;
    wire N__42420;
    wire N__42419;
    wire N__42416;
    wire N__42413;
    wire N__42410;
    wire N__42403;
    wire N__42400;
    wire N__42397;
    wire N__42396;
    wire N__42393;
    wire N__42390;
    wire N__42387;
    wire N__42384;
    wire N__42379;
    wire N__42378;
    wire N__42375;
    wire N__42374;
    wire N__42371;
    wire N__42368;
    wire N__42365;
    wire N__42362;
    wire N__42359;
    wire N__42356;
    wire N__42351;
    wire N__42346;
    wire N__42343;
    wire N__42340;
    wire N__42339;
    wire N__42336;
    wire N__42333;
    wire N__42328;
    wire N__42325;
    wire N__42322;
    wire N__42319;
    wire N__42316;
    wire N__42315;
    wire N__42312;
    wire N__42309;
    wire N__42306;
    wire N__42303;
    wire N__42298;
    wire N__42297;
    wire N__42294;
    wire N__42291;
    wire N__42288;
    wire N__42285;
    wire N__42282;
    wire N__42277;
    wire N__42274;
    wire N__42271;
    wire N__42270;
    wire N__42269;
    wire N__42266;
    wire N__42261;
    wire N__42256;
    wire N__42255;
    wire N__42252;
    wire N__42251;
    wire N__42248;
    wire N__42245;
    wire N__42240;
    wire N__42235;
    wire N__42234;
    wire N__42231;
    wire N__42228;
    wire N__42225;
    wire N__42224;
    wire N__42221;
    wire N__42218;
    wire N__42215;
    wire N__42208;
    wire N__42207;
    wire N__42206;
    wire N__42205;
    wire N__42204;
    wire N__42199;
    wire N__42198;
    wire N__42197;
    wire N__42194;
    wire N__42193;
    wire N__42192;
    wire N__42189;
    wire N__42186;
    wire N__42183;
    wire N__42180;
    wire N__42179;
    wire N__42176;
    wire N__42173;
    wire N__42172;
    wire N__42171;
    wire N__42170;
    wire N__42167;
    wire N__42166;
    wire N__42163;
    wire N__42162;
    wire N__42157;
    wire N__42156;
    wire N__42155;
    wire N__42150;
    wire N__42147;
    wire N__42144;
    wire N__42141;
    wire N__42138;
    wire N__42135;
    wire N__42132;
    wire N__42123;
    wire N__42120;
    wire N__42115;
    wire N__42106;
    wire N__42091;
    wire N__42090;
    wire N__42089;
    wire N__42084;
    wire N__42081;
    wire N__42080;
    wire N__42079;
    wire N__42078;
    wire N__42075;
    wire N__42072;
    wire N__42071;
    wire N__42068;
    wire N__42067;
    wire N__42064;
    wire N__42061;
    wire N__42056;
    wire N__42049;
    wire N__42044;
    wire N__42037;
    wire N__42034;
    wire N__42031;
    wire N__42028;
    wire N__42027;
    wire N__42024;
    wire N__42021;
    wire N__42016;
    wire N__42013;
    wire N__42010;
    wire N__42007;
    wire N__42004;
    wire N__42001;
    wire N__41998;
    wire N__41995;
    wire N__41992;
    wire N__41989;
    wire N__41988;
    wire N__41985;
    wire N__41984;
    wire N__41983;
    wire N__41982;
    wire N__41979;
    wire N__41976;
    wire N__41971;
    wire N__41966;
    wire N__41959;
    wire N__41956;
    wire N__41953;
    wire N__41950;
    wire N__41949;
    wire N__41946;
    wire N__41943;
    wire N__41940;
    wire N__41937;
    wire N__41932;
    wire N__41929;
    wire N__41926;
    wire N__41923;
    wire N__41920;
    wire N__41917;
    wire N__41914;
    wire N__41911;
    wire N__41908;
    wire N__41905;
    wire N__41902;
    wire N__41899;
    wire N__41896;
    wire N__41893;
    wire N__41890;
    wire N__41887;
    wire N__41884;
    wire N__41881;
    wire N__41880;
    wire N__41877;
    wire N__41874;
    wire N__41873;
    wire N__41870;
    wire N__41867;
    wire N__41864;
    wire N__41859;
    wire N__41858;
    wire N__41855;
    wire N__41852;
    wire N__41849;
    wire N__41842;
    wire N__41839;
    wire N__41836;
    wire N__41833;
    wire N__41830;
    wire N__41827;
    wire N__41824;
    wire N__41821;
    wire N__41818;
    wire N__41815;
    wire N__41812;
    wire N__41809;
    wire N__41806;
    wire N__41803;
    wire N__41800;
    wire N__41797;
    wire N__41794;
    wire N__41791;
    wire N__41790;
    wire N__41789;
    wire N__41788;
    wire N__41787;
    wire N__41786;
    wire N__41783;
    wire N__41780;
    wire N__41777;
    wire N__41776;
    wire N__41773;
    wire N__41772;
    wire N__41771;
    wire N__41766;
    wire N__41761;
    wire N__41760;
    wire N__41759;
    wire N__41758;
    wire N__41755;
    wire N__41752;
    wire N__41749;
    wire N__41744;
    wire N__41741;
    wire N__41738;
    wire N__41735;
    wire N__41732;
    wire N__41729;
    wire N__41722;
    wire N__41717;
    wire N__41704;
    wire N__41701;
    wire N__41698;
    wire N__41695;
    wire N__41692;
    wire N__41689;
    wire N__41686;
    wire N__41683;
    wire N__41680;
    wire N__41677;
    wire N__41674;
    wire N__41671;
    wire N__41668;
    wire N__41665;
    wire N__41662;
    wire N__41659;
    wire N__41656;
    wire N__41653;
    wire N__41650;
    wire N__41647;
    wire N__41644;
    wire N__41641;
    wire N__41638;
    wire N__41635;
    wire N__41632;
    wire N__41629;
    wire N__41628;
    wire N__41627;
    wire N__41624;
    wire N__41623;
    wire N__41620;
    wire N__41617;
    wire N__41614;
    wire N__41611;
    wire N__41608;
    wire N__41601;
    wire N__41596;
    wire N__41593;
    wire N__41590;
    wire N__41587;
    wire N__41584;
    wire N__41583;
    wire N__41580;
    wire N__41579;
    wire N__41574;
    wire N__41573;
    wire N__41572;
    wire N__41571;
    wire N__41568;
    wire N__41565;
    wire N__41558;
    wire N__41551;
    wire N__41548;
    wire N__41547;
    wire N__41544;
    wire N__41541;
    wire N__41538;
    wire N__41533;
    wire N__41530;
    wire N__41527;
    wire N__41524;
    wire N__41521;
    wire N__41518;
    wire N__41515;
    wire N__41512;
    wire N__41509;
    wire N__41506;
    wire N__41503;
    wire N__41500;
    wire N__41497;
    wire N__41494;
    wire N__41491;
    wire N__41488;
    wire N__41485;
    wire N__41482;
    wire N__41479;
    wire N__41476;
    wire N__41473;
    wire N__41470;
    wire N__41467;
    wire N__41464;
    wire N__41461;
    wire N__41458;
    wire N__41455;
    wire N__41452;
    wire N__41449;
    wire N__41446;
    wire N__41443;
    wire N__41440;
    wire N__41437;
    wire N__41434;
    wire N__41431;
    wire N__41428;
    wire N__41425;
    wire N__41422;
    wire N__41419;
    wire N__41416;
    wire N__41413;
    wire N__41410;
    wire N__41407;
    wire N__41404;
    wire N__41401;
    wire N__41400;
    wire N__41399;
    wire N__41398;
    wire N__41397;
    wire N__41396;
    wire N__41395;
    wire N__41392;
    wire N__41391;
    wire N__41390;
    wire N__41379;
    wire N__41376;
    wire N__41373;
    wire N__41368;
    wire N__41365;
    wire N__41356;
    wire N__41353;
    wire N__41350;
    wire N__41349;
    wire N__41348;
    wire N__41347;
    wire N__41346;
    wire N__41343;
    wire N__41332;
    wire N__41331;
    wire N__41330;
    wire N__41329;
    wire N__41326;
    wire N__41321;
    wire N__41318;
    wire N__41313;
    wire N__41308;
    wire N__41307;
    wire N__41306;
    wire N__41305;
    wire N__41302;
    wire N__41299;
    wire N__41292;
    wire N__41287;
    wire N__41286;
    wire N__41285;
    wire N__41284;
    wire N__41283;
    wire N__41280;
    wire N__41277;
    wire N__41274;
    wire N__41271;
    wire N__41268;
    wire N__41265;
    wire N__41262;
    wire N__41257;
    wire N__41254;
    wire N__41245;
    wire N__41242;
    wire N__41239;
    wire N__41238;
    wire N__41235;
    wire N__41232;
    wire N__41227;
    wire N__41226;
    wire N__41223;
    wire N__41220;
    wire N__41219;
    wire N__41218;
    wire N__41217;
    wire N__41212;
    wire N__41209;
    wire N__41204;
    wire N__41197;
    wire N__41194;
    wire N__41193;
    wire N__41188;
    wire N__41185;
    wire N__41182;
    wire N__41179;
    wire N__41176;
    wire N__41173;
    wire N__41172;
    wire N__41169;
    wire N__41166;
    wire N__41161;
    wire N__41158;
    wire N__41157;
    wire N__41156;
    wire N__41153;
    wire N__41150;
    wire N__41147;
    wire N__41142;
    wire N__41137;
    wire N__41134;
    wire N__41131;
    wire N__41128;
    wire N__41125;
    wire N__41122;
    wire N__41119;
    wire N__41118;
    wire N__41117;
    wire N__41116;
    wire N__41113;
    wire N__41108;
    wire N__41103;
    wire N__41098;
    wire N__41095;
    wire N__41092;
    wire N__41089;
    wire N__41086;
    wire N__41083;
    wire N__41080;
    wire N__41077;
    wire N__41074;
    wire N__41071;
    wire N__41068;
    wire N__41065;
    wire N__41062;
    wire N__41059;
    wire N__41056;
    wire N__41055;
    wire N__41050;
    wire N__41047;
    wire N__41044;
    wire N__41041;
    wire N__41038;
    wire N__41035;
    wire N__41032;
    wire N__41029;
    wire N__41026;
    wire N__41023;
    wire N__41020;
    wire N__41019;
    wire N__41018;
    wire N__41015;
    wire N__41012;
    wire N__41007;
    wire N__41002;
    wire N__40999;
    wire N__40996;
    wire N__40993;
    wire N__40990;
    wire N__40987;
    wire N__40984;
    wire N__40981;
    wire N__40978;
    wire N__40977;
    wire N__40976;
    wire N__40969;
    wire N__40966;
    wire N__40963;
    wire N__40960;
    wire N__40957;
    wire N__40954;
    wire N__40951;
    wire N__40948;
    wire N__40945;
    wire N__40942;
    wire N__40941;
    wire N__40938;
    wire N__40935;
    wire N__40930;
    wire N__40927;
    wire N__40924;
    wire N__40921;
    wire N__40920;
    wire N__40917;
    wire N__40914;
    wire N__40911;
    wire N__40908;
    wire N__40905;
    wire N__40900;
    wire N__40897;
    wire N__40894;
    wire N__40891;
    wire N__40888;
    wire N__40885;
    wire N__40882;
    wire N__40879;
    wire N__40876;
    wire N__40873;
    wire N__40870;
    wire N__40867;
    wire N__40864;
    wire N__40861;
    wire N__40858;
    wire N__40855;
    wire N__40854;
    wire N__40851;
    wire N__40848;
    wire N__40845;
    wire N__40842;
    wire N__40837;
    wire N__40834;
    wire N__40831;
    wire N__40830;
    wire N__40829;
    wire N__40824;
    wire N__40821;
    wire N__40818;
    wire N__40813;
    wire N__40810;
    wire N__40809;
    wire N__40808;
    wire N__40805;
    wire N__40802;
    wire N__40799;
    wire N__40796;
    wire N__40793;
    wire N__40790;
    wire N__40787;
    wire N__40784;
    wire N__40777;
    wire N__40776;
    wire N__40775;
    wire N__40772;
    wire N__40769;
    wire N__40766;
    wire N__40763;
    wire N__40758;
    wire N__40755;
    wire N__40752;
    wire N__40747;
    wire N__40744;
    wire N__40741;
    wire N__40738;
    wire N__40735;
    wire N__40732;
    wire N__40729;
    wire N__40726;
    wire N__40723;
    wire N__40720;
    wire N__40717;
    wire N__40714;
    wire N__40711;
    wire N__40708;
    wire N__40705;
    wire N__40702;
    wire N__40699;
    wire N__40696;
    wire N__40693;
    wire N__40692;
    wire N__40689;
    wire N__40686;
    wire N__40685;
    wire N__40682;
    wire N__40679;
    wire N__40676;
    wire N__40673;
    wire N__40670;
    wire N__40663;
    wire N__40660;
    wire N__40657;
    wire N__40654;
    wire N__40651;
    wire N__40650;
    wire N__40649;
    wire N__40646;
    wire N__40643;
    wire N__40640;
    wire N__40637;
    wire N__40634;
    wire N__40631;
    wire N__40628;
    wire N__40623;
    wire N__40620;
    wire N__40615;
    wire N__40612;
    wire N__40609;
    wire N__40606;
    wire N__40603;
    wire N__40600;
    wire N__40597;
    wire N__40594;
    wire N__40591;
    wire N__40588;
    wire N__40585;
    wire N__40582;
    wire N__40579;
    wire N__40576;
    wire N__40573;
    wire N__40570;
    wire N__40567;
    wire N__40564;
    wire N__40563;
    wire N__40558;
    wire N__40557;
    wire N__40554;
    wire N__40551;
    wire N__40546;
    wire N__40543;
    wire N__40540;
    wire N__40537;
    wire N__40534;
    wire N__40531;
    wire N__40530;
    wire N__40527;
    wire N__40524;
    wire N__40521;
    wire N__40516;
    wire N__40515;
    wire N__40514;
    wire N__40513;
    wire N__40512;
    wire N__40511;
    wire N__40510;
    wire N__40509;
    wire N__40508;
    wire N__40507;
    wire N__40506;
    wire N__40505;
    wire N__40504;
    wire N__40503;
    wire N__40502;
    wire N__40501;
    wire N__40500;
    wire N__40499;
    wire N__40498;
    wire N__40497;
    wire N__40496;
    wire N__40495;
    wire N__40450;
    wire N__40447;
    wire N__40444;
    wire N__40441;
    wire N__40438;
    wire N__40435;
    wire N__40432;
    wire N__40429;
    wire N__40426;
    wire N__40423;
    wire N__40420;
    wire N__40417;
    wire N__40416;
    wire N__40415;
    wire N__40412;
    wire N__40411;
    wire N__40408;
    wire N__40405;
    wire N__40402;
    wire N__40399;
    wire N__40396;
    wire N__40391;
    wire N__40386;
    wire N__40381;
    wire N__40380;
    wire N__40377;
    wire N__40374;
    wire N__40373;
    wire N__40366;
    wire N__40363;
    wire N__40362;
    wire N__40359;
    wire N__40356;
    wire N__40353;
    wire N__40348;
    wire N__40345;
    wire N__40342;
    wire N__40339;
    wire N__40336;
    wire N__40333;
    wire N__40330;
    wire N__40327;
    wire N__40324;
    wire N__40321;
    wire N__40318;
    wire N__40315;
    wire N__40312;
    wire N__40309;
    wire N__40306;
    wire N__40303;
    wire N__40300;
    wire N__40297;
    wire N__40296;
    wire N__40293;
    wire N__40290;
    wire N__40287;
    wire N__40284;
    wire N__40281;
    wire N__40278;
    wire N__40275;
    wire N__40272;
    wire N__40267;
    wire N__40264;
    wire N__40263;
    wire N__40260;
    wire N__40257;
    wire N__40252;
    wire N__40249;
    wire N__40246;
    wire N__40243;
    wire N__40240;
    wire N__40237;
    wire N__40234;
    wire N__40231;
    wire N__40228;
    wire N__40225;
    wire N__40222;
    wire N__40219;
    wire N__40218;
    wire N__40217;
    wire N__40216;
    wire N__40213;
    wire N__40208;
    wire N__40205;
    wire N__40200;
    wire N__40197;
    wire N__40192;
    wire N__40191;
    wire N__40188;
    wire N__40185;
    wire N__40182;
    wire N__40179;
    wire N__40176;
    wire N__40171;
    wire N__40170;
    wire N__40167;
    wire N__40164;
    wire N__40163;
    wire N__40162;
    wire N__40157;
    wire N__40152;
    wire N__40147;
    wire N__40144;
    wire N__40141;
    wire N__40138;
    wire N__40135;
    wire N__40132;
    wire N__40129;
    wire N__40128;
    wire N__40125;
    wire N__40122;
    wire N__40119;
    wire N__40114;
    wire N__40111;
    wire N__40108;
    wire N__40105;
    wire N__40104;
    wire N__40101;
    wire N__40098;
    wire N__40093;
    wire N__40092;
    wire N__40089;
    wire N__40086;
    wire N__40083;
    wire N__40078;
    wire N__40077;
    wire N__40074;
    wire N__40071;
    wire N__40068;
    wire N__40065;
    wire N__40062;
    wire N__40057;
    wire N__40056;
    wire N__40055;
    wire N__40048;
    wire N__40045;
    wire N__40042;
    wire N__40039;
    wire N__40036;
    wire N__40033;
    wire N__40030;
    wire N__40029;
    wire N__40024;
    wire N__40021;
    wire N__40020;
    wire N__40015;
    wire N__40012;
    wire N__40009;
    wire N__40006;
    wire N__40003;
    wire N__40000;
    wire N__39997;
    wire N__39994;
    wire N__39993;
    wire N__39990;
    wire N__39987;
    wire N__39984;
    wire N__39981;
    wire N__39976;
    wire N__39975;
    wire N__39970;
    wire N__39967;
    wire N__39964;
    wire N__39961;
    wire N__39958;
    wire N__39957;
    wire N__39956;
    wire N__39953;
    wire N__39948;
    wire N__39945;
    wire N__39942;
    wire N__39939;
    wire N__39936;
    wire N__39931;
    wire N__39928;
    wire N__39925;
    wire N__39922;
    wire N__39919;
    wire N__39916;
    wire N__39913;
    wire N__39910;
    wire N__39907;
    wire N__39904;
    wire N__39901;
    wire N__39898;
    wire N__39895;
    wire N__39892;
    wire N__39889;
    wire N__39886;
    wire N__39883;
    wire N__39880;
    wire N__39877;
    wire N__39874;
    wire N__39871;
    wire N__39870;
    wire N__39869;
    wire N__39868;
    wire N__39867;
    wire N__39862;
    wire N__39859;
    wire N__39854;
    wire N__39847;
    wire N__39844;
    wire N__39843;
    wire N__39840;
    wire N__39837;
    wire N__39834;
    wire N__39831;
    wire N__39826;
    wire N__39823;
    wire N__39822;
    wire N__39817;
    wire N__39814;
    wire N__39811;
    wire N__39808;
    wire N__39805;
    wire N__39804;
    wire N__39801;
    wire N__39798;
    wire N__39793;
    wire N__39790;
    wire N__39787;
    wire N__39786;
    wire N__39785;
    wire N__39782;
    wire N__39781;
    wire N__39780;
    wire N__39777;
    wire N__39776;
    wire N__39773;
    wire N__39772;
    wire N__39769;
    wire N__39768;
    wire N__39767;
    wire N__39766;
    wire N__39755;
    wire N__39752;
    wire N__39749;
    wire N__39742;
    wire N__39739;
    wire N__39736;
    wire N__39727;
    wire N__39724;
    wire N__39723;
    wire N__39722;
    wire N__39719;
    wire N__39716;
    wire N__39715;
    wire N__39714;
    wire N__39711;
    wire N__39708;
    wire N__39707;
    wire N__39704;
    wire N__39699;
    wire N__39694;
    wire N__39691;
    wire N__39686;
    wire N__39683;
    wire N__39676;
    wire N__39675;
    wire N__39674;
    wire N__39673;
    wire N__39670;
    wire N__39669;
    wire N__39668;
    wire N__39667;
    wire N__39666;
    wire N__39665;
    wire N__39664;
    wire N__39663;
    wire N__39656;
    wire N__39653;
    wire N__39642;
    wire N__39637;
    wire N__39628;
    wire N__39627;
    wire N__39624;
    wire N__39621;
    wire N__39618;
    wire N__39615;
    wire N__39612;
    wire N__39609;
    wire N__39604;
    wire N__39601;
    wire N__39598;
    wire N__39595;
    wire N__39594;
    wire N__39593;
    wire N__39590;
    wire N__39587;
    wire N__39584;
    wire N__39579;
    wire N__39576;
    wire N__39573;
    wire N__39568;
    wire N__39567;
    wire N__39566;
    wire N__39563;
    wire N__39560;
    wire N__39557;
    wire N__39556;
    wire N__39553;
    wire N__39550;
    wire N__39547;
    wire N__39544;
    wire N__39541;
    wire N__39538;
    wire N__39535;
    wire N__39532;
    wire N__39523;
    wire N__39520;
    wire N__39517;
    wire N__39516;
    wire N__39513;
    wire N__39510;
    wire N__39507;
    wire N__39504;
    wire N__39501;
    wire N__39498;
    wire N__39495;
    wire N__39490;
    wire N__39487;
    wire N__39486;
    wire N__39483;
    wire N__39480;
    wire N__39477;
    wire N__39472;
    wire N__39471;
    wire N__39466;
    wire N__39465;
    wire N__39462;
    wire N__39459;
    wire N__39454;
    wire N__39451;
    wire N__39448;
    wire N__39445;
    wire N__39442;
    wire N__39439;
    wire N__39436;
    wire N__39433;
    wire N__39432;
    wire N__39431;
    wire N__39428;
    wire N__39423;
    wire N__39420;
    wire N__39417;
    wire N__39414;
    wire N__39411;
    wire N__39406;
    wire N__39403;
    wire N__39402;
    wire N__39399;
    wire N__39396;
    wire N__39393;
    wire N__39390;
    wire N__39385;
    wire N__39384;
    wire N__39379;
    wire N__39376;
    wire N__39373;
    wire N__39372;
    wire N__39371;
    wire N__39366;
    wire N__39363;
    wire N__39360;
    wire N__39357;
    wire N__39352;
    wire N__39351;
    wire N__39350;
    wire N__39345;
    wire N__39342;
    wire N__39339;
    wire N__39336;
    wire N__39331;
    wire N__39330;
    wire N__39329;
    wire N__39326;
    wire N__39323;
    wire N__39318;
    wire N__39315;
    wire N__39312;
    wire N__39309;
    wire N__39304;
    wire N__39303;
    wire N__39298;
    wire N__39297;
    wire N__39294;
    wire N__39291;
    wire N__39286;
    wire N__39285;
    wire N__39284;
    wire N__39279;
    wire N__39276;
    wire N__39271;
    wire N__39268;
    wire N__39265;
    wire N__39264;
    wire N__39263;
    wire N__39258;
    wire N__39255;
    wire N__39252;
    wire N__39249;
    wire N__39244;
    wire N__39243;
    wire N__39240;
    wire N__39237;
    wire N__39232;
    wire N__39229;
    wire N__39228;
    wire N__39223;
    wire N__39220;
    wire N__39217;
    wire N__39214;
    wire N__39211;
    wire N__39208;
    wire N__39205;
    wire N__39202;
    wire N__39199;
    wire N__39196;
    wire N__39193;
    wire N__39190;
    wire N__39187;
    wire N__39184;
    wire N__39181;
    wire N__39178;
    wire N__39175;
    wire N__39172;
    wire N__39169;
    wire N__39166;
    wire N__39163;
    wire N__39160;
    wire N__39157;
    wire N__39154;
    wire N__39151;
    wire N__39148;
    wire N__39145;
    wire N__39142;
    wire N__39139;
    wire N__39136;
    wire N__39133;
    wire N__39130;
    wire N__39127;
    wire N__39124;
    wire N__39121;
    wire N__39118;
    wire N__39115;
    wire N__39112;
    wire N__39109;
    wire N__39106;
    wire N__39103;
    wire N__39100;
    wire N__39097;
    wire N__39094;
    wire N__39091;
    wire N__39088;
    wire N__39085;
    wire N__39082;
    wire N__39079;
    wire N__39076;
    wire N__39075;
    wire N__39072;
    wire N__39069;
    wire N__39066;
    wire N__39063;
    wire N__39058;
    wire N__39055;
    wire N__39052;
    wire N__39049;
    wire N__39046;
    wire N__39043;
    wire N__39042;
    wire N__39041;
    wire N__39038;
    wire N__39035;
    wire N__39032;
    wire N__39029;
    wire N__39022;
    wire N__39019;
    wire N__39016;
    wire N__39013;
    wire N__39010;
    wire N__39007;
    wire N__39004;
    wire N__39001;
    wire N__38998;
    wire N__38995;
    wire N__38994;
    wire N__38991;
    wire N__38990;
    wire N__38983;
    wire N__38980;
    wire N__38977;
    wire N__38974;
    wire N__38971;
    wire N__38968;
    wire N__38965;
    wire N__38962;
    wire N__38959;
    wire N__38956;
    wire N__38953;
    wire N__38952;
    wire N__38951;
    wire N__38950;
    wire N__38949;
    wire N__38948;
    wire N__38947;
    wire N__38944;
    wire N__38941;
    wire N__38938;
    wire N__38933;
    wire N__38928;
    wire N__38917;
    wire N__38916;
    wire N__38915;
    wire N__38914;
    wire N__38911;
    wire N__38904;
    wire N__38899;
    wire N__38898;
    wire N__38897;
    wire N__38896;
    wire N__38893;
    wire N__38886;
    wire N__38881;
    wire N__38878;
    wire N__38875;
    wire N__38872;
    wire N__38869;
    wire N__38866;
    wire N__38865;
    wire N__38862;
    wire N__38861;
    wire N__38858;
    wire N__38855;
    wire N__38852;
    wire N__38849;
    wire N__38846;
    wire N__38843;
    wire N__38840;
    wire N__38837;
    wire N__38830;
    wire N__38827;
    wire N__38824;
    wire N__38823;
    wire N__38820;
    wire N__38817;
    wire N__38812;
    wire N__38809;
    wire N__38808;
    wire N__38807;
    wire N__38806;
    wire N__38805;
    wire N__38804;
    wire N__38795;
    wire N__38792;
    wire N__38789;
    wire N__38782;
    wire N__38779;
    wire N__38776;
    wire N__38773;
    wire N__38772;
    wire N__38769;
    wire N__38766;
    wire N__38763;
    wire N__38760;
    wire N__38757;
    wire N__38754;
    wire N__38751;
    wire N__38748;
    wire N__38743;
    wire N__38742;
    wire N__38739;
    wire N__38736;
    wire N__38733;
    wire N__38730;
    wire N__38725;
    wire N__38722;
    wire N__38721;
    wire N__38718;
    wire N__38715;
    wire N__38710;
    wire N__38707;
    wire N__38704;
    wire N__38701;
    wire N__38700;
    wire N__38699;
    wire N__38696;
    wire N__38691;
    wire N__38686;
    wire N__38683;
    wire N__38682;
    wire N__38679;
    wire N__38676;
    wire N__38675;
    wire N__38672;
    wire N__38669;
    wire N__38666;
    wire N__38659;
    wire N__38658;
    wire N__38657;
    wire N__38652;
    wire N__38649;
    wire N__38646;
    wire N__38641;
    wire N__38638;
    wire N__38635;
    wire N__38634;
    wire N__38633;
    wire N__38630;
    wire N__38625;
    wire N__38620;
    wire N__38617;
    wire N__38616;
    wire N__38615;
    wire N__38612;
    wire N__38609;
    wire N__38608;
    wire N__38605;
    wire N__38602;
    wire N__38599;
    wire N__38596;
    wire N__38593;
    wire N__38590;
    wire N__38587;
    wire N__38584;
    wire N__38581;
    wire N__38580;
    wire N__38571;
    wire N__38568;
    wire N__38563;
    wire N__38560;
    wire N__38557;
    wire N__38554;
    wire N__38551;
    wire N__38548;
    wire N__38545;
    wire N__38544;
    wire N__38543;
    wire N__38540;
    wire N__38537;
    wire N__38534;
    wire N__38529;
    wire N__38526;
    wire N__38523;
    wire N__38520;
    wire N__38517;
    wire N__38514;
    wire N__38509;
    wire N__38506;
    wire N__38505;
    wire N__38504;
    wire N__38501;
    wire N__38498;
    wire N__38495;
    wire N__38492;
    wire N__38489;
    wire N__38486;
    wire N__38483;
    wire N__38480;
    wire N__38477;
    wire N__38474;
    wire N__38471;
    wire N__38464;
    wire N__38461;
    wire N__38458;
    wire N__38455;
    wire N__38454;
    wire N__38453;
    wire N__38450;
    wire N__38447;
    wire N__38444;
    wire N__38439;
    wire N__38436;
    wire N__38433;
    wire N__38430;
    wire N__38427;
    wire N__38424;
    wire N__38419;
    wire N__38416;
    wire N__38413;
    wire N__38410;
    wire N__38409;
    wire N__38408;
    wire N__38405;
    wire N__38402;
    wire N__38399;
    wire N__38394;
    wire N__38391;
    wire N__38388;
    wire N__38385;
    wire N__38382;
    wire N__38379;
    wire N__38374;
    wire N__38371;
    wire N__38368;
    wire N__38367;
    wire N__38366;
    wire N__38363;
    wire N__38360;
    wire N__38357;
    wire N__38354;
    wire N__38351;
    wire N__38348;
    wire N__38345;
    wire N__38342;
    wire N__38339;
    wire N__38334;
    wire N__38331;
    wire N__38326;
    wire N__38323;
    wire N__38320;
    wire N__38319;
    wire N__38318;
    wire N__38315;
    wire N__38312;
    wire N__38309;
    wire N__38306;
    wire N__38303;
    wire N__38300;
    wire N__38297;
    wire N__38294;
    wire N__38291;
    wire N__38286;
    wire N__38283;
    wire N__38278;
    wire N__38275;
    wire N__38272;
    wire N__38271;
    wire N__38270;
    wire N__38267;
    wire N__38264;
    wire N__38261;
    wire N__38258;
    wire N__38255;
    wire N__38252;
    wire N__38249;
    wire N__38246;
    wire N__38243;
    wire N__38238;
    wire N__38235;
    wire N__38230;
    wire N__38227;
    wire N__38226;
    wire N__38223;
    wire N__38222;
    wire N__38219;
    wire N__38216;
    wire N__38213;
    wire N__38210;
    wire N__38207;
    wire N__38204;
    wire N__38201;
    wire N__38198;
    wire N__38195;
    wire N__38192;
    wire N__38185;
    wire N__38182;
    wire N__38179;
    wire N__38176;
    wire N__38173;
    wire N__38172;
    wire N__38171;
    wire N__38168;
    wire N__38165;
    wire N__38162;
    wire N__38157;
    wire N__38154;
    wire N__38151;
    wire N__38148;
    wire N__38145;
    wire N__38142;
    wire N__38137;
    wire N__38134;
    wire N__38131;
    wire N__38130;
    wire N__38127;
    wire N__38124;
    wire N__38123;
    wire N__38120;
    wire N__38117;
    wire N__38114;
    wire N__38107;
    wire N__38106;
    wire N__38105;
    wire N__38102;
    wire N__38099;
    wire N__38096;
    wire N__38093;
    wire N__38086;
    wire N__38083;
    wire N__38082;
    wire N__38081;
    wire N__38078;
    wire N__38075;
    wire N__38072;
    wire N__38069;
    wire N__38066;
    wire N__38061;
    wire N__38058;
    wire N__38055;
    wire N__38052;
    wire N__38047;
    wire N__38044;
    wire N__38041;
    wire N__38038;
    wire N__38035;
    wire N__38034;
    wire N__38031;
    wire N__38028;
    wire N__38027;
    wire N__38022;
    wire N__38019;
    wire N__38016;
    wire N__38013;
    wire N__38010;
    wire N__38007;
    wire N__38002;
    wire N__37999;
    wire N__37996;
    wire N__37993;
    wire N__37990;
    wire N__37989;
    wire N__37988;
    wire N__37985;
    wire N__37982;
    wire N__37979;
    wire N__37974;
    wire N__37971;
    wire N__37968;
    wire N__37965;
    wire N__37962;
    wire N__37959;
    wire N__37954;
    wire N__37951;
    wire N__37948;
    wire N__37947;
    wire N__37946;
    wire N__37943;
    wire N__37940;
    wire N__37937;
    wire N__37934;
    wire N__37931;
    wire N__37928;
    wire N__37925;
    wire N__37922;
    wire N__37919;
    wire N__37914;
    wire N__37911;
    wire N__37906;
    wire N__37903;
    wire N__37900;
    wire N__37897;
    wire N__37896;
    wire N__37895;
    wire N__37892;
    wire N__37889;
    wire N__37886;
    wire N__37883;
    wire N__37880;
    wire N__37877;
    wire N__37872;
    wire N__37869;
    wire N__37866;
    wire N__37863;
    wire N__37858;
    wire N__37855;
    wire N__37852;
    wire N__37849;
    wire N__37848;
    wire N__37847;
    wire N__37844;
    wire N__37841;
    wire N__37838;
    wire N__37833;
    wire N__37830;
    wire N__37827;
    wire N__37824;
    wire N__37821;
    wire N__37818;
    wire N__37813;
    wire N__37810;
    wire N__37807;
    wire N__37806;
    wire N__37803;
    wire N__37802;
    wire N__37799;
    wire N__37796;
    wire N__37793;
    wire N__37790;
    wire N__37787;
    wire N__37784;
    wire N__37781;
    wire N__37776;
    wire N__37773;
    wire N__37768;
    wire N__37765;
    wire N__37764;
    wire N__37763;
    wire N__37760;
    wire N__37755;
    wire N__37752;
    wire N__37749;
    wire N__37744;
    wire N__37741;
    wire N__37738;
    wire N__37737;
    wire N__37736;
    wire N__37733;
    wire N__37728;
    wire N__37723;
    wire N__37720;
    wire N__37717;
    wire N__37714;
    wire N__37711;
    wire N__37708;
    wire N__37705;
    wire N__37702;
    wire N__37699;
    wire N__37698;
    wire N__37695;
    wire N__37692;
    wire N__37689;
    wire N__37686;
    wire N__37683;
    wire N__37678;
    wire N__37675;
    wire N__37672;
    wire N__37669;
    wire N__37668;
    wire N__37665;
    wire N__37662;
    wire N__37659;
    wire N__37656;
    wire N__37653;
    wire N__37650;
    wire N__37645;
    wire N__37644;
    wire N__37639;
    wire N__37636;
    wire N__37635;
    wire N__37634;
    wire N__37631;
    wire N__37626;
    wire N__37623;
    wire N__37620;
    wire N__37615;
    wire N__37612;
    wire N__37609;
    wire N__37606;
    wire N__37605;
    wire N__37602;
    wire N__37599;
    wire N__37594;
    wire N__37593;
    wire N__37592;
    wire N__37585;
    wire N__37582;
    wire N__37579;
    wire N__37576;
    wire N__37573;
    wire N__37570;
    wire N__37567;
    wire N__37566;
    wire N__37563;
    wire N__37560;
    wire N__37557;
    wire N__37554;
    wire N__37551;
    wire N__37548;
    wire N__37545;
    wire N__37540;
    wire N__37537;
    wire N__37534;
    wire N__37531;
    wire N__37528;
    wire N__37525;
    wire N__37522;
    wire N__37521;
    wire N__37518;
    wire N__37515;
    wire N__37512;
    wire N__37507;
    wire N__37504;
    wire N__37501;
    wire N__37498;
    wire N__37495;
    wire N__37492;
    wire N__37491;
    wire N__37488;
    wire N__37485;
    wire N__37482;
    wire N__37477;
    wire N__37474;
    wire N__37471;
    wire N__37468;
    wire N__37465;
    wire N__37462;
    wire N__37459;
    wire N__37456;
    wire N__37453;
    wire N__37450;
    wire N__37447;
    wire N__37444;
    wire N__37441;
    wire N__37438;
    wire N__37435;
    wire N__37432;
    wire N__37431;
    wire N__37428;
    wire N__37425;
    wire N__37422;
    wire N__37419;
    wire N__37416;
    wire N__37413;
    wire N__37410;
    wire N__37405;
    wire N__37402;
    wire N__37399;
    wire N__37396;
    wire N__37393;
    wire N__37390;
    wire N__37387;
    wire N__37384;
    wire N__37381;
    wire N__37378;
    wire N__37375;
    wire N__37372;
    wire N__37369;
    wire N__37366;
    wire N__37365;
    wire N__37364;
    wire N__37361;
    wire N__37356;
    wire N__37351;
    wire N__37350;
    wire N__37345;
    wire N__37342;
    wire N__37339;
    wire N__37336;
    wire N__37333;
    wire N__37330;
    wire N__37327;
    wire N__37324;
    wire N__37321;
    wire N__37318;
    wire N__37315;
    wire N__37312;
    wire N__37309;
    wire N__37306;
    wire N__37303;
    wire N__37300;
    wire N__37299;
    wire N__37296;
    wire N__37293;
    wire N__37290;
    wire N__37285;
    wire N__37282;
    wire N__37279;
    wire N__37276;
    wire N__37275;
    wire N__37272;
    wire N__37269;
    wire N__37266;
    wire N__37263;
    wire N__37260;
    wire N__37257;
    wire N__37254;
    wire N__37249;
    wire N__37246;
    wire N__37243;
    wire N__37240;
    wire N__37239;
    wire N__37236;
    wire N__37233;
    wire N__37230;
    wire N__37227;
    wire N__37222;
    wire N__37219;
    wire N__37216;
    wire N__37213;
    wire N__37210;
    wire N__37209;
    wire N__37206;
    wire N__37203;
    wire N__37200;
    wire N__37195;
    wire N__37192;
    wire N__37189;
    wire N__37186;
    wire N__37183;
    wire N__37182;
    wire N__37179;
    wire N__37176;
    wire N__37173;
    wire N__37170;
    wire N__37165;
    wire N__37162;
    wire N__37159;
    wire N__37156;
    wire N__37153;
    wire N__37150;
    wire N__37147;
    wire N__37144;
    wire N__37143;
    wire N__37140;
    wire N__37137;
    wire N__37134;
    wire N__37131;
    wire N__37126;
    wire N__37123;
    wire N__37122;
    wire N__37119;
    wire N__37116;
    wire N__37113;
    wire N__37110;
    wire N__37107;
    wire N__37102;
    wire N__37099;
    wire N__37096;
    wire N__37093;
    wire N__37090;
    wire N__37087;
    wire N__37084;
    wire N__37081;
    wire N__37078;
    wire N__37075;
    wire N__37072;
    wire N__37071;
    wire N__37070;
    wire N__37067;
    wire N__37064;
    wire N__37061;
    wire N__37058;
    wire N__37055;
    wire N__37052;
    wire N__37049;
    wire N__37042;
    wire N__37041;
    wire N__37038;
    wire N__37035;
    wire N__37030;
    wire N__37027;
    wire N__37024;
    wire N__37021;
    wire N__37020;
    wire N__37017;
    wire N__37014;
    wire N__37013;
    wire N__37010;
    wire N__37007;
    wire N__37004;
    wire N__37001;
    wire N__36998;
    wire N__36995;
    wire N__36992;
    wire N__36985;
    wire N__36984;
    wire N__36981;
    wire N__36978;
    wire N__36975;
    wire N__36972;
    wire N__36967;
    wire N__36964;
    wire N__36961;
    wire N__36958;
    wire N__36957;
    wire N__36954;
    wire N__36951;
    wire N__36946;
    wire N__36943;
    wire N__36940;
    wire N__36937;
    wire N__36934;
    wire N__36931;
    wire N__36928;
    wire N__36927;
    wire N__36924;
    wire N__36921;
    wire N__36918;
    wire N__36913;
    wire N__36910;
    wire N__36907;
    wire N__36904;
    wire N__36903;
    wire N__36900;
    wire N__36897;
    wire N__36894;
    wire N__36891;
    wire N__36886;
    wire N__36883;
    wire N__36880;
    wire N__36877;
    wire N__36874;
    wire N__36871;
    wire N__36870;
    wire N__36867;
    wire N__36864;
    wire N__36861;
    wire N__36858;
    wire N__36853;
    wire N__36850;
    wire N__36847;
    wire N__36846;
    wire N__36843;
    wire N__36840;
    wire N__36835;
    wire N__36832;
    wire N__36831;
    wire N__36828;
    wire N__36827;
    wire N__36820;
    wire N__36817;
    wire N__36816;
    wire N__36813;
    wire N__36810;
    wire N__36805;
    wire N__36802;
    wire N__36799;
    wire N__36796;
    wire N__36795;
    wire N__36792;
    wire N__36789;
    wire N__36786;
    wire N__36783;
    wire N__36778;
    wire N__36775;
    wire N__36772;
    wire N__36769;
    wire N__36766;
    wire N__36763;
    wire N__36762;
    wire N__36759;
    wire N__36756;
    wire N__36753;
    wire N__36750;
    wire N__36747;
    wire N__36744;
    wire N__36741;
    wire N__36736;
    wire N__36735;
    wire N__36730;
    wire N__36727;
    wire N__36724;
    wire N__36721;
    wire N__36718;
    wire N__36715;
    wire N__36712;
    wire N__36711;
    wire N__36706;
    wire N__36703;
    wire N__36700;
    wire N__36697;
    wire N__36696;
    wire N__36693;
    wire N__36692;
    wire N__36689;
    wire N__36686;
    wire N__36683;
    wire N__36676;
    wire N__36675;
    wire N__36672;
    wire N__36671;
    wire N__36668;
    wire N__36665;
    wire N__36662;
    wire N__36659;
    wire N__36656;
    wire N__36649;
    wire N__36648;
    wire N__36645;
    wire N__36644;
    wire N__36643;
    wire N__36642;
    wire N__36639;
    wire N__36638;
    wire N__36625;
    wire N__36622;
    wire N__36619;
    wire N__36616;
    wire N__36613;
    wire N__36610;
    wire N__36607;
    wire N__36604;
    wire N__36601;
    wire N__36598;
    wire N__36595;
    wire N__36592;
    wire N__36589;
    wire N__36586;
    wire N__36583;
    wire N__36580;
    wire N__36577;
    wire N__36574;
    wire N__36571;
    wire N__36568;
    wire N__36567;
    wire N__36564;
    wire N__36561;
    wire N__36560;
    wire N__36557;
    wire N__36554;
    wire N__36551;
    wire N__36544;
    wire N__36541;
    wire N__36540;
    wire N__36537;
    wire N__36534;
    wire N__36531;
    wire N__36526;
    wire N__36523;
    wire N__36520;
    wire N__36517;
    wire N__36514;
    wire N__36511;
    wire N__36508;
    wire N__36505;
    wire N__36502;
    wire N__36499;
    wire N__36496;
    wire N__36493;
    wire N__36490;
    wire N__36487;
    wire N__36484;
    wire N__36481;
    wire N__36478;
    wire N__36475;
    wire N__36472;
    wire N__36469;
    wire N__36466;
    wire N__36463;
    wire N__36460;
    wire N__36457;
    wire N__36454;
    wire N__36451;
    wire N__36450;
    wire N__36449;
    wire N__36446;
    wire N__36443;
    wire N__36440;
    wire N__36435;
    wire N__36430;
    wire N__36429;
    wire N__36426;
    wire N__36423;
    wire N__36420;
    wire N__36415;
    wire N__36414;
    wire N__36411;
    wire N__36410;
    wire N__36405;
    wire N__36402;
    wire N__36399;
    wire N__36396;
    wire N__36393;
    wire N__36388;
    wire N__36385;
    wire N__36382;
    wire N__36379;
    wire N__36376;
    wire N__36373;
    wire N__36370;
    wire N__36367;
    wire N__36364;
    wire N__36361;
    wire N__36358;
    wire N__36355;
    wire N__36352;
    wire N__36349;
    wire N__36346;
    wire N__36343;
    wire N__36340;
    wire N__36337;
    wire N__36334;
    wire N__36331;
    wire N__36328;
    wire N__36325;
    wire N__36322;
    wire N__36319;
    wire N__36316;
    wire N__36313;
    wire N__36310;
    wire N__36307;
    wire N__36304;
    wire N__36301;
    wire N__36298;
    wire N__36295;
    wire N__36292;
    wire N__36289;
    wire N__36286;
    wire N__36283;
    wire N__36280;
    wire N__36277;
    wire N__36274;
    wire N__36271;
    wire N__36268;
    wire N__36265;
    wire N__36262;
    wire N__36259;
    wire N__36256;
    wire N__36253;
    wire N__36250;
    wire N__36247;
    wire N__36244;
    wire N__36241;
    wire N__36238;
    wire N__36237;
    wire N__36232;
    wire N__36229;
    wire N__36226;
    wire N__36225;
    wire N__36224;
    wire N__36221;
    wire N__36216;
    wire N__36213;
    wire N__36210;
    wire N__36205;
    wire N__36202;
    wire N__36199;
    wire N__36198;
    wire N__36197;
    wire N__36194;
    wire N__36189;
    wire N__36184;
    wire N__36181;
    wire N__36180;
    wire N__36175;
    wire N__36172;
    wire N__36169;
    wire N__36166;
    wire N__36165;
    wire N__36164;
    wire N__36161;
    wire N__36156;
    wire N__36151;
    wire N__36150;
    wire N__36145;
    wire N__36142;
    wire N__36139;
    wire N__36138;
    wire N__36137;
    wire N__36134;
    wire N__36129;
    wire N__36124;
    wire N__36121;
    wire N__36118;
    wire N__36115;
    wire N__36114;
    wire N__36113;
    wire N__36110;
    wire N__36105;
    wire N__36100;
    wire N__36097;
    wire N__36096;
    wire N__36095;
    wire N__36092;
    wire N__36087;
    wire N__36082;
    wire N__36079;
    wire N__36076;
    wire N__36075;
    wire N__36072;
    wire N__36069;
    wire N__36064;
    wire N__36061;
    wire N__36060;
    wire N__36057;
    wire N__36054;
    wire N__36049;
    wire N__36046;
    wire N__36045;
    wire N__36044;
    wire N__36041;
    wire N__36038;
    wire N__36035;
    wire N__36028;
    wire N__36027;
    wire N__36026;
    wire N__36025;
    wire N__36022;
    wire N__36021;
    wire N__36020;
    wire N__36017;
    wire N__36014;
    wire N__36005;
    wire N__35998;
    wire N__35995;
    wire N__35994;
    wire N__35993;
    wire N__35990;
    wire N__35987;
    wire N__35984;
    wire N__35977;
    wire N__35976;
    wire N__35975;
    wire N__35974;
    wire N__35973;
    wire N__35970;
    wire N__35969;
    wire N__35966;
    wire N__35965;
    wire N__35962;
    wire N__35961;
    wire N__35960;
    wire N__35957;
    wire N__35944;
    wire N__35941;
    wire N__35938;
    wire N__35929;
    wire N__35926;
    wire N__35923;
    wire N__35922;
    wire N__35921;
    wire N__35920;
    wire N__35917;
    wire N__35914;
    wire N__35909;
    wire N__35902;
    wire N__35901;
    wire N__35898;
    wire N__35895;
    wire N__35892;
    wire N__35889;
    wire N__35884;
    wire N__35881;
    wire N__35878;
    wire N__35875;
    wire N__35872;
    wire N__35869;
    wire N__35866;
    wire N__35863;
    wire N__35860;
    wire N__35859;
    wire N__35854;
    wire N__35851;
    wire N__35850;
    wire N__35849;
    wire N__35844;
    wire N__35841;
    wire N__35836;
    wire N__35833;
    wire N__35830;
    wire N__35829;
    wire N__35826;
    wire N__35823;
    wire N__35818;
    wire N__35817;
    wire N__35816;
    wire N__35809;
    wire N__35808;
    wire N__35805;
    wire N__35804;
    wire N__35801;
    wire N__35800;
    wire N__35797;
    wire N__35794;
    wire N__35791;
    wire N__35788;
    wire N__35779;
    wire N__35778;
    wire N__35777;
    wire N__35776;
    wire N__35769;
    wire N__35766;
    wire N__35765;
    wire N__35764;
    wire N__35763;
    wire N__35758;
    wire N__35751;
    wire N__35746;
    wire N__35743;
    wire N__35740;
    wire N__35737;
    wire N__35736;
    wire N__35735;
    wire N__35734;
    wire N__35733;
    wire N__35730;
    wire N__35729;
    wire N__35726;
    wire N__35723;
    wire N__35720;
    wire N__35717;
    wire N__35712;
    wire N__35705;
    wire N__35702;
    wire N__35699;
    wire N__35692;
    wire N__35689;
    wire N__35688;
    wire N__35687;
    wire N__35686;
    wire N__35685;
    wire N__35684;
    wire N__35681;
    wire N__35674;
    wire N__35671;
    wire N__35668;
    wire N__35659;
    wire N__35656;
    wire N__35655;
    wire N__35654;
    wire N__35651;
    wire N__35646;
    wire N__35641;
    wire N__35640;
    wire N__35639;
    wire N__35636;
    wire N__35631;
    wire N__35628;
    wire N__35625;
    wire N__35620;
    wire N__35619;
    wire N__35614;
    wire N__35611;
    wire N__35608;
    wire N__35605;
    wire N__35602;
    wire N__35599;
    wire N__35596;
    wire N__35593;
    wire N__35590;
    wire N__35587;
    wire N__35584;
    wire N__35581;
    wire N__35580;
    wire N__35579;
    wire N__35574;
    wire N__35571;
    wire N__35568;
    wire N__35565;
    wire N__35562;
    wire N__35559;
    wire N__35556;
    wire N__35551;
    wire N__35548;
    wire N__35547;
    wire N__35542;
    wire N__35539;
    wire N__35536;
    wire N__35533;
    wire N__35530;
    wire N__35527;
    wire N__35526;
    wire N__35521;
    wire N__35518;
    wire N__35515;
    wire N__35512;
    wire N__35509;
    wire N__35506;
    wire N__35503;
    wire N__35502;
    wire N__35497;
    wire N__35494;
    wire N__35491;
    wire N__35488;
    wire N__35485;
    wire N__35482;
    wire N__35479;
    wire N__35478;
    wire N__35477;
    wire N__35474;
    wire N__35469;
    wire N__35464;
    wire N__35463;
    wire N__35458;
    wire N__35455;
    wire N__35454;
    wire N__35449;
    wire N__35446;
    wire N__35443;
    wire N__35440;
    wire N__35437;
    wire N__35436;
    wire N__35435;
    wire N__35430;
    wire N__35427;
    wire N__35422;
    wire N__35419;
    wire N__35416;
    wire N__35413;
    wire N__35410;
    wire N__35409;
    wire N__35404;
    wire N__35401;
    wire N__35398;
    wire N__35395;
    wire N__35392;
    wire N__35389;
    wire N__35386;
    wire N__35383;
    wire N__35382;
    wire N__35377;
    wire N__35374;
    wire N__35373;
    wire N__35368;
    wire N__35365;
    wire N__35362;
    wire N__35359;
    wire N__35356;
    wire N__35355;
    wire N__35354;
    wire N__35347;
    wire N__35344;
    wire N__35341;
    wire N__35338;
    wire N__35335;
    wire N__35332;
    wire N__35329;
    wire N__35328;
    wire N__35323;
    wire N__35320;
    wire N__35319;
    wire N__35314;
    wire N__35311;
    wire N__35308;
    wire N__35307;
    wire N__35302;
    wire N__35299;
    wire N__35296;
    wire N__35293;
    wire N__35290;
    wire N__35287;
    wire N__35286;
    wire N__35285;
    wire N__35278;
    wire N__35275;
    wire N__35272;
    wire N__35269;
    wire N__35266;
    wire N__35263;
    wire N__35260;
    wire N__35259;
    wire N__35254;
    wire N__35251;
    wire N__35248;
    wire N__35245;
    wire N__35242;
    wire N__35241;
    wire N__35240;
    wire N__35237;
    wire N__35234;
    wire N__35231;
    wire N__35226;
    wire N__35221;
    wire N__35218;
    wire N__35217;
    wire N__35214;
    wire N__35211;
    wire N__35206;
    wire N__35203;
    wire N__35202;
    wire N__35199;
    wire N__35196;
    wire N__35193;
    wire N__35190;
    wire N__35187;
    wire N__35182;
    wire N__35179;
    wire N__35176;
    wire N__35173;
    wire N__35172;
    wire N__35167;
    wire N__35164;
    wire N__35163;
    wire N__35160;
    wire N__35157;
    wire N__35154;
    wire N__35149;
    wire N__35148;
    wire N__35145;
    wire N__35142;
    wire N__35139;
    wire N__35136;
    wire N__35131;
    wire N__35130;
    wire N__35127;
    wire N__35126;
    wire N__35123;
    wire N__35120;
    wire N__35117;
    wire N__35114;
    wire N__35107;
    wire N__35104;
    wire N__35101;
    wire N__35098;
    wire N__35097;
    wire N__35092;
    wire N__35089;
    wire N__35088;
    wire N__35087;
    wire N__35082;
    wire N__35079;
    wire N__35076;
    wire N__35073;
    wire N__35070;
    wire N__35067;
    wire N__35064;
    wire N__35061;
    wire N__35056;
    wire N__35055;
    wire N__35052;
    wire N__35049;
    wire N__35044;
    wire N__35043;
    wire N__35038;
    wire N__35035;
    wire N__35032;
    wire N__35031;
    wire N__35026;
    wire N__35023;
    wire N__35020;
    wire N__35019;
    wire N__35014;
    wire N__35011;
    wire N__35008;
    wire N__35005;
    wire N__35002;
    wire N__34999;
    wire N__34998;
    wire N__34995;
    wire N__34992;
    wire N__34989;
    wire N__34986;
    wire N__34983;
    wire N__34980;
    wire N__34977;
    wire N__34972;
    wire N__34971;
    wire N__34968;
    wire N__34965;
    wire N__34962;
    wire N__34957;
    wire N__34956;
    wire N__34951;
    wire N__34948;
    wire N__34947;
    wire N__34944;
    wire N__34941;
    wire N__34936;
    wire N__34933;
    wire N__34930;
    wire N__34929;
    wire N__34924;
    wire N__34921;
    wire N__34918;
    wire N__34915;
    wire N__34912;
    wire N__34909;
    wire N__34906;
    wire N__34903;
    wire N__34900;
    wire N__34897;
    wire N__34894;
    wire N__34891;
    wire N__34888;
    wire N__34885;
    wire N__34882;
    wire N__34879;
    wire N__34876;
    wire N__34873;
    wire N__34870;
    wire N__34867;
    wire N__34864;
    wire N__34861;
    wire N__34858;
    wire N__34855;
    wire N__34852;
    wire N__34849;
    wire N__34846;
    wire N__34843;
    wire N__34842;
    wire N__34839;
    wire N__34836;
    wire N__34831;
    wire N__34828;
    wire N__34825;
    wire N__34822;
    wire N__34819;
    wire N__34816;
    wire N__34813;
    wire N__34810;
    wire N__34807;
    wire N__34804;
    wire N__34801;
    wire N__34798;
    wire N__34795;
    wire N__34792;
    wire N__34789;
    wire N__34786;
    wire N__34783;
    wire N__34780;
    wire N__34777;
    wire N__34774;
    wire N__34771;
    wire N__34768;
    wire N__34765;
    wire N__34762;
    wire N__34759;
    wire N__34756;
    wire N__34753;
    wire N__34750;
    wire N__34747;
    wire N__34744;
    wire N__34741;
    wire N__34738;
    wire N__34737;
    wire N__34736;
    wire N__34735;
    wire N__34734;
    wire N__34733;
    wire N__34732;
    wire N__34731;
    wire N__34730;
    wire N__34729;
    wire N__34728;
    wire N__34727;
    wire N__34726;
    wire N__34725;
    wire N__34724;
    wire N__34723;
    wire N__34690;
    wire N__34687;
    wire N__34684;
    wire N__34681;
    wire N__34680;
    wire N__34677;
    wire N__34674;
    wire N__34671;
    wire N__34666;
    wire N__34663;
    wire N__34662;
    wire N__34659;
    wire N__34656;
    wire N__34653;
    wire N__34648;
    wire N__34645;
    wire N__34642;
    wire N__34639;
    wire N__34636;
    wire N__34633;
    wire N__34630;
    wire N__34627;
    wire N__34624;
    wire N__34621;
    wire N__34618;
    wire N__34615;
    wire N__34612;
    wire N__34611;
    wire N__34610;
    wire N__34603;
    wire N__34600;
    wire N__34597;
    wire N__34596;
    wire N__34591;
    wire N__34588;
    wire N__34585;
    wire N__34582;
    wire N__34579;
    wire N__34576;
    wire N__34573;
    wire N__34570;
    wire N__34567;
    wire N__34566;
    wire N__34565;
    wire N__34562;
    wire N__34559;
    wire N__34556;
    wire N__34549;
    wire N__34548;
    wire N__34545;
    wire N__34542;
    wire N__34539;
    wire N__34534;
    wire N__34533;
    wire N__34530;
    wire N__34527;
    wire N__34524;
    wire N__34519;
    wire N__34518;
    wire N__34515;
    wire N__34512;
    wire N__34509;
    wire N__34504;
    wire N__34503;
    wire N__34500;
    wire N__34497;
    wire N__34494;
    wire N__34489;
    wire N__34488;
    wire N__34485;
    wire N__34482;
    wire N__34479;
    wire N__34474;
    wire N__34473;
    wire N__34470;
    wire N__34467;
    wire N__34462;
    wire N__34459;
    wire N__34456;
    wire N__34453;
    wire N__34450;
    wire N__34447;
    wire N__34444;
    wire N__34441;
    wire N__34438;
    wire N__34435;
    wire N__34432;
    wire N__34429;
    wire N__34426;
    wire N__34423;
    wire N__34420;
    wire N__34417;
    wire N__34414;
    wire N__34411;
    wire N__34408;
    wire N__34405;
    wire N__34402;
    wire N__34399;
    wire N__34396;
    wire N__34393;
    wire N__34390;
    wire N__34387;
    wire N__34384;
    wire N__34381;
    wire N__34378;
    wire N__34375;
    wire N__34372;
    wire N__34369;
    wire N__34366;
    wire N__34363;
    wire N__34360;
    wire N__34357;
    wire N__34354;
    wire N__34351;
    wire N__34348;
    wire N__34345;
    wire N__34342;
    wire N__34339;
    wire N__34336;
    wire N__34333;
    wire N__34330;
    wire N__34327;
    wire N__34324;
    wire N__34321;
    wire N__34318;
    wire N__34315;
    wire N__34312;
    wire N__34309;
    wire N__34306;
    wire N__34303;
    wire N__34300;
    wire N__34297;
    wire N__34294;
    wire N__34291;
    wire N__34288;
    wire N__34285;
    wire N__34282;
    wire N__34279;
    wire N__34276;
    wire N__34273;
    wire N__34270;
    wire N__34267;
    wire N__34264;
    wire N__34261;
    wire N__34258;
    wire N__34255;
    wire N__34252;
    wire N__34249;
    wire N__34246;
    wire N__34243;
    wire N__34240;
    wire N__34237;
    wire N__34234;
    wire N__34231;
    wire N__34228;
    wire N__34225;
    wire N__34222;
    wire N__34219;
    wire N__34216;
    wire N__34213;
    wire N__34210;
    wire N__34207;
    wire N__34204;
    wire N__34201;
    wire N__34198;
    wire N__34195;
    wire N__34192;
    wire N__34189;
    wire N__34186;
    wire N__34183;
    wire N__34180;
    wire N__34179;
    wire N__34178;
    wire N__34175;
    wire N__34170;
    wire N__34165;
    wire N__34162;
    wire N__34159;
    wire N__34156;
    wire N__34153;
    wire N__34150;
    wire N__34147;
    wire N__34144;
    wire N__34141;
    wire N__34138;
    wire N__34135;
    wire N__34132;
    wire N__34129;
    wire N__34126;
    wire N__34123;
    wire N__34120;
    wire N__34117;
    wire N__34114;
    wire N__34113;
    wire N__34112;
    wire N__34105;
    wire N__34102;
    wire N__34101;
    wire N__34098;
    wire N__34097;
    wire N__34090;
    wire N__34087;
    wire N__34086;
    wire N__34085;
    wire N__34084;
    wire N__34081;
    wire N__34074;
    wire N__34069;
    wire N__34066;
    wire N__34063;
    wire N__34060;
    wire N__34057;
    wire N__34054;
    wire N__34053;
    wire N__34052;
    wire N__34049;
    wire N__34044;
    wire N__34039;
    wire N__34038;
    wire N__34035;
    wire N__34032;
    wire N__34027;
    wire N__34024;
    wire N__34021;
    wire N__34018;
    wire N__34015;
    wire N__34014;
    wire N__34011;
    wire N__34008;
    wire N__34003;
    wire N__34000;
    wire N__33997;
    wire N__33994;
    wire N__33993;
    wire N__33990;
    wire N__33987;
    wire N__33982;
    wire N__33979;
    wire N__33978;
    wire N__33975;
    wire N__33974;
    wire N__33971;
    wire N__33968;
    wire N__33965;
    wire N__33962;
    wire N__33959;
    wire N__33954;
    wire N__33949;
    wire N__33948;
    wire N__33945;
    wire N__33942;
    wire N__33939;
    wire N__33936;
    wire N__33931;
    wire N__33928;
    wire N__33925;
    wire N__33922;
    wire N__33919;
    wire N__33916;
    wire N__33913;
    wire N__33910;
    wire N__33907;
    wire N__33904;
    wire N__33901;
    wire N__33898;
    wire N__33895;
    wire N__33892;
    wire N__33889;
    wire N__33886;
    wire N__33883;
    wire N__33880;
    wire N__33877;
    wire N__33874;
    wire N__33871;
    wire N__33870;
    wire N__33867;
    wire N__33864;
    wire N__33859;
    wire N__33856;
    wire N__33853;
    wire N__33850;
    wire N__33847;
    wire N__33844;
    wire N__33843;
    wire N__33838;
    wire N__33835;
    wire N__33832;
    wire N__33829;
    wire N__33826;
    wire N__33823;
    wire N__33820;
    wire N__33817;
    wire N__33814;
    wire N__33811;
    wire N__33808;
    wire N__33805;
    wire N__33802;
    wire N__33799;
    wire N__33796;
    wire N__33793;
    wire N__33790;
    wire N__33787;
    wire N__33784;
    wire N__33781;
    wire N__33778;
    wire N__33775;
    wire N__33772;
    wire N__33769;
    wire N__33766;
    wire N__33763;
    wire N__33760;
    wire N__33757;
    wire N__33754;
    wire N__33751;
    wire N__33748;
    wire N__33745;
    wire N__33742;
    wire N__33739;
    wire N__33736;
    wire N__33733;
    wire N__33730;
    wire N__33727;
    wire N__33724;
    wire N__33721;
    wire N__33718;
    wire N__33715;
    wire N__33712;
    wire N__33709;
    wire N__33706;
    wire N__33703;
    wire N__33700;
    wire N__33697;
    wire N__33694;
    wire N__33691;
    wire N__33688;
    wire N__33687;
    wire N__33682;
    wire N__33679;
    wire N__33676;
    wire N__33673;
    wire N__33670;
    wire N__33667;
    wire N__33664;
    wire N__33661;
    wire N__33660;
    wire N__33655;
    wire N__33652;
    wire N__33649;
    wire N__33646;
    wire N__33643;
    wire N__33640;
    wire N__33637;
    wire N__33634;
    wire N__33631;
    wire N__33628;
    wire N__33627;
    wire N__33626;
    wire N__33623;
    wire N__33618;
    wire N__33613;
    wire N__33610;
    wire N__33607;
    wire N__33606;
    wire N__33601;
    wire N__33598;
    wire N__33595;
    wire N__33592;
    wire N__33589;
    wire N__33586;
    wire N__33585;
    wire N__33580;
    wire N__33577;
    wire N__33574;
    wire N__33571;
    wire N__33568;
    wire N__33565;
    wire N__33562;
    wire N__33559;
    wire N__33556;
    wire N__33553;
    wire N__33550;
    wire N__33547;
    wire N__33544;
    wire N__33541;
    wire N__33538;
    wire N__33535;
    wire N__33532;
    wire N__33529;
    wire N__33526;
    wire N__33523;
    wire N__33520;
    wire N__33517;
    wire N__33514;
    wire N__33511;
    wire N__33508;
    wire N__33507;
    wire N__33504;
    wire N__33501;
    wire N__33496;
    wire N__33493;
    wire N__33490;
    wire N__33487;
    wire N__33484;
    wire N__33483;
    wire N__33478;
    wire N__33475;
    wire N__33472;
    wire N__33469;
    wire N__33466;
    wire N__33465;
    wire N__33460;
    wire N__33457;
    wire N__33454;
    wire N__33451;
    wire N__33448;
    wire N__33445;
    wire N__33442;
    wire N__33439;
    wire N__33436;
    wire N__33435;
    wire N__33430;
    wire N__33427;
    wire N__33424;
    wire N__33421;
    wire N__33420;
    wire N__33419;
    wire N__33414;
    wire N__33411;
    wire N__33408;
    wire N__33403;
    wire N__33400;
    wire N__33399;
    wire N__33394;
    wire N__33391;
    wire N__33390;
    wire N__33389;
    wire N__33382;
    wire N__33379;
    wire N__33376;
    wire N__33373;
    wire N__33370;
    wire N__33367;
    wire N__33364;
    wire N__33361;
    wire N__33358;
    wire N__33355;
    wire N__33354;
    wire N__33353;
    wire N__33346;
    wire N__33343;
    wire N__33340;
    wire N__33337;
    wire N__33334;
    wire N__33331;
    wire N__33328;
    wire N__33325;
    wire N__33322;
    wire N__33319;
    wire N__33316;
    wire N__33313;
    wire N__33310;
    wire N__33307;
    wire N__33304;
    wire N__33301;
    wire N__33298;
    wire N__33295;
    wire N__33292;
    wire N__33289;
    wire N__33286;
    wire N__33283;
    wire N__33280;
    wire N__33277;
    wire N__33274;
    wire N__33271;
    wire N__33268;
    wire N__33265;
    wire N__33262;
    wire N__33259;
    wire N__33256;
    wire N__33253;
    wire N__33250;
    wire N__33247;
    wire N__33244;
    wire N__33241;
    wire N__33238;
    wire N__33235;
    wire N__33232;
    wire N__33229;
    wire N__33226;
    wire N__33223;
    wire N__33220;
    wire N__33217;
    wire N__33214;
    wire N__33211;
    wire N__33208;
    wire N__33205;
    wire N__33202;
    wire N__33199;
    wire N__33196;
    wire N__33193;
    wire N__33190;
    wire N__33187;
    wire N__33184;
    wire N__33181;
    wire N__33178;
    wire N__33175;
    wire N__33172;
    wire N__33169;
    wire N__33166;
    wire N__33163;
    wire N__33160;
    wire N__33157;
    wire N__33154;
    wire N__33151;
    wire N__33148;
    wire N__33145;
    wire N__33142;
    wire N__33139;
    wire N__33136;
    wire N__33133;
    wire N__33130;
    wire N__33127;
    wire N__33124;
    wire N__33121;
    wire N__33118;
    wire N__33115;
    wire N__33112;
    wire N__33109;
    wire N__33106;
    wire N__33103;
    wire N__33100;
    wire N__33097;
    wire N__33094;
    wire N__33091;
    wire N__33088;
    wire N__33085;
    wire N__33082;
    wire N__33079;
    wire N__33076;
    wire N__33073;
    wire N__33070;
    wire N__33067;
    wire N__33064;
    wire N__33061;
    wire N__33058;
    wire N__33055;
    wire N__33052;
    wire N__33049;
    wire N__33046;
    wire N__33043;
    wire N__33040;
    wire N__33037;
    wire N__33034;
    wire N__33031;
    wire N__33028;
    wire N__33025;
    wire N__33022;
    wire N__33019;
    wire N__33016;
    wire N__33013;
    wire N__33010;
    wire N__33007;
    wire N__33004;
    wire N__33001;
    wire N__32998;
    wire N__32995;
    wire N__32992;
    wire N__32989;
    wire N__32986;
    wire N__32983;
    wire N__32980;
    wire N__32977;
    wire N__32974;
    wire N__32971;
    wire N__32968;
    wire N__32965;
    wire N__32962;
    wire N__32959;
    wire \Pc2drone_pll_inst.clk_system_pll ;
    wire GNDG0;
    wire VCCG0;
    wire \pid_alt.O_3_12 ;
    wire \pid_alt.O_3_14 ;
    wire \pid_alt.O_3_8 ;
    wire \pid_alt.O_3_18 ;
    wire \pid_alt.O_3_22 ;
    wire \pid_alt.O_3_20 ;
    wire \pid_alt.O_3_19 ;
    wire \pid_alt.O_3_21 ;
    wire \pid_alt.O_3_17 ;
    wire \pid_alt.O_3_24 ;
    wire \pid_alt.O_3_7 ;
    wire \pid_alt.O_3_15 ;
    wire \pid_alt.O_3_9 ;
    wire \pid_alt.O_3_10 ;
    wire \pid_alt.O_3_11 ;
    wire \pid_alt.O_3_13 ;
    wire \pid_alt.O_3_16 ;
    wire \pid_alt.O_4_13 ;
    wire \pid_alt.O_4_18 ;
    wire \pid_alt.O_4_19 ;
    wire \pid_alt.O_4_20 ;
    wire \pid_alt.O_4_16 ;
    wire \pid_alt.O_4_17 ;
    wire \pid_alt.O_4_23 ;
    wire \pid_alt.O_4_22 ;
    wire \pid_alt.O_4_24 ;
    wire \pid_alt.O_4_7 ;
    wire \pid_alt.O_4_15 ;
    wire \pid_alt.O_4_10 ;
    wire \pid_alt.O_4_11 ;
    wire \pid_alt.O_4_21 ;
    wire \pid_alt.O_3_4 ;
    wire \pid_alt.O_5_5 ;
    wire \pid_alt.O_4_6 ;
    wire \pid_alt.O_5_6 ;
    wire \pid_alt.O_3_6 ;
    wire \pid_alt.O_5_8 ;
    wire \pid_alt.error_p_reg_esr_RNIOI4PZ0Z_0_cascade_ ;
    wire \pid_alt.error_d_regZ0Z_0 ;
    wire \pid_front.O_0_23 ;
    wire \pid_alt.O_4_5 ;
    wire \pid_alt.O_4_8 ;
    wire \pid_alt.O_4_9 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIGDHM_0Z0Z_11_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNIDAHMZ0Z_10 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIGDHM_0Z0Z_11 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIDAHMZ0Z_10_cascade_ ;
    wire \pid_alt.error_d_reg_prevZ0Z_10 ;
    wire \pid_alt.error_d_regZ0Z_10 ;
    wire \pid_alt.error_d_reg_prevZ0Z_11 ;
    wire \pid_alt.error_d_regZ0Z_11 ;
    wire \pid_alt.O_5_24 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIL8611Z0Z_9_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNIL8611Z0Z_9 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIDAHM_0Z0Z_10 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI20IM_0Z0Z_17 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI20IM_0Z0Z_17_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNIVSHMZ0Z_16 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16_cascade_ ;
    wire \pid_alt.error_d_regZ0Z_16 ;
    wire \pid_alt.error_d_reg_prevZ0Z_16 ;
    wire \pid_alt.O_5_4 ;
    wire \pid_alt.error_p_regZ0Z_0 ;
    wire \pid_alt.O_5_10 ;
    wire \pid_alt.O_5_22 ;
    wire \pid_alt.O_5_23 ;
    wire \pid_alt.O_5_17 ;
    wire \pid_alt.O_5_9 ;
    wire \pid_alt.O_5_21 ;
    wire \pid_alt.error_p_regZ0Z_17 ;
    wire \pid_alt.O_5_11 ;
    wire \pid_alt.O_5_12 ;
    wire \pid_alt.O_5_13 ;
    wire \pid_alt.O_5_7 ;
    wire \pid_alt.O_5_15 ;
    wire \pid_alt.error_p_regZ0Z_11 ;
    wire \pid_alt.O_5_16 ;
    wire \pid_alt.O_5_14 ;
    wire \pid_alt.error_p_regZ0Z_10 ;
    wire \pid_alt.O_5_18 ;
    wire \pid_alt.O_5_19 ;
    wire \pid_alt.O_5_20 ;
    wire \pid_alt.error_p_regZ0Z_16 ;
    wire \pid_alt.O_3_5 ;
    wire alt_kd_0;
    wire alt_kd_1;
    wire alt_kd_2;
    wire alt_kd_3;
    wire alt_kd_4;
    wire alt_kd_5;
    wire alt_kd_6;
    wire alt_kd_7;
    wire \pid_alt.O_4_12 ;
    wire \pid_alt.O_4_14 ;
    wire \pid_alt.O_4_4 ;
    wire alt_ki_5;
    wire alt_ki_6;
    wire \pid_alt.error_p_regZ0Z_2 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI0J511_0Z0Z_2_cascade_ ;
    wire \pid_alt.error_p_regZ0Z_1 ;
    wire \pid_alt.error_d_reg_prevZ0Z_1 ;
    wire \pid_alt.error_d_regZ0Z_1 ;
    wire \pid_alt.un1_pid_prereg_16_0 ;
    wire \pid_alt.error_d_reg_prev_esr_RNITF511_0Z0Z_1_cascade_ ;
    wire \pid_alt.error_d_regZ0Z_2 ;
    wire \pid_alt.error_d_reg_prevZ0Z_2 ;
    wire \pid_alt.error_d_reg_prevZ0Z_0 ;
    wire \pid_alt.error_d_reg_prev_esr_RNITF511Z0Z_1 ;
    wire \pid_alt.error_p_reg_esr_RNIOI4PZ0Z_0 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI0J511_0Z0Z_2 ;
    wire \pid_alt.error_d_reg_prev_esr_RNITF511_0Z0Z_1 ;
    wire \pid_alt.error_d_regZ0Z_17 ;
    wire \pid_alt.error_d_reg_prevZ0Z_17 ;
    wire bfn_2_16_0_;
    wire \pid_alt.error_i_regZ0Z_1 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_0 ;
    wire \pid_alt.error_i_regZ0Z_2 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_1 ;
    wire \pid_alt.error_i_regZ0Z_3 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_2 ;
    wire \pid_alt.error_i_regZ0Z_4 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_3 ;
    wire \pid_alt.error_i_regZ0Z_5 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_4 ;
    wire \pid_alt.error_i_regZ0Z_6 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_5 ;
    wire \pid_alt.error_i_regZ0Z_7 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_6 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_7 ;
    wire \pid_alt.error_i_regZ0Z_8 ;
    wire bfn_2_17_0_;
    wire \pid_alt.error_i_regZ0Z_9 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_8 ;
    wire \pid_alt.error_i_regZ0Z_10 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_9 ;
    wire \pid_alt.error_i_regZ0Z_11 ;
    wire \pid_alt.error_i_reg_esr_RNI4NMPZ0Z_11 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_10 ;
    wire \pid_alt.error_i_regZ0Z_12 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_11 ;
    wire \pid_alt.error_i_regZ0Z_13 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_12 ;
    wire \pid_alt.error_i_regZ0Z_14 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_13 ;
    wire \pid_alt.error_i_regZ0Z_15 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_14 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_15 ;
    wire \pid_alt.error_i_regZ0Z_16 ;
    wire bfn_2_18_0_;
    wire \pid_alt.error_i_regZ0Z_17 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_16 ;
    wire \pid_alt.error_i_regZ0Z_18 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_17 ;
    wire \pid_alt.error_i_regZ0Z_19 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_18 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_19 ;
    wire \pid_alt.error_i_regZ0Z_20 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_20 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16 ;
    wire \pid_alt.error_i_reg_esr_RNI5BMJZ0Z_16 ;
    wire \pid_alt.error_i_acummZ0Z_10 ;
    wire \pid_alt.error_i_acummZ0Z_11 ;
    wire \pid_alt.error_i_acummZ0Z_6 ;
    wire \pid_alt.error_i_acummZ0Z_7 ;
    wire \pid_alt.error_i_acummZ0Z_8 ;
    wire \pid_alt.error_i_acummZ0Z_9 ;
    wire \pid_alt.error_i_acummZ0Z_12 ;
    wire \pid_alt.error_i_acummZ0Z_5 ;
    wire \pid_alt.error_i_acummZ0Z_3 ;
    wire \pid_alt.error_i_acummZ0Z_1 ;
    wire \pid_alt.error_i_acummZ0Z_2 ;
    wire \pid_alt.error_i_acumm_prereg_esr_RNICB6L2_0Z0Z_5_cascade_ ;
    wire \pid_alt.error_i_acumm_prereg_esr_RNICB6L2Z0Z_5 ;
    wire \pid_alt.N_159 ;
    wire \pid_alt.N_159_cascade_ ;
    wire \pid_alt.error_i_acummZ0Z_4 ;
    wire alt_kp_6;
    wire alt_kp_1;
    wire alt_kp_3;
    wire \pid_front.O_0_9 ;
    wire \pid_alt.O_3_23 ;
    wire \pid_alt.N_933_0_g ;
    wire alt_ki_0;
    wire alt_ki_1;
    wire alt_ki_2;
    wire alt_ki_3;
    wire alt_ki_4;
    wire alt_ki_7;
    wire \pid_alt.error_p_regZ0Z_3 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI3M511Z0Z_3 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI3M511Z0Z_3_cascade_ ;
    wire \pid_alt.error_p_regZ0Z_4 ;
    wire \pid_alt.error_d_reg_prevZ0Z_4 ;
    wire \pid_alt.error_d_regZ0Z_4 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI6P511_0Z0Z_4 ;
    wire \pid_alt.error_d_regZ0Z_3 ;
    wire \pid_alt.error_d_reg_prevZ0Z_3 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI3M511_0Z0Z_3 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI0J511Z0Z_2 ;
    wire \pid_alt.error_d_reg_prev_esr_RNII5LS3Z0Z_1 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI9S511Z0Z_5 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI9S511Z0Z_5_cascade_ ;
    wire \pid_alt.error_p_regZ0Z_6 ;
    wire \pid_alt.error_d_reg_prevZ0Z_6 ;
    wire \pid_alt.error_d_regZ0Z_6 ;
    wire \pid_alt.error_d_reg_prev_esr_RNICV511_0Z0Z_6 ;
    wire \pid_alt.error_d_reg_prevZ0Z_5 ;
    wire \pid_alt.error_p_regZ0Z_5 ;
    wire \pid_alt.error_d_regZ0Z_5 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI9S511_0Z0Z_5 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI6P511Z0Z_4 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI9S511_0Z0Z_5_cascade_ ;
    wire \pid_alt.error_d_regZ0Z_13 ;
    wire \pid_alt.error_d_reg_prevZ0Z_13 ;
    wire \pid_alt.error_p_regZ0Z_13 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIMJHM_0Z0Z_13 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIMJHM_0Z0Z_13_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12 ;
    wire \pid_alt.error_d_reg_prevZ0Z_12 ;
    wire \pid_alt.error_p_regZ0Z_12 ;
    wire \pid_alt.error_d_regZ0Z_12 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIGDHMZ0Z_11 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNISPHM_0Z0Z_15 ;
    wire \pid_alt.error_d_reg_prev_esr_RNISPHM_0Z0Z_15_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNIPMHMZ0Z_14 ;
    wire \pid_alt.error_p_regZ0Z_14 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14_cascade_ ;
    wire \pid_alt.error_d_regZ0Z_14 ;
    wire \pid_alt.error_d_reg_prevZ0Z_14 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIMJHMZ0Z_13 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNI86IM_0Z0Z_19 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI86IM_0Z0Z_19_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18 ;
    wire \pid_alt.error_d_regZ0Z_18 ;
    wire \pid_alt.error_p_regZ0Z_18 ;
    wire \pid_alt.error_d_reg_prevZ0Z_18 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI20IMZ0Z_17 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18_cascade_ ;
    wire \pid_alt.error_i_reg_esr_RNI9HOJZ0Z_18 ;
    wire \pid_alt.error_p_regZ0Z_19 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI86IMZ0Z_19_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNI86IMZ0Z_19 ;
    wire \pid_alt.un1_pid_prereg_236_1 ;
    wire \pid_alt.error_d_regZ0Z_19 ;
    wire \pid_alt.error_d_reg_prevZ0Z_19 ;
    wire \pid_alt.error_d_reg_prevZ0Z_20 ;
    wire \pid_alt.error_d_regZ0Z_20 ;
    wire \pid_alt.error_p_regZ0Z_20 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_20_c_RNISVKK ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_9_c_RNIQN3F ;
    wire \pid_alt.error_i_reg_esr_RNI7RNPZ0Z_12 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_10 ;
    wire \pid_alt.m21_e_2_cascade_ ;
    wire \pid_alt.error_i_acumm_preregZ0Z_2 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_3 ;
    wire \pid_alt.m35_e_3 ;
    wire \pid_alt.N_62_mux ;
    wire \pid_alt.N_545_cascade_ ;
    wire \pid_alt.error_i_acumm7lto12 ;
    wire \pid_alt.N_158 ;
    wire \pid_alt.error_i_acumm_prereg_esr_RNIFJA3Z0Z_14_cascade_ ;
    wire \pid_alt.N_9_0 ;
    wire \pid_alt.N_9_0_cascade_ ;
    wire \pid_alt.m21_e_10 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_18 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_16 ;
    wire \pid_alt.m7_e_4 ;
    wire \pid_alt.error_i_acumm_esr_RNI33H91Z0Z_4 ;
    wire \pid_alt.error_i_reg_esr_RNI7ENJZ0Z_17 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_17 ;
    wire \pid_alt.error_i_reg_esr_RNI38LJZ0Z_15 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_15 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ ;
    wire \pid_alt.error_i_acumm_preregZ0Z_20 ;
    wire \pid_alt.error_i_acumm_esr_RNIJ6LMZ0Z_13 ;
    wire alt_kp_5;
    wire alt_kp_7;
    wire alt_kp_0;
    wire \ppm_encoder_1.pulses2count_9_i_3_1_2_cascade_ ;
    wire \ppm_encoder_1.pulses2count_9_0_0_1 ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_5 ;
    wire \ppm_encoder_1.N_513_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_2 ;
    wire \ppm_encoder_1.un2_throttle_0_0_2_5_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_0_0_5 ;
    wire \ppm_encoder_1.pulses2count_9_0_1_1 ;
    wire \ppm_encoder_1.rudderZ0Z_5 ;
    wire \ppm_encoder_1.N_507_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_0_1_2_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_2_cascade_ ;
    wire \ppm_encoder_1.N_264_i_i_cascade_ ;
    wire \ppm_encoder_1.N_465_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_0_2_8_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_8 ;
    wire \ppm_encoder_1.throttleZ0Z_2 ;
    wire \ppm_encoder_1.aileronZ0Z_5 ;
    wire \ppm_encoder_1.throttleZ0Z_1 ;
    wire \ppm_encoder_1.throttleZ0Z_5 ;
    wire bfn_4_9_0_;
    wire \ppm_encoder_1.un1_throttle_cry_0_THRU_CO ;
    wire \ppm_encoder_1.un1_throttle_cry_0 ;
    wire \ppm_encoder_1.un1_throttle_cry_1_THRU_CO ;
    wire \ppm_encoder_1.un1_throttle_cry_1 ;
    wire \ppm_encoder_1.un1_throttle_cry_2_THRU_CO ;
    wire \ppm_encoder_1.un1_throttle_cry_2 ;
    wire \ppm_encoder_1.un1_throttle_cry_3_THRU_CO ;
    wire \ppm_encoder_1.un1_throttle_cry_3 ;
    wire \ppm_encoder_1.un1_throttle_cry_4_THRU_CO ;
    wire \ppm_encoder_1.un1_throttle_cry_4 ;
    wire \ppm_encoder_1.un1_throttle_cry_5_THRU_CO ;
    wire \ppm_encoder_1.un1_throttle_cry_5 ;
    wire \ppm_encoder_1.un1_throttle_cry_6 ;
    wire \ppm_encoder_1.un1_throttle_cry_7 ;
    wire bfn_4_10_0_;
    wire \ppm_encoder_1.un1_throttle_cry_8 ;
    wire \ppm_encoder_1.un1_throttle_cry_9_THRU_CO ;
    wire \ppm_encoder_1.un1_throttle_cry_9 ;
    wire \ppm_encoder_1.un1_throttle_cry_10_THRU_CO ;
    wire \ppm_encoder_1.un1_throttle_cry_10 ;
    wire \ppm_encoder_1.un1_throttle_cry_11 ;
    wire \ppm_encoder_1.un1_throttle_cry_12_THRU_CO ;
    wire \ppm_encoder_1.un1_throttle_cry_12 ;
    wire \ppm_encoder_1.un1_throttle_cry_13 ;
    wire throttle_order_10;
    wire \pid_alt.source_pid_1_sqmuxa_0_a2_1_4_cascade_ ;
    wire throttle_order_11;
    wire throttle_order_6;
    wire \pid_alt.source_pid_9_0_tz_6 ;
    wire \pid_alt.N_52_cascade_ ;
    wire \pid_alt.N_54_cascade_ ;
    wire throttle_order_1;
    wire throttle_order_2;
    wire \pid_alt.N_54 ;
    wire throttle_order_3;
    wire \pid_alt.error_d_reg_prev_i_0 ;
    wire bfn_4_13_0_;
    wire \pid_alt.error_p_reg_esr_RNI3SMI1Z0Z_0 ;
    wire \pid_alt.un1_pid_prereg_0 ;
    wire \pid_alt.pid_preregZ0Z_0 ;
    wire \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CO ;
    wire \pid_alt.error_d_reg_prev_esr_RNIFPN33Z0Z_1 ;
    wire \pid_alt.pid_preregZ0Z_1 ;
    wire \pid_alt.un1_pid_prereg_0_cry_0 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIF0465Z0Z_1 ;
    wire \pid_alt.error_i_acumm_esr_RNITQE91Z0Z_2 ;
    wire \pid_alt.pid_preregZ0Z_2 ;
    wire \pid_alt.un1_pid_prereg_0_cry_1 ;
    wire \pid_alt.error_d_reg_prev_esr_RNILDG87Z0Z_2 ;
    wire \pid_alt.error_i_acumm_esr_RNI0VF91Z0Z_3 ;
    wire \pid_alt.pid_preregZ0Z_3 ;
    wire \pid_alt.un1_pid_prereg_0_cry_2 ;
    wire \pid_alt.error_d_reg_prev_esr_RNILE0V5Z0Z_2 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI11TA9Z0Z_3 ;
    wire \pid_alt.un1_pid_prereg_0_cry_3 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIOGSO6Z0Z_4 ;
    wire \pid_alt.error_d_reg_prev_esr_RNICISB3Z0Z_3 ;
    wire \pid_alt.un1_pid_prereg_0_cry_4 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI171A6Z0Z_5 ;
    wire \pid_alt.error_d_reg_prev_esr_RNICUVC3Z0Z_4 ;
    wire \pid_alt.un1_pid_prereg_0_cry_5 ;
    wire \pid_alt.un1_pid_prereg_0_cry_6 ;
    wire bfn_4_14_0_;
    wire \pid_alt.un1_pid_prereg_0_cry_7 ;
    wire \pid_alt.un1_pid_prereg_0_cry_8 ;
    wire \pid_alt.error_d_reg_prev_esr_RNICI045Z0Z_9 ;
    wire \pid_alt.un1_pid_prereg_0_cry_9 ;
    wire \pid_alt.error_d_reg_prev_esr_RNITPKD4Z0Z_10 ;
    wire \pid_alt.error_d_reg_prev_esr_RNISAR62Z0Z_9 ;
    wire \pid_alt.un1_pid_prereg_0_cry_10 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIB8KD4Z0Z_11 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI1FP62Z0Z_10 ;
    wire \pid_alt.un1_pid_prereg_0_cry_11 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI64JA4Z0Z_12 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIAPQ62Z0Z_11 ;
    wire \pid_alt.un1_pid_prereg_0_cry_12 ;
    wire \pid_alt.error_d_reg_prev_esr_RNICQF44Z0Z_13 ;
    wire \pid_alt.error_d_reg_prev_esr_RNISAO32Z0Z_12 ;
    wire \pid_alt.un1_pid_prereg_0_cry_13 ;
    wire \pid_alt.un1_pid_prereg_0_cry_14 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI88G14Z0Z_14 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIGFN02Z0Z_13 ;
    wire bfn_4_15_0_;
    wire \pid_alt.error_d_reg_prev_esr_RNIOQI14Z0Z_15 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIOOO02Z0Z_14 ;
    wire \pid_alt.un1_pid_prereg_0_cry_15 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI02Q02Z0Z_15 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI8DL14Z0Z_16 ;
    wire \pid_alt.un1_pid_prereg_0_cry_16 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIOVN14Z0Z_17 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI8BR02Z0Z_16 ;
    wire \pid_alt.un1_pid_prereg_0_cry_17 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI8IQ14Z0Z_18 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIGKS02Z0Z_17 ;
    wire \pid_alt.un1_pid_prereg_0_cry_18 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIK3024Z0Z_19 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIOTT02Z0Z_18 ;
    wire \pid_alt.un1_pid_prereg_0_cry_19 ;
    wire \pid_alt.error_d_reg_prev_esr_RNICG9B1_0Z0Z_20 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIS5212Z0Z_19 ;
    wire \pid_alt.un1_pid_prereg_0_cry_20 ;
    wire \pid_alt.error_d_reg_prev_esr_RNICG9B1_1Z0Z_20 ;
    wire \pid_alt.un1_pid_prereg_0_cry_21 ;
    wire \pid_alt.un1_pid_prereg_0_cry_22 ;
    wire \pid_alt.error_d_reg_prev_esr_RNICG9B1Z0Z_20 ;
    wire \pid_alt.error_d_reg_prev_esr_RNICG9B1_2Z0Z_20 ;
    wire bfn_4_16_0_;
    wire \pid_alt.un1_pid_prereg_0_axb_24 ;
    wire \pid_alt.un1_pid_prereg_0_cry_23 ;
    wire \pid_alt.error_i_reg_esr_RNI15KJZ0Z_14 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_14 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ ;
    wire \pid_alt.error_i_reg_esr_RNIBKPJZ0Z_19 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_19 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIN49Q5Z0Z_8 ;
    wire \pid_alt.error_p_regZ0Z_9 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNIG75T2Z0Z_8 ;
    wire \pid_alt.error_d_reg_prev_esr_RNII5611Z0Z_8 ;
    wire \pid_alt.error_d_regZ0Z_9 ;
    wire \pid_alt.error_d_reg_prevZ0Z_9 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_8_c_RNI9POQ ;
    wire \pid_alt.error_i_acumm_preregZ0Z_9 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_8 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_11 ;
    wire \pid_alt.m21_e_8 ;
    wire bfn_4_18_0_;
    wire \pid_alt.error_1 ;
    wire \pid_alt.error_cry_0 ;
    wire \pid_alt.error_2 ;
    wire \pid_alt.error_cry_1 ;
    wire \pid_alt.error_3 ;
    wire \pid_alt.error_cry_2 ;
    wire \pid_alt.error_4 ;
    wire \pid_alt.error_cry_3 ;
    wire \pid_alt.error_5 ;
    wire \pid_alt.error_cry_4 ;
    wire \pid_alt.error_6 ;
    wire \pid_alt.error_cry_5 ;
    wire \pid_alt.error_7 ;
    wire \pid_alt.error_cry_6 ;
    wire \pid_alt.error_cry_7 ;
    wire \pid_alt.error_8 ;
    wire bfn_4_19_0_;
    wire \pid_alt.error_9 ;
    wire \pid_alt.error_cry_8 ;
    wire \pid_alt.error_10 ;
    wire \pid_alt.error_cry_9 ;
    wire \pid_alt.error_11 ;
    wire \pid_alt.error_cry_10 ;
    wire \pid_alt.error_12 ;
    wire \pid_alt.error_cry_11 ;
    wire \pid_alt.error_13 ;
    wire \pid_alt.error_cry_12 ;
    wire \pid_alt.error_14 ;
    wire \pid_alt.error_cry_13 ;
    wire \pid_alt.error_cry_14 ;
    wire \pid_alt.error_15 ;
    wire \pid_alt.error_i_acumm_esr_RNIQMD91Z0Z_1 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_1 ;
    wire \pid_alt.m21_e_0_cascade_ ;
    wire \pid_alt.error_i_acumm7lto4 ;
    wire \pid_alt.m21_e_9 ;
    wire \pid_alt.error_i_regZ0Z_0 ;
    wire \pid_alt.error_i_acummZ0Z_0 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_0 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_7 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_6 ;
    wire \pid_alt.m35_e_2 ;
    wire \pid_alt.error_i_reg_esr_RNIT8KA1Z0Z_5 ;
    wire \pid_alt.error_i_acumm7lto5 ;
    wire \pid_front.O_0_20 ;
    wire \ppm_encoder_1.PPM_STATE_fastZ0Z_0 ;
    wire \ppm_encoder_1.PPM_STATE_fast_RNICIABZ0Z_0_cascade_ ;
    wire \ppm_encoder_1.aileron_RNI7E8E1Z0Z_1_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_0_1_1_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_0_0_1 ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_1_cascade_ ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI6LFQZ0Z_0_cascade_ ;
    wire \ppm_encoder_1.N_303_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_0_2_2 ;
    wire \ppm_encoder_1.N_448_cascade_ ;
    wire \ppm_encoder_1.elevatorZ0Z_12 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_2_3_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_0_1_3 ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_3_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_0_1_8 ;
    wire \ppm_encoder_1.throttleZ0Z_4 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_1_4 ;
    wire \ppm_encoder_1.N_260_i_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_4_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_0_2_9_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_9_cascade_ ;
    wire \ppm_encoder_1.N_454 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_1_9 ;
    wire \ppm_encoder_1.throttleZ0Z_13 ;
    wire \pid_alt.source_pid_1_sqmuxa_0_a2_0_3_cascade_ ;
    wire \pid_alt.N_57_cascade_ ;
    wire \pid_alt.un1_reset_1_cascade_ ;
    wire \pid_alt.un1_reset_0_i_cascade_ ;
    wire \pid_alt.pid_preregZ0Z_8 ;
    wire \pid_alt.pid_preregZ0Z_7 ;
    wire \pid_alt.pid_preregZ0Z_9 ;
    wire \pid_alt.pid_preregZ0Z_6 ;
    wire \pid_alt.pid_preregZ0Z_11 ;
    wire \pid_alt.source_pid_1_sqmuxa_0_o2_3_cascade_ ;
    wire \pid_alt.pid_preregZ0Z_10 ;
    wire \pid_alt.N_51 ;
    wire \pid_alt.source_pid_1_sqmuxa_0_a2_0_2 ;
    wire \pid_alt.source_pid_1_sqmuxa_0_a2_1_5 ;
    wire \pid_alt.source_pid_1_sqmuxa_0_a2_1_7 ;
    wire \pid_alt.pid_preregZ0Z_22 ;
    wire \pid_alt.pid_preregZ0Z_19 ;
    wire \pid_alt.pid_preregZ0Z_20 ;
    wire \pid_alt.pid_preregZ0Z_17 ;
    wire \pid_alt.pid_preregZ0Z_23 ;
    wire \pid_alt.pid_preregZ0Z_18 ;
    wire \pid_alt.pid_preregZ0Z_21 ;
    wire \pid_alt.pid_preregZ0Z_15 ;
    wire \pid_alt.pid_preregZ0Z_16 ;
    wire \pid_alt.pid_preregZ0Z_14 ;
    wire \pid_alt.source_pid_1_sqmuxa_0_a2_2_5_cascade_ ;
    wire \pid_alt.source_pid_1_sqmuxa_0_a2_2_6 ;
    wire \pid_alt.N_539_cascade_ ;
    wire \pid_alt.pid_preregZ0Z_4 ;
    wire \pid_alt.source_pid_9_0_0_4_cascade_ ;
    wire throttle_order_4;
    wire \pid_alt.N_52 ;
    wire throttle_order_5;
    wire \pid_alt.pid_preregZ0Z_24 ;
    wire \pid_alt.pid_preregZ0Z_13 ;
    wire \pid_alt.N_539 ;
    wire throttle_order_13;
    wire \pid_alt.N_72_i_1 ;
    wire \pid_alt.un1_reset_0_i ;
    wire \pid_alt.error_d_reg_prev_esr_RNI5G6Q5Z0Z_7 ;
    wire \pid_alt.error_p_regZ0Z_8 ;
    wire \pid_alt.error_d_reg_prevZ0Z_8 ;
    wire \pid_alt.error_d_regZ0Z_8 ;
    wire \pid_alt.error_d_reg_prev_esr_RNII5611_0Z0Z_8 ;
    wire \pid_alt.error_d_reg_prev_esr_RNII5611_0Z0Z_8_cascade_ ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ ;
    wire \pid_alt.error_d_reg_prev_esr_RNI7T3T2Z0Z_7 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIF2611Z0Z_7 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIUI2T2Z0Z_6 ;
    wire \pid_alt.error_d_regZ0Z_7 ;
    wire \pid_alt.error_d_reg_prevZ0Z_7 ;
    wire \pid_alt.error_p_regZ0Z_7 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIF2611_0Z0Z_7 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIL81T2Z0Z_5 ;
    wire \pid_alt.error_d_reg_prev_esr_RNICV511Z0Z_6 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIF2611_0Z0Z_7_cascade_ ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ ;
    wire \pid_alt.error_d_reg_prev_esr_RNIJR3Q5Z0Z_6 ;
    wire \pid_front.O_0_21 ;
    wire \pid_front.O_0_7 ;
    wire \pid_front.O_0_11 ;
    wire \pid_front.O_0_12 ;
    wire uart_input_pc_c;
    wire \uart_pc_sync.aux_0__0_Z0Z_0 ;
    wire \pid_alt.pid_preregZ0Z_12 ;
    wire \pid_alt.pid_preregZ0Z_5 ;
    wire \pid_alt.N_154 ;
    wire \pid_alt.state_1_0_0 ;
    wire \Commands_frame_decoder.source_CH1data8_cascade_ ;
    wire alt_command_1;
    wire \Commands_frame_decoder.source_CH1data8lto7Z0Z_2 ;
    wire alt_command_3;
    wire alt_command_0;
    wire \Commands_frame_decoder.source_CH1data8 ;
    wire alt_command_2;
    wire \Commands_frame_decoder.state_ns_i_a2_0_2_0_cascade_ ;
    wire alt_command_4;
    wire alt_command_5;
    wire alt_command_6;
    wire alt_kp_2;
    wire drone_altitude_i_8;
    wire \pid_alt.error_p_regZ0Z_15 ;
    wire \pid_alt.error_d_reg_prev_esr_RNISPHMZ0Z_15 ;
    wire \pid_alt.error_d_regZ0Z_15 ;
    wire \pid_alt.error_d_reg_prevZ0Z_15 ;
    wire \pid_alt.state_0_g_0 ;
    wire \pid_alt.N_111 ;
    wire \pid_alt.un1_reset_1_0_i_cascade_ ;
    wire alt_command_7;
    wire \ppm_encoder_1.init_pulsesZ0Z_1 ;
    wire uart_input_drone_c;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_13 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_0_13_cascade_ ;
    wire \ppm_encoder_1.N_516 ;
    wire \ppm_encoder_1.N_440 ;
    wire \ppm_encoder_1.N_516_cascade_ ;
    wire \uart_drone_sync.aux_0__0__0_0 ;
    wire \ppm_encoder_1.throttleZ0Z_11 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_1_11 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_0_11_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_0_0_4 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_2_10_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_10_cascade_ ;
    wire \ppm_encoder_1.N_458 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_1_10 ;
    wire \ppm_encoder_1.elevatorZ0Z_1 ;
    wire \ppm_encoder_1.elevatorZ0Z_11 ;
    wire \ppm_encoder_1.elevatorZ0Z_2 ;
    wire \ppm_encoder_1.rudderZ0Z_11 ;
    wire bfn_7_9_0_;
    wire \ppm_encoder_1.un1_rudder_cry_6_THRU_CO ;
    wire \ppm_encoder_1.un1_rudder_cry_6 ;
    wire \ppm_encoder_1.un1_rudder_cry_7 ;
    wire \ppm_encoder_1.un1_rudder_cry_8_THRU_CO ;
    wire \ppm_encoder_1.un1_rudder_cry_8 ;
    wire \ppm_encoder_1.un1_rudder_cry_9 ;
    wire \ppm_encoder_1.un1_rudder_cry_10_THRU_CO ;
    wire \ppm_encoder_1.un1_rudder_cry_10 ;
    wire \ppm_encoder_1.un1_rudder_cry_11 ;
    wire \ppm_encoder_1.un1_rudder_cry_12 ;
    wire \ppm_encoder_1.un1_rudder_cry_13 ;
    wire bfn_7_10_0_;
    wire bfn_7_11_0_;
    wire \scaler_4.un2_source_data_0_cry_1 ;
    wire scaler_4_data_7;
    wire \scaler_4.un2_source_data_0_cry_2 ;
    wire \scaler_4.un2_source_data_0_cry_3 ;
    wire scaler_4_data_9;
    wire \scaler_4.un2_source_data_0_cry_4 ;
    wire \scaler_4.un2_source_data_0_cry_5 ;
    wire scaler_4_data_11;
    wire \scaler_4.un2_source_data_0_cry_6 ;
    wire \scaler_4.un2_source_data_0_cry_7 ;
    wire \scaler_4.un2_source_data_0_cry_8 ;
    wire bfn_7_12_0_;
    wire \scaler_4.un2_source_data_0_cry_9 ;
    wire scaler_4_data_14;
    wire \Commands_frame_decoder.preinit_RNIHOVZ0Z81_cascade_ ;
    wire \Commands_frame_decoder.WDT_RNIHV6PZ0Z_11_cascade_ ;
    wire \Commands_frame_decoder.WDT_RNIET8A1_0Z0Z_4 ;
    wire \Commands_frame_decoder.WDT_RNI30853Z0Z_10 ;
    wire \Commands_frame_decoder.preinitZ0 ;
    wire \Commands_frame_decoder.WDT_RNI2VDI1Z0Z_10 ;
    wire \Commands_frame_decoder.WDT_RNITK4L_0Z0Z_8 ;
    wire \Commands_frame_decoder.WDT_RNIET8A1Z0Z_4_cascade_ ;
    wire \Commands_frame_decoder.WDT_RNIHV6P_0Z0Z_11 ;
    wire \Commands_frame_decoder.WDT8lt14_0_cascade_ ;
    wire \Commands_frame_decoder.N_365_0_cascade_ ;
    wire \Commands_frame_decoder.WDT_RNITK4LZ0Z_8 ;
    wire \pid_front.O_0_13 ;
    wire \uart_pc.stateZ0Z_1 ;
    wire \uart_pc.state_srsts_i_0_2_cascade_ ;
    wire \uart_pc.N_144_1_cascade_ ;
    wire \Commands_frame_decoder.count_1_sqmuxa ;
    wire \uart_pc.stateZ0Z_2 ;
    wire \uart_pc.N_145 ;
    wire \Commands_frame_decoder.N_370_2 ;
    wire \Commands_frame_decoder.N_371 ;
    wire \Commands_frame_decoder.N_370_2_cascade_ ;
    wire \Commands_frame_decoder.state_ns_i_0_0_cascade_ ;
    wire \Commands_frame_decoder.N_372 ;
    wire \Commands_frame_decoder.state_RNO_0Z0Z_14_cascade_ ;
    wire \Commands_frame_decoder.N_365_0 ;
    wire \Commands_frame_decoder.stateZ0Z_2 ;
    wire \uart_pc.state_srsts_0_0_0_cascade_ ;
    wire \uart_pc.stateZ0Z_0 ;
    wire \uart_pc.N_126_li_cascade_ ;
    wire bfn_7_19_0_;
    wire \uart_pc.timer_CountZ1Z_2 ;
    wire \uart_pc.timer_Count_RNO_0Z0Z_2 ;
    wire \uart_pc.un4_timer_Count_1_cry_1 ;
    wire \uart_pc.un4_timer_Count_1_cry_2 ;
    wire \uart_pc.un4_timer_Count_1_cry_3 ;
    wire \uart_pc.timer_Count_RNO_0Z0Z_4 ;
    wire \uart_pc.timer_CountZ0Z_4 ;
    wire \uart_pc.timer_Count_RNO_0Z0Z_3 ;
    wire \uart_pc.timer_CountZ1Z_3 ;
    wire \uart_pc.timer_CountZ0Z_0 ;
    wire \uart_pc.timer_Count_0_sqmuxa ;
    wire \uart_pc.timer_Count_RNO_0Z0Z_1_cascade_ ;
    wire \uart_pc.timer_CountZ1Z_1 ;
    wire \Commands_frame_decoder.stateZ0Z_14 ;
    wire \Commands_frame_decoder.countZ0Z_0 ;
    wire \uart_pc.N_144_1 ;
    wire \uart_pc.N_143 ;
    wire \Commands_frame_decoder.stateZ0Z_0 ;
    wire \Commands_frame_decoder.state_ns_0_a3_3_1 ;
    wire \pid_front.state_0_0 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5I0L2Z0Z_3 ;
    wire bfn_8_1_0_;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_1 ;
    wire \ppm_encoder_1.un1_init_pulses_11_1 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_0 ;
    wire \ppm_encoder_1.init_pulses_RNIHGIP3Z0Z_2 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_1 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_3 ;
    wire \ppm_encoder_1.un1_init_pulses_11_3 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_2 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_4 ;
    wire \ppm_encoder_1.un1_init_pulses_11_4 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_3 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_5 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_4 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_5 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_7 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_6 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_7 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_8 ;
    wire bfn_8_2_0_;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_9 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_8 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_10 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_9 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_10 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_12 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_11 ;
    wire \ppm_encoder_1.init_pulses_RNIOHJF3Z0Z_13 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_12 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_14 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_13 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_15 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_14 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_15 ;
    wire bfn_8_3_0_;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_16 ;
    wire \ppm_encoder_1.PPM_STATE_RNIMINSZ0Z_0 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_17 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_11 ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_13 ;
    wire \ppm_encoder_1.N_254_i_i_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_17 ;
    wire \ppm_encoder_1.un1_init_pulses_11_16 ;
    wire \ppm_encoder_1.un1_init_pulses_11_10 ;
    wire \ppm_encoder_1.N_298_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_11_17 ;
    wire \ppm_encoder_1.un1_init_pulses_11_18 ;
    wire \ppm_encoder_1.un1_init_pulses_11_13 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_13 ;
    wire \ppm_encoder_1.un1_init_pulses_11_14 ;
    wire \ppm_encoder_1.un1_init_pulses_11_15 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3 ;
    wire \ppm_encoder_1.N_257_i_i_cascade_ ;
    wire throttle_order_0;
    wire \ppm_encoder_1.N_266_i ;
    wire \ppm_encoder_1.aileronZ0Z_0 ;
    wire \ppm_encoder_1.throttleZ0Z_0 ;
    wire \ppm_encoder_1.aileronZ0Z_10 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ;
    wire \ppm_encoder_1.N_508_cascade_ ;
    wire throttle_order_12;
    wire \ppm_encoder_1.un1_throttle_cry_11_THRU_CO ;
    wire \ppm_encoder_1.elevatorZ0Z_10 ;
    wire \ppm_encoder_1.un1_rudder_cry_7_THRU_CO ;
    wire scaler_4_data_8;
    wire \ppm_encoder_1.elevatorZ0Z_13 ;
    wire \ppm_encoder_1.un1_rudder_cry_9_THRU_CO ;
    wire scaler_4_data_10;
    wire \ppm_encoder_1.un1_rudder_cry_12_THRU_CO ;
    wire scaler_4_data_13;
    wire \ppm_encoder_1.rudderZ0Z_13 ;
    wire scaler_4_data_12;
    wire \ppm_encoder_1.un1_rudder_cry_11_THRU_CO ;
    wire \ppm_encoder_1.rudderZ0Z_12 ;
    wire bfn_8_11_0_;
    wire frame_decoder_CH4data_1;
    wire \scaler_4.un3_source_data_0_cry_0 ;
    wire frame_decoder_CH4data_2;
    wire \scaler_4.un3_source_data_0_cry_1_c_RNI74CL ;
    wire \scaler_4.un3_source_data_0_cry_1 ;
    wire frame_decoder_CH4data_3;
    wire \scaler_4.un3_source_data_0_cry_2_c_RNIA8DL ;
    wire \scaler_4.un3_source_data_0_cry_2 ;
    wire frame_decoder_CH4data_4;
    wire \scaler_4.un3_source_data_0_cry_3_c_RNIDCEL ;
    wire \scaler_4.un3_source_data_0_cry_3 ;
    wire frame_decoder_CH4data_5;
    wire \scaler_4.un3_source_data_0_cry_4_c_RNIGGFL ;
    wire \scaler_4.un3_source_data_0_cry_4 ;
    wire frame_decoder_CH4data_6;
    wire \scaler_4.un3_source_data_0_cry_5_c_RNIJKGL ;
    wire \scaler_4.un3_source_data_0_cry_5 ;
    wire \scaler_4.un3_source_data_0_cry_6_c_RNIOUNN ;
    wire \scaler_4.un3_source_data_0_cry_6 ;
    wire \scaler_4.un3_source_data_0_cry_7 ;
    wire \scaler_4.un3_source_data_0_cry_7_c_RNIP0PN ;
    wire bfn_8_12_0_;
    wire \scaler_4.un3_source_data_0_cry_8 ;
    wire \scaler_4.un3_source_data_0_cry_8_c_RNIS918 ;
    wire \Commands_frame_decoder.state_RNIQRI31Z0Z_10 ;
    wire \scaler_4.un3_source_data_0_axb_7 ;
    wire \Commands_frame_decoder.state_0_sqmuxa ;
    wire \Commands_frame_decoder.WDTZ0Z_0 ;
    wire bfn_8_13_0_;
    wire \Commands_frame_decoder.WDTZ0Z_1 ;
    wire \Commands_frame_decoder.un1_WDT_cry_0 ;
    wire \Commands_frame_decoder.WDTZ0Z_2 ;
    wire \Commands_frame_decoder.un1_WDT_cry_1 ;
    wire \Commands_frame_decoder.WDTZ0Z_3 ;
    wire \Commands_frame_decoder.un1_WDT_cry_2 ;
    wire \Commands_frame_decoder.WDTZ0Z_4 ;
    wire \Commands_frame_decoder.un1_WDT_cry_3 ;
    wire \Commands_frame_decoder.WDTZ0Z_5 ;
    wire \Commands_frame_decoder.un1_WDT_cry_4 ;
    wire \Commands_frame_decoder.WDTZ0Z_6 ;
    wire \Commands_frame_decoder.un1_WDT_cry_5 ;
    wire \Commands_frame_decoder.WDTZ0Z_7 ;
    wire \Commands_frame_decoder.un1_WDT_cry_6 ;
    wire \Commands_frame_decoder.un1_WDT_cry_7 ;
    wire \Commands_frame_decoder.WDTZ0Z_8 ;
    wire bfn_8_14_0_;
    wire \Commands_frame_decoder.WDTZ0Z_9 ;
    wire \Commands_frame_decoder.un1_WDT_cry_8 ;
    wire \Commands_frame_decoder.WDTZ0Z_10 ;
    wire \Commands_frame_decoder.un1_WDT_cry_9 ;
    wire \Commands_frame_decoder.WDTZ0Z_11 ;
    wire \Commands_frame_decoder.un1_WDT_cry_10 ;
    wire \Commands_frame_decoder.WDTZ0Z_12 ;
    wire \Commands_frame_decoder.un1_WDT_cry_11 ;
    wire \Commands_frame_decoder.WDTZ0Z_13 ;
    wire \Commands_frame_decoder.un1_WDT_cry_12 ;
    wire \Commands_frame_decoder.un1_WDT_cry_13 ;
    wire \Commands_frame_decoder.un1_WDT_cry_14 ;
    wire scaler_4_data_5;
    wire \uart_pc.N_152_cascade_ ;
    wire \uart_pc.CO0_cascade_ ;
    wire \uart_pc.un1_state_7_0 ;
    wire \uart_pc.un1_state_4_0 ;
    wire \uart_pc.bit_CountZ0Z_0 ;
    wire \uart_pc.bit_CountZ0Z_1 ;
    wire \uart_pc.bit_CountZ0Z_2 ;
    wire \uart_pc.timer_Count_RNILR1B2Z0Z_2_cascade_ ;
    wire \Commands_frame_decoder.state_ns_i_a2_2_1Z0Z_0_cascade_ ;
    wire \Commands_frame_decoder.N_410 ;
    wire \uart_pc.timer_Count_RNIMQ8T1Z0Z_2_cascade_ ;
    wire \dron_frame_decoder_1.WDTZ0Z_0 ;
    wire bfn_8_18_0_;
    wire \dron_frame_decoder_1.WDTZ0Z_1 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_0 ;
    wire \dron_frame_decoder_1.WDTZ0Z_2 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_1 ;
    wire \dron_frame_decoder_1.WDTZ0Z_3 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_2 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_3 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_4 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_5 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_6 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_7 ;
    wire bfn_8_19_0_;
    wire \dron_frame_decoder_1.un1_WDT_cry_8 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_9 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_10 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_11 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_12 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_13 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_14 ;
    wire \dron_frame_decoder_1.source_data_valid_2_sqmuxa_iZ0 ;
    wire \dron_frame_decoder_1.WDTZ0Z_6 ;
    wire \dron_frame_decoder_1.WDTZ0Z_7 ;
    wire \dron_frame_decoder_1.WDTZ0Z_10 ;
    wire \dron_frame_decoder_1.WDT10lt12_0_cascade_ ;
    wire \dron_frame_decoder_1.WDT10_0_i ;
    wire \dron_frame_decoder_1.WDT10_0_i_1 ;
    wire \dron_frame_decoder_1.WDTZ0Z_8 ;
    wire \dron_frame_decoder_1.WDTZ0Z_5 ;
    wire \dron_frame_decoder_1.WDTZ0Z_9 ;
    wire \dron_frame_decoder_1.WDTZ0Z_4 ;
    wire \dron_frame_decoder_1.WDT10lto9_3 ;
    wire \dron_frame_decoder_1.WDTZ0Z_11 ;
    wire \dron_frame_decoder_1.WDTZ0Z_12 ;
    wire \dron_frame_decoder_1.WDTZ0Z_13 ;
    wire \dron_frame_decoder_1.WDT10lt12_0 ;
    wire \dron_frame_decoder_1.WDTZ0Z_14 ;
    wire \dron_frame_decoder_1.WDT10lt14_0_cascade_ ;
    wire \dron_frame_decoder_1.WDTZ0Z_15 ;
    wire \dron_frame_decoder_1.N_218_cascade_ ;
    wire \dron_frame_decoder_1.stateZ0Z_2 ;
    wire \ppm_encoder_1.N_262_i_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_6_cascade_ ;
    wire \ppm_encoder_1.elevatorZ0Z_6 ;
    wire scaler_4_data_6;
    wire \ppm_encoder_1.rudderZ0Z_6 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z1 ;
    wire \ppm_encoder_1.N_262_i_i_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_6 ;
    wire \ppm_encoder_1.init_pulses_RNIQOIP3Z0Z_6 ;
    wire bfn_9_2_0_;
    wire \ppm_encoder_1.init_pulses_RNI29LM5Z0Z_1 ;
    wire \ppm_encoder_1.N_258_i_i ;
    wire \ppm_encoder_1.un1_init_pulses_10_1 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_0 ;
    wire \ppm_encoder_1.init_pulses_RNIIIS46Z0Z_2 ;
    wire \ppm_encoder_1.N_259_i_i ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_1 ;
    wire \ppm_encoder_1.init_pulses_RNINNS46Z0Z_3 ;
    wire \ppm_encoder_1.N_256_i_i ;
    wire \ppm_encoder_1.un1_init_pulses_10_3 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_2 ;
    wire \ppm_encoder_1.init_pulses_RNIFTCL6Z0Z_4 ;
    wire \ppm_encoder_1.N_260_i_i ;
    wire \ppm_encoder_1.un1_init_pulses_10_4 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_3 ;
    wire \ppm_encoder_1.init_pulses_RNI3K6R5Z0Z_5 ;
    wire \ppm_encoder_1.N_261_i_i ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_4 ;
    wire \ppm_encoder_1.init_pulses_RNI20JF6Z0Z_6 ;
    wire \ppm_encoder_1.N_262_i_i ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_5 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_6 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_7 ;
    wire \ppm_encoder_1.init_pulses_RNIL76H6Z0Z_8 ;
    wire \ppm_encoder_1.N_264_i_i ;
    wire bfn_9_3_0_;
    wire \ppm_encoder_1.init_pulses_RNIOCUG6Z0Z_9 ;
    wire \ppm_encoder_1.N_265_i_i ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_8 ;
    wire \ppm_encoder_1.init_pulses_RNI8E326Z0Z_10 ;
    wire \ppm_encoder_1.N_255_i_i ;
    wire \ppm_encoder_1.un1_init_pulses_10_10 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_9 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_10 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_11 ;
    wire \ppm_encoder_1.init_pulses_RNI8L3H5Z0Z_13 ;
    wire \ppm_encoder_1.N_268_i_i ;
    wire \ppm_encoder_1.un1_init_pulses_10_13 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_12 ;
    wire \ppm_encoder_1.un1_init_pulses_10_14 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_13 ;
    wire \ppm_encoder_1.init_pulses_RNILFR51Z0Z_15 ;
    wire \ppm_encoder_1.N_254_i_i ;
    wire \ppm_encoder_1.un1_init_pulses_10_15 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_14 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_15 ;
    wire \ppm_encoder_1.un1_init_pulses_10_16 ;
    wire bfn_9_4_0_;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_17 ;
    wire \ppm_encoder_1.un1_init_pulses_10_17 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_16 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_17 ;
    wire \ppm_encoder_1.un1_init_pulses_10_18 ;
    wire \ppm_encoder_1.init_pulses_4_sqmuxa_i_0_0_0 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_1_0 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_0_0 ;
    wire \ppm_encoder_1.N_257_i_i ;
    wire \ppm_encoder_1.throttle_RNI0EA05Z0Z_0 ;
    wire \ppm_encoder_1.N_266_i_i ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_11 ;
    wire \ppm_encoder_1.init_pulses_RNIU1F76Z0Z_11 ;
    wire \ppm_encoder_1.N_263_i_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_7_cascade_ ;
    wire \ppm_encoder_1.init_pulses_RNISD9M6Z0Z_7 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_0_0_7 ;
    wire \ppm_encoder_1.rudderZ0Z_7 ;
    wire \ppm_encoder_1.N_263_i_i ;
    wire \ppm_encoder_1.N_293 ;
    wire \ppm_encoder_1.N_507 ;
    wire \ppm_encoder_1.N_509 ;
    wire \ppm_encoder_1.un2_throttle_iv_i_i_0_14_cascade_ ;
    wire \ppm_encoder_1.N_303 ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_14_cascade_ ;
    wire \ppm_encoder_1.init_pulses_RNIP98N6Z0Z_14 ;
    wire \ppm_encoder_1.rudderZ0Z_14 ;
    wire \ppm_encoder_1.N_269_i_i ;
    wire \ppm_encoder_1.pulses2count_9_0_0_11 ;
    wire \ppm_encoder_1.N_431 ;
    wire \ppm_encoder_1.N_269_i ;
    wire \ppm_encoder_1.throttleZ0Z_6 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_3 ;
    wire \ppm_encoder_1.aileronZ0Z_8 ;
    wire \ppm_encoder_1.elevatorZ0Z_8 ;
    wire \ppm_encoder_1.aileronZ0Z_9 ;
    wire \ppm_encoder_1.pulses2count_9_i_1_9 ;
    wire \ppm_encoder_1.elevatorZ0Z_9 ;
    wire \ppm_encoder_1.un1_throttle_cry_6_THRU_CO ;
    wire throttle_order_7;
    wire throttle_order_8;
    wire \ppm_encoder_1.un1_throttle_cry_7_THRU_CO ;
    wire \ppm_encoder_1.throttleZ0Z_8 ;
    wire throttle_order_9;
    wire \ppm_encoder_1.un1_throttle_cry_8_THRU_CO ;
    wire \ppm_encoder_1.throttleZ0Z_9 ;
    wire \ppm_encoder_1.aileronZ0Z_6 ;
    wire \uart_drone.N_126_li_cascade_ ;
    wire \uart_drone.N_143_cascade_ ;
    wire \scaler_4.un2_source_data_0 ;
    wire frame_decoder_CH4data_0;
    wire \scaler_4.un2_source_data_0_cry_1_c_RNOZ0 ;
    wire \pid_alt.N_933_0 ;
    wire frame_decoder_OFF4data_0;
    wire frame_decoder_OFF4data_1;
    wire frame_decoder_OFF4data_2;
    wire frame_decoder_OFF4data_3;
    wire frame_decoder_OFF4data_4;
    wire frame_decoder_OFF4data_5;
    wire frame_decoder_OFF4data_6;
    wire xy_kp_0;
    wire xy_kp_1;
    wire xy_kp_2;
    wire xy_kp_3;
    wire xy_kp_5;
    wire xy_kp_6;
    wire xy_kp_7;
    wire \uart_pc.N_152 ;
    wire \uart_pc.data_AuxZ0Z_7 ;
    wire \Commands_frame_decoder.un1_sink_data_valid_2_0_0 ;
    wire \Commands_frame_decoder.source_offset4data_1_sqmuxa ;
    wire \Commands_frame_decoder.source_offset4data_1_sqmuxa_cascade_ ;
    wire \Commands_frame_decoder.source_offset4data_1_sqmuxa_0 ;
    wire \Commands_frame_decoder.source_CH4data_1_sqmuxa_0 ;
    wire \uart_pc.N_126_li ;
    wire \uart_pc.stateZ0Z_4 ;
    wire \uart_pc.un1_state_2_0_a3_0 ;
    wire \uart_pc.stateZ0Z_3 ;
    wire \uart_pc.un1_state_2_0_cascade_ ;
    wire \uart_pc.data_Auxce_0_0_0 ;
    wire \uart_pc.data_Auxce_0_1 ;
    wire \uart_pc.data_Auxce_0_0_2 ;
    wire \uart_pc.data_Auxce_0_3 ;
    wire \uart_pc.data_AuxZ0Z_3 ;
    wire \uart_pc.data_Auxce_0_0_4 ;
    wire \uart_pc.data_AuxZ0Z_4 ;
    wire \uart_pc.data_Auxce_0_5 ;
    wire \uart_pc.un1_state_2_0 ;
    wire \uart_pc.data_Auxce_0_6 ;
    wire \uart_pc.data_AuxZ0Z_6 ;
    wire \uart_pc.state_RNIEAGSZ0Z_4 ;
    wire \uart_pc.data_AuxZ1Z_2 ;
    wire \Commands_frame_decoder.state_ns_0_a3_0_1Z0Z_2_cascade_ ;
    wire \Commands_frame_decoder.stateZ0Z_1 ;
    wire \Commands_frame_decoder.N_406 ;
    wire \uart_pc.data_AuxZ1Z_0 ;
    wire \uart_pc.data_AuxZ0Z_5 ;
    wire \uart_pc.timer_Count_RNILR1B2Z0Z_2 ;
    wire \uart_pc.timer_Count_RNIMQ8T1Z0Z_2 ;
    wire \uart_pc.data_AuxZ1Z_1 ;
    wire \pid_alt.drone_altitude_i_0 ;
    wire frame_decoder_OFF4data_7;
    wire frame_decoder_CH4data_7;
    wire \scaler_4.N_2928_i_l_ofxZ0 ;
    wire drone_altitude_i_4;
    wire drone_altitude_i_5;
    wire drone_altitude_i_6;
    wire drone_altitude_i_7;
    wire xy_kd_1;
    wire drone_altitude_i_9;
    wire \dron_frame_decoder_1.state_RNI4N6KZ0Z_2 ;
    wire \dron_frame_decoder_1.un1_sink_data_valid_5_i_0 ;
    wire \dron_frame_decoder_1.un1_sink_data_valid_5_i_0_cascade_ ;
    wire \dron_frame_decoder_1.stateZ0Z_4 ;
    wire \dron_frame_decoder_1.stateZ0Z_5 ;
    wire \dron_frame_decoder_1.state_ns_0_i_a2_0_2_3_cascade_ ;
    wire \dron_frame_decoder_1.stateZ0Z_3 ;
    wire \dron_frame_decoder_1.state_ns_0_i_a2_0_3_3 ;
    wire \dron_frame_decoder_1.stateZ0Z_6 ;
    wire \pid_alt.state_RNIFCSD1Z0Z_0 ;
    wire \Commands_frame_decoder.state_ns_0_a3_0_1 ;
    wire \pid_front.O_0_6 ;
    wire bfn_10_1_0_;
    wire \ppm_encoder_1.counter24_0_data_tmp_0 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_1 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_2 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_3 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_4 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_5 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_6 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_7 ;
    wire bfn_10_2_0_;
    wire \ppm_encoder_1.counter24_0_data_tmp_8 ;
    wire \ppm_encoder_1.counter24_0_N_2 ;
    wire \ppm_encoder_1.counter24_0_I_51_c_RNOZ0 ;
    wire \ppm_encoder_1.counter24_0_I_39_c_RNOZ0 ;
    wire \ppm_encoder_1.un1_init_pulses_11_2 ;
    wire \ppm_encoder_1.un1_init_pulses_10_2 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_2 ;
    wire \ppm_encoder_1.un1_init_pulses_11_5 ;
    wire \ppm_encoder_1.un1_init_pulses_10_5 ;
    wire \ppm_encoder_1.un1_init_pulses_11_6 ;
    wire \ppm_encoder_1.un1_init_pulses_10_6 ;
    wire \ppm_encoder_1.un1_init_pulses_11_7 ;
    wire \ppm_encoder_1.un1_init_pulses_10_7 ;
    wire \ppm_encoder_1.un1_init_pulses_10_9 ;
    wire \ppm_encoder_1.un1_init_pulses_11_9 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_9 ;
    wire \ppm_encoder_1.throttleZ0Z_10 ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_16 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_16 ;
    wire \ppm_encoder_1.un1_init_pulses_11_8 ;
    wire \ppm_encoder_1.un1_init_pulses_10_8 ;
    wire \ppm_encoder_1.un1_init_pulses_11_11 ;
    wire \ppm_encoder_1.un1_init_pulses_10_11 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_11 ;
    wire \ppm_encoder_1.un1_init_pulses_11_12 ;
    wire \ppm_encoder_1.un1_init_pulses_10_12 ;
    wire \ppm_encoder_1.aileronZ0Z_4 ;
    wire \ppm_encoder_1.elevatorZ0Z_4 ;
    wire \ppm_encoder_1.elevatorZ0Z_0 ;
    wire \ppm_encoder_1.N_393 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_ns_0 ;
    wire \ppm_encoder_1.N_56 ;
    wire \ppm_encoder_1.N_378 ;
    wire \ppm_encoder_1.rudderZ0Z_10 ;
    wire \ppm_encoder_1.N_406 ;
    wire scaler_4_data_4;
    wire \ppm_encoder_1.rudderZ0Z_4 ;
    wire \ppm_encoder_1.N_420 ;
    wire \ppm_encoder_1.rudderZ0Z_8 ;
    wire \ppm_encoder_1.rudderZ0Z_9 ;
    wire \ppm_encoder_1.N_425 ;
    wire \ppm_encoder_1.pulses2count_9_i_2_9 ;
    wire \ppm_encoder_1.N_275 ;
    wire \ppm_encoder_1.elevatorZ0Z_3 ;
    wire \ppm_encoder_1.N_513 ;
    wire \ppm_encoder_1.N_300 ;
    wire \ppm_encoder_1.pulses2count_9_0_0_0_3 ;
    wire bfn_10_7_0_;
    wire \ppm_encoder_1.un1_elevator_cry_0_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_0 ;
    wire \ppm_encoder_1.un1_elevator_cry_1_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_1 ;
    wire \ppm_encoder_1.un1_elevator_cry_2_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_2 ;
    wire \ppm_encoder_1.un1_elevator_cry_3_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_3 ;
    wire \ppm_encoder_1.un1_elevator_cry_4 ;
    wire \ppm_encoder_1.un1_elevator_cry_5_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_5 ;
    wire \ppm_encoder_1.un1_elevator_cry_6 ;
    wire \ppm_encoder_1.un1_elevator_cry_7 ;
    wire \ppm_encoder_1.un1_elevator_cry_7_THRU_CO ;
    wire bfn_10_8_0_;
    wire \ppm_encoder_1.un1_elevator_cry_8_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_8 ;
    wire \ppm_encoder_1.un1_elevator_cry_9_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_9 ;
    wire \ppm_encoder_1.un1_elevator_cry_10_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_10 ;
    wire \ppm_encoder_1.un1_elevator_cry_11_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_11 ;
    wire \ppm_encoder_1.un1_elevator_cry_12_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_12 ;
    wire \ppm_encoder_1.un1_elevator_cry_13 ;
    wire \ppm_encoder_1.elevatorZ0Z_14 ;
    wire \uart_drone.N_152_cascade_ ;
    wire \uart_drone.un1_state_7_0 ;
    wire \uart_drone.CO0 ;
    wire \ppm_encoder_1.throttleZ0Z_12 ;
    wire bfn_10_10_0_;
    wire \ppm_encoder_1.un1_aileron_cry_0_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_0 ;
    wire \ppm_encoder_1.un1_aileron_cry_1_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_1 ;
    wire \ppm_encoder_1.un1_aileron_cry_2_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_2 ;
    wire \ppm_encoder_1.un1_aileron_cry_3_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_3 ;
    wire \ppm_encoder_1.un1_aileron_cry_4_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_4 ;
    wire \ppm_encoder_1.un1_aileron_cry_5_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_5 ;
    wire \ppm_encoder_1.un1_aileron_cry_6_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_6 ;
    wire \ppm_encoder_1.un1_aileron_cry_7 ;
    wire \ppm_encoder_1.un1_aileron_cry_7_THRU_CO ;
    wire bfn_10_11_0_;
    wire \ppm_encoder_1.un1_aileron_cry_8_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_8 ;
    wire \ppm_encoder_1.un1_aileron_cry_9_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_9 ;
    wire \ppm_encoder_1.un1_aileron_cry_10_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_10 ;
    wire \ppm_encoder_1.un1_aileron_cry_11_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_11 ;
    wire \ppm_encoder_1.un1_aileron_cry_12 ;
    wire \ppm_encoder_1.un1_aileron_cry_13 ;
    wire \ppm_encoder_1.pid_altitude_dv_0 ;
    wire \uart_drone.timer_CountZ0Z_0 ;
    wire bfn_10_12_0_;
    wire \uart_drone.timer_CountZ1Z_2 ;
    wire \uart_drone.timer_Count_RNO_0_0_2 ;
    wire \uart_drone.un4_timer_Count_1_cry_1 ;
    wire \uart_drone.un4_timer_Count_1_cry_2 ;
    wire \uart_drone.un4_timer_Count_1_cry_3 ;
    wire \uart_drone.data_rdyc_1 ;
    wire \uart_drone.timer_Count_RNO_0_0_4 ;
    wire \uart_drone.timer_Count_RNO_0_0_3 ;
    wire \uart_drone_sync.aux_1__0__0_0 ;
    wire \uart_pc_sync.aux_1__0_Z0Z_0 ;
    wire \uart_pc_sync.aux_2__0_Z0Z_0 ;
    wire \uart_pc_sync.aux_3__0_Z0Z_0 ;
    wire debug_CH3_20A_c;
    wire \scaler_4.debug_CH3_20A_c_0 ;
    wire \Commands_frame_decoder.state_RNIG48SZ0Z_7 ;
    wire \Commands_frame_decoder.WDT8lt14_0 ;
    wire \Commands_frame_decoder.WDTZ0Z_15 ;
    wire \Commands_frame_decoder.WDTZ0Z_14 ;
    wire \Commands_frame_decoder.stateZ0Z_10 ;
    wire \Commands_frame_decoder.N_403_cascade_ ;
    wire \Commands_frame_decoder.stateZ0Z_8 ;
    wire \Commands_frame_decoder.stateZ0Z_9 ;
    wire \pid_alt.error_axbZ0Z_1 ;
    wire \pid_alt.error_axbZ0Z_12 ;
    wire drone_altitude_0;
    wire drone_altitude_1;
    wire \dron_frame_decoder_1.drone_altitude_4 ;
    wire \dron_frame_decoder_1.drone_altitude_5 ;
    wire \dron_frame_decoder_1.drone_altitude_6 ;
    wire \dron_frame_decoder_1.drone_altitude_7 ;
    wire \dron_frame_decoder_1.N_740_0 ;
    wire drone_altitude_12;
    wire drone_altitude_15;
    wire \dron_frame_decoder_1.drone_altitude_8 ;
    wire \dron_frame_decoder_1.drone_altitude_9 ;
    wire \Commands_frame_decoder.state_RNIF38SZ0Z_6 ;
    wire \dron_frame_decoder_1.state_RNI3T3K1Z0Z_7 ;
    wire \dron_frame_decoder_1.drone_altitude_10 ;
    wire drone_altitude_i_10;
    wire \Commands_frame_decoder.stateZ0Z_13 ;
    wire \Commands_frame_decoder.stateZ0Z_12 ;
    wire \Commands_frame_decoder.source_xy_ki_1_sqmuxa ;
    wire \Commands_frame_decoder.source_xy_ki_1_sqmuxa_cascade_ ;
    wire \dron_frame_decoder_1.N_230_5 ;
    wire \dron_frame_decoder_1.N_230_5_cascade_ ;
    wire uart_drone_data_rdy;
    wire \dron_frame_decoder_1.state_ns_i_a2_0_1_0 ;
    wire \dron_frame_decoder_1.N_224_cascade_ ;
    wire \dron_frame_decoder_1.state_ns_i_a2_1_1Z0Z_0_cascade_ ;
    wire \dron_frame_decoder_1.N_220 ;
    wire \dron_frame_decoder_1.N_224 ;
    wire \dron_frame_decoder_1.N_220_cascade_ ;
    wire \dron_frame_decoder_1.stateZ0Z_1 ;
    wire \dron_frame_decoder_1.N_200 ;
    wire \dron_frame_decoder_1.N_198 ;
    wire \dron_frame_decoder_1.stateZ0Z_0 ;
    wire \dron_frame_decoder_1.state_ns_i_a2_0_2_0 ;
    wire \ppm_encoder_1.counter24_0_I_15_c_RNOZ0 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_15 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_14 ;
    wire \ppm_encoder_1.N_309 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_16 ;
    wire \ppm_encoder_1.pulses2countZ0Z_16 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_17 ;
    wire \ppm_encoder_1.pulses2countZ0Z_17 ;
    wire \ppm_encoder_1.counter24_0_I_21_c_RNOZ0 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_6 ;
    wire \ppm_encoder_1.N_306 ;
    wire \ppm_encoder_1.pulses2countZ0Z_6 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_7 ;
    wire \ppm_encoder_1.N_310 ;
    wire \ppm_encoder_1.pulses2countZ0Z_7 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_18 ;
    wire \ppm_encoder_1.pulses2countZ0Z_18 ;
    wire \ppm_encoder_1.counter24_0_I_57_c_RNOZ0 ;
    wire \ppm_encoder_1.pulses2count_9_i_2_8 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_8 ;
    wire \ppm_encoder_1.pulses2count_9_i_1_8 ;
    wire \ppm_encoder_1.pulses2countZ0Z_8 ;
    wire \ppm_encoder_1.pulses2countZ0Z_9 ;
    wire \ppm_encoder_1.counter24_0_I_27_c_RNOZ0 ;
    wire \ppm_encoder_1.counter24_0_I_57_c_RNIJMMDZ0 ;
    wire \ppm_encoder_1.counter24_0_I_57_c_RNIJMMDZ0_cascade_ ;
    wire \ppm_encoder_1.N_500 ;
    wire ppm_output_c;
    wire \ppm_encoder_1.N_486_9 ;
    wire \ppm_encoder_1.PPM_STATEZ0Z_1 ;
    wire \ppm_encoder_1.N_486 ;
    wire \ppm_encoder_1.N_486_cascade_ ;
    wire \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ;
    wire \ppm_encoder_1.counter24_0_N_2_THRU_CO ;
    wire \ppm_encoder_1.PPM_STATEZ0Z_0 ;
    wire \ppm_encoder_1.N_374 ;
    wire \ppm_encoder_1.N_298 ;
    wire \ppm_encoder_1.un1_init_pulses_11_0 ;
    wire \ppm_encoder_1.N_374_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_10_0 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_0 ;
    wire \ppm_encoder_1.counter24_0_I_1_c_RNOZ0 ;
    wire \ppm_encoder_1.pulses2count_9_0_3_1 ;
    wire \ppm_encoder_1.aileronZ0Z_1 ;
    wire \ppm_encoder_1.pulses2countZ0Z_1 ;
    wire \ppm_encoder_1.pulses2count_9_0_3_11 ;
    wire \ppm_encoder_1.aileronZ0Z_11 ;
    wire \ppm_encoder_1.pulses2countZ0Z_11 ;
    wire \ppm_encoder_1.counter24_0_I_33_c_RNOZ0 ;
    wire \ppm_encoder_1.pulses2count_9_i_0_2_10 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_10 ;
    wire \ppm_encoder_1.pulses2count_9_i_0_1_10 ;
    wire \ppm_encoder_1.pulses2countZ0Z_10 ;
    wire \ppm_encoder_1.pulses2count_9_0_0_0 ;
    wire \ppm_encoder_1.pulses2count_9_0_2_0 ;
    wire \ppm_encoder_1.pulses2countZ0Z_0 ;
    wire \ppm_encoder_1.pulses2count_9_i_2_4 ;
    wire \ppm_encoder_1.pulses2count_9_i_1_4 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_4 ;
    wire \ppm_encoder_1.pulses2countZ0Z_4 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_5 ;
    wire \ppm_encoder_1.N_307 ;
    wire \ppm_encoder_1.pulses2countZ0Z_5 ;
    wire \ppm_encoder_1.pulses2count_9_0_1_13 ;
    wire \ppm_encoder_1.un2_throttle_0_2_13 ;
    wire \ppm_encoder_1.pulses2countZ0Z_13 ;
    wire \ppm_encoder_1.aileronZ0Z_12 ;
    wire \ppm_encoder_1.pulses2countZ0Z_12 ;
    wire \ppm_encoder_1.pulses2count_9_i_3_2 ;
    wire \ppm_encoder_1.aileronZ0Z_2 ;
    wire \ppm_encoder_1.pulses2count_9_0_0_1_3 ;
    wire \ppm_encoder_1.N_514 ;
    wire \ppm_encoder_1.throttleZ0Z_3 ;
    wire \ppm_encoder_1.N_529 ;
    wire \ppm_encoder_1.N_304 ;
    wire \ppm_encoder_1.pulses2count_9_0_0_3_3_cascade_ ;
    wire \ppm_encoder_1.aileronZ0Z_3 ;
    wire \ppm_encoder_1.N_295_i_0 ;
    wire \ppm_encoder_1.pulses2countZ0Z_2 ;
    wire \ppm_encoder_1.pulses2countZ0Z_3 ;
    wire \ppm_encoder_1.counter24_0_I_9_c_RNOZ0 ;
    wire \ppm_encoder_1.un1_elevator_cry_6_THRU_CO ;
    wire \ppm_encoder_1.elevatorZ0Z_7 ;
    wire \ppm_encoder_1.un1_aileron_cry_12_THRU_CO ;
    wire \ppm_encoder_1.aileronZ0Z_13 ;
    wire \ppm_encoder_1.un1_elevator_cry_4_THRU_CO ;
    wire pid_altitude_dv;
    wire \ppm_encoder_1.elevatorZ0Z_5 ;
    wire \uart_drone.timer_Count_RNO_0_0_1 ;
    wire \uart_drone.timer_CountZ1Z_1 ;
    wire \uart_drone.N_144_1_cascade_ ;
    wire \uart_drone.N_145 ;
    wire \ppm_encoder_1.N_436 ;
    wire \ppm_encoder_1.N_508 ;
    wire \ppm_encoder_1.pulses2count_9_0_0_12 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_12 ;
    wire \ppm_encoder_1.pulses2count_9_0_3_12 ;
    wire \uart_drone.N_144_1 ;
    wire \uart_drone.N_143 ;
    wire \uart_drone.state_srsts_i_0_2_cascade_ ;
    wire \Commands_frame_decoder.stateZ0Z_11 ;
    wire \Commands_frame_decoder.state_RNIRSI31Z0Z_11 ;
    wire \uart_drone.stateZ0Z_2 ;
    wire \uart_drone.timer_Count_0_sqmuxa ;
    wire \uart_drone.timer_CountZ1Z_3 ;
    wire \uart_drone.un1_state_4_0 ;
    wire \uart_drone.stateZ0Z_1 ;
    wire \uart_drone_sync.aux_2__0__0_0 ;
    wire \uart_drone_sync.aux_3__0__0_0 ;
    wire \uart_drone.un1_state_2_0_a3_0 ;
    wire \reset_module_System.count_1_1_cascade_ ;
    wire \reset_module_System.reset6_19_cascade_ ;
    wire \reset_module_System.reset_isoZ0 ;
    wire \reset_module_System.reset6_13_cascade_ ;
    wire \reset_module_System.reset6_3 ;
    wire \reset_module_System.reset6_17 ;
    wire \reset_module_System.countZ0Z_0 ;
    wire \reset_module_System.countZ0Z_1 ;
    wire bfn_11_13_0_;
    wire \reset_module_System.count_1_cry_1 ;
    wire \reset_module_System.count_1_cry_2 ;
    wire \reset_module_System.countZ0Z_4 ;
    wire \reset_module_System.count_1_cry_3 ;
    wire \reset_module_System.countZ0Z_5 ;
    wire \reset_module_System.count_1_cry_4 ;
    wire \reset_module_System.count_1_cry_5 ;
    wire \reset_module_System.countZ0Z_7 ;
    wire \reset_module_System.count_1_cry_6 ;
    wire \reset_module_System.countZ0Z_8 ;
    wire \reset_module_System.count_1_cry_7 ;
    wire \reset_module_System.count_1_cry_8 ;
    wire \reset_module_System.countZ0Z_9 ;
    wire bfn_11_14_0_;
    wire \reset_module_System.countZ0Z_10 ;
    wire \reset_module_System.count_1_cry_9 ;
    wire \reset_module_System.countZ0Z_11 ;
    wire \reset_module_System.count_1_cry_10 ;
    wire \reset_module_System.countZ0Z_12 ;
    wire \reset_module_System.count_1_cry_11 ;
    wire \reset_module_System.count_1_cry_12 ;
    wire \reset_module_System.countZ0Z_14 ;
    wire \reset_module_System.count_1_cry_13 ;
    wire \reset_module_System.count_1_cry_14 ;
    wire \reset_module_System.countZ0Z_16 ;
    wire \reset_module_System.count_1_cry_15 ;
    wire \reset_module_System.count_1_cry_16 ;
    wire \reset_module_System.countZ0Z_17 ;
    wire bfn_11_15_0_;
    wire \reset_module_System.countZ0Z_18 ;
    wire \reset_module_System.count_1_cry_17 ;
    wire \reset_module_System.count_1_cry_18 ;
    wire \reset_module_System.count_1_cry_19 ;
    wire \reset_module_System.count_1_cry_20 ;
    wire \dron_frame_decoder_1.drone_H_disp_side_7 ;
    wire \Commands_frame_decoder.source_CH4data_1_sqmuxa ;
    wire \dron_frame_decoder_1.drone_H_disp_side_10 ;
    wire \dron_frame_decoder_1.drone_H_disp_side_8 ;
    wire \dron_frame_decoder_1.drone_H_disp_side_9 ;
    wire \dron_frame_decoder_1.N_716_0 ;
    wire debug_CH2_18A_c;
    wire \uart_pc.data_rdyc_1 ;
    wire \Commands_frame_decoder.stateZ0Z_6 ;
    wire alt_kp_4;
    wire \Commands_frame_decoder.stateZ0Z_7 ;
    wire xy_kp_4;
    wire \Commands_frame_decoder.un1_sink_data_valid_2_0 ;
    wire \Commands_frame_decoder.stateZ0Z_3 ;
    wire \Commands_frame_decoder.source_CH2data_1_sqmuxa ;
    wire \Commands_frame_decoder.stateZ0Z_4 ;
    wire \pid_alt.error_axbZ0Z_13 ;
    wire drone_altitude_13;
    wire \pid_alt.error_axbZ0Z_14 ;
    wire drone_altitude_14;
    wire \dron_frame_decoder_1.N_732_0 ;
    wire drone_altitude_2;
    wire \pid_alt.error_axbZ0Z_2 ;
    wire drone_altitude_3;
    wire \pid_alt.error_axbZ0Z_3 ;
    wire drone_H_disp_front_1;
    wire \dron_frame_decoder_1.drone_altitude_11 ;
    wire drone_altitude_i_11;
    wire \dron_frame_decoder_1.drone_H_disp_front_5 ;
    wire \dron_frame_decoder_1.drone_H_disp_front_6 ;
    wire bfn_11_22_0_;
    wire \pid_front.un11lto30_i_a2 ;
    wire \pid_front.un11lto30_i_a2_0 ;
    wire \pid_front.un11lto30_i_a2_1 ;
    wire \pid_front.un11lto30_i_a2_2 ;
    wire \pid_front.un11lto30_i_a2_3 ;
    wire \pid_front.un11lto30_i_a2_4 ;
    wire \pid_front.un11lto30_i_a2_5 ;
    wire \pid_front.un11lto30_i_a2_6 ;
    wire bfn_11_23_0_;
    wire \pid_front.un11lto30_i_a2_0_and ;
    wire \pid_front.un1_reset_i_a2_3_4_cascade_ ;
    wire \pid_front.N_593_cascade_ ;
    wire front_order_5;
    wire \pid_front.N_11_i ;
    wire \ppm_encoder_1.pulses2countZ0Z_14 ;
    wire \ppm_encoder_1.pulses2countZ0Z_15 ;
    wire \ppm_encoder_1.counter24_0_I_45_c_RNOZ0 ;
    wire \ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_a2_18_8_cascade_ ;
    wire \ppm_encoder_1.N_486_18 ;
    wire \ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_a2_18_10 ;
    wire \ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_a2_18_11 ;
    wire \ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_a2_18_9 ;
    wire \ppm_encoder_1.PPM_STATE_fast_RNICIABZ0Z_0 ;
    wire \ppm_encoder_1.counterZ0Z_0 ;
    wire bfn_12_2_0_;
    wire \ppm_encoder_1.counterZ0Z_1 ;
    wire \ppm_encoder_1.un1_counter_13_cry_0 ;
    wire \ppm_encoder_1.counterZ0Z_2 ;
    wire \ppm_encoder_1.un1_counter_13_cry_1 ;
    wire \ppm_encoder_1.counterZ0Z_3 ;
    wire \ppm_encoder_1.un1_counter_13_cry_2 ;
    wire \ppm_encoder_1.counterZ0Z_4 ;
    wire \ppm_encoder_1.un1_counter_13_cry_3 ;
    wire \ppm_encoder_1.counterZ0Z_5 ;
    wire \ppm_encoder_1.un1_counter_13_cry_4 ;
    wire \ppm_encoder_1.counterZ0Z_6 ;
    wire \ppm_encoder_1.un1_counter_13_cry_5 ;
    wire \ppm_encoder_1.counterZ0Z_7 ;
    wire \ppm_encoder_1.un1_counter_13_cry_6 ;
    wire \ppm_encoder_1.un1_counter_13_cry_7 ;
    wire \ppm_encoder_1.counterZ0Z_8 ;
    wire bfn_12_3_0_;
    wire \ppm_encoder_1.counterZ0Z_9 ;
    wire \ppm_encoder_1.un1_counter_13_cry_8 ;
    wire \ppm_encoder_1.counterZ0Z_10 ;
    wire \ppm_encoder_1.un1_counter_13_cry_9 ;
    wire \ppm_encoder_1.counterZ0Z_11 ;
    wire \ppm_encoder_1.un1_counter_13_cry_10 ;
    wire \ppm_encoder_1.counterZ0Z_12 ;
    wire \ppm_encoder_1.un1_counter_13_cry_11 ;
    wire \ppm_encoder_1.counterZ0Z_13 ;
    wire \ppm_encoder_1.un1_counter_13_cry_12 ;
    wire \ppm_encoder_1.counterZ0Z_14 ;
    wire \ppm_encoder_1.un1_counter_13_cry_13 ;
    wire \ppm_encoder_1.counterZ0Z_15 ;
    wire \ppm_encoder_1.un1_counter_13_cry_14 ;
    wire \ppm_encoder_1.un1_counter_13_cry_15 ;
    wire \ppm_encoder_1.counterZ0Z_16 ;
    wire bfn_12_4_0_;
    wire \ppm_encoder_1.counterZ0Z_17 ;
    wire \ppm_encoder_1.un1_counter_13_cry_16 ;
    wire \ppm_encoder_1.un1_counter_13_cry_17 ;
    wire \ppm_encoder_1.counterZ0Z_18 ;
    wire \ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83 ;
    wire side_order_12;
    wire side_order_13;
    wire \ppm_encoder_1.aileronZ0Z_14 ;
    wire \ppm_encoder_1.throttleZ0Z_14 ;
    wire \ppm_encoder_1.pulses2count_9_i_0_14_cascade_ ;
    wire \ppm_encoder_1.pulses2count_9_i_1_14 ;
    wire \ppm_encoder_1.un2_throttle_0_0_2_5 ;
    wire \ppm_encoder_1.pulses2count_9_i_0_5 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z2 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z2 ;
    wire \ppm_encoder_1.N_301_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_0_2_6 ;
    wire \ppm_encoder_1.pulses2count_9_0_0_6 ;
    wire \ppm_encoder_1.N_301 ;
    wire \ppm_encoder_1.pulses2count_9_i_1_7 ;
    wire side_order_10;
    wire side_order_11;
    wire side_order_6;
    wire side_order_7;
    wire side_order_8;
    wire side_order_9;
    wire \ppm_encoder_1.throttleZ0Z_7 ;
    wire \ppm_encoder_1.aileronZ0Z_7 ;
    wire \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ;
    wire \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ;
    wire \ppm_encoder_1.pulses2count_9_i_0_7 ;
    wire \uart_drone.stateZ0Z_3 ;
    wire \uart_drone.stateZ0Z_4 ;
    wire \uart_drone.timer_CountZ0Z_4 ;
    wire \uart_drone.state_srsts_0_0_0_cascade_ ;
    wire \uart_drone.N_126_li ;
    wire \uart_drone.stateZ0Z_0 ;
    wire \pid_side.error_i_acumm_13_0_a2_3_0_2 ;
    wire front_order_10;
    wire front_order_11;
    wire front_order_6;
    wire front_order_7;
    wire front_order_8;
    wire front_order_9;
    wire front_order_1;
    wire front_order_4;
    wire \reset_module_System.count_1_2 ;
    wire \reset_module_System.reset6_14 ;
    wire \reset_module_System.reset6_19 ;
    wire \reset_module_System.countZ0Z_6 ;
    wire \reset_module_System.countZ0Z_3 ;
    wire \reset_module_System.countZ0Z_20 ;
    wire \reset_module_System.countZ0Z_2 ;
    wire \reset_module_System.reset6_11 ;
    wire \pid_front.state_RNIVIRQZ0Z_0 ;
    wire uart_pc_data_rdy;
    wire \Commands_frame_decoder.un1_state57_iZ0 ;
    wire \pid_side.state_RNINK4UZ0Z_0_cascade_ ;
    wire \reset_module_System.countZ0Z_19 ;
    wire \reset_module_System.countZ0Z_15 ;
    wire \reset_module_System.countZ0Z_21 ;
    wire \reset_module_System.countZ0Z_13 ;
    wire \reset_module_System.reset6_15 ;
    wire \pid_front.m64_i_o2_0_cascade_ ;
    wire \pid_front.error_i_reg_esr_RNO_4_0_14_cascade_ ;
    wire \pid_front.m64_i_o2_0 ;
    wire \pid_front.m9_2_03_3_i_0_o2_0_1_cascade_ ;
    wire \pid_front.m9_2_03_3_i_0_o2_0_cascade_ ;
    wire drone_H_disp_front_3;
    wire drone_H_disp_front_2;
    wire \dron_frame_decoder_1.drone_H_disp_front_4 ;
    wire \pid_front.error_axb_0 ;
    wire bfn_12_18_0_;
    wire \pid_front.error_axbZ0Z_1 ;
    wire \pid_front.error_cry_0 ;
    wire \pid_front.error_axbZ0Z_2 ;
    wire \pid_front.error_cry_1 ;
    wire \pid_front.error_axbZ0Z_3 ;
    wire \pid_front.error_cry_2 ;
    wire drone_H_disp_front_i_4;
    wire \pid_front.error_cry_3 ;
    wire drone_H_disp_front_i_5;
    wire \pid_front.error_cry_0_0 ;
    wire drone_H_disp_front_i_6;
    wire \pid_front.error_cry_1_0 ;
    wire \pid_front.error_cry_2_0 ;
    wire \pid_front.error_cry_3_0 ;
    wire bfn_12_19_0_;
    wire \pid_front.error_cry_4 ;
    wire drone_H_disp_front_i_10;
    wire \pid_front.error_cry_5 ;
    wire \pid_front.error_cry_6 ;
    wire \pid_front.error_cry_7 ;
    wire \pid_front.error_cry_8 ;
    wire drone_H_disp_front_i_13;
    wire \pid_front.error_cry_9 ;
    wire \pid_front.error_cry_10 ;
    wire front_command_0;
    wire front_command_1;
    wire front_command_2;
    wire front_command_3;
    wire front_command_4;
    wire front_command_5;
    wire front_command_6;
    wire \Commands_frame_decoder.source_CH3data_1_sqmuxa_0 ;
    wire drone_H_disp_front_14;
    wire \dron_frame_decoder_1.drone_H_disp_front_10 ;
    wire \pid_front.un11lto30_i_a2_4_and ;
    wire \pid_front.N_175_cascade_ ;
    wire \pid_front.N_593 ;
    wire \pid_front.N_277_cascade_ ;
    wire \pid_front.N_291 ;
    wire \pid_front.un1_reset_i_o3_0_cascade_ ;
    wire \pid_front.N_342 ;
    wire \pid_front.un1_reset_0_i_3_cascade_ ;
    wire front_order_13;
    wire \pid_front.N_277 ;
    wire front_order_12;
    wire \pid_front.N_2364_i_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNIBG6FZ0Z_7 ;
    wire \pid_front.error_p_reg_esr_RNIGL6F_0Z0Z_8 ;
    wire \pid_front.error_p_reg_esr_RNIBG6FZ0Z_7_cascade_ ;
    wire \pid_front.error_d_reg_prevZ0Z_7 ;
    wire \pid_front.error_p_regZ0Z_8 ;
    wire \pid_front.error_p_reg_esr_RNIGL6FZ0Z_8_cascade_ ;
    wire \pid_front.un11lto30_i_a2_3_and ;
    wire \pid_front.un11lto30_i_a2_2_and ;
    wire \pid_front.pid_preregZ0Z_14 ;
    wire \pid_front.source_pid_9_i_0_o3_0_11 ;
    wire \pid_front.source_pid_9_i_0_o3_0_11_cascade_ ;
    wire \pid_front.N_175 ;
    wire \pid_front.un1_pid_prereg_0_9_cascade_ ;
    wire \pid_front.un1_pid_prereg_0_10_cascade_ ;
    wire \pid_front.un1_pid_prereg_0_8 ;
    wire \pid_front.un1_pid_prereg_0_8_cascade_ ;
    wire \pid_front.un1_pid_prereg_0_9 ;
    wire \pid_front.un11lto30_i_a2_5_and ;
    wire \pid_front.N_2364_i ;
    wire \pid_front.error_p_regZ0Z_7 ;
    wire \pid_front.error_p_reg_esr_RNIBG6F_0Z0Z_7_cascade_ ;
    wire \pid_front.un11lto30_i_a2_6_and ;
    wire \pid_front.error_d_reg_prev_esr_RNIQHN6Z0Z_1_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNI2BC9_0Z0Z_1_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNI2BC9Z0Z_1 ;
    wire \pid_front.O_0_10 ;
    wire \pid_side.error_i_acumm_13_i_o2_0_7_3_cascade_ ;
    wire \pid_side.un1_reset_i_a2_4_cascade_ ;
    wire \pid_side.N_342_cascade_ ;
    wire \pid_side.un1_reset_0_i_3_cascade_ ;
    wire side_order_1;
    wire side_order_2;
    wire side_order_3;
    wire \pid_side.state_0_0 ;
    wire \pid_side.source_pid_9_i_0_o3_0_11_cascade_ ;
    wire \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ;
    wire \ppm_encoder_1.N_267_i ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_12_1 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_2_12 ;
    wire \ppm_encoder_1.N_267_i_i ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_12_cascade_ ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_RNI1TA86Z0Z_2 ;
    wire \pid_side.N_531_cascade_ ;
    wire \pid_side.N_544_cascade_ ;
    wire \pid_side.N_603 ;
    wire \pid_side.N_181_cascade_ ;
    wire \pid_side.error_i_acumm_13_i_0_1_3_cascade_ ;
    wire \pid_side.error_i_acumm_13_i_0_3_cascade_ ;
    wire \pid_side.N_177 ;
    wire \pid_side.N_544 ;
    wire \pid_side.N_233_cascade_ ;
    wire \pid_side.N_251_cascade_ ;
    wire \uart_drone.bit_CountZ0Z_0 ;
    wire \uart_drone.bit_CountZ0Z_1 ;
    wire \uart_drone.bit_CountZ0Z_2 ;
    wire \uart_drone.data_Auxce_0_0_0 ;
    wire \uart_drone.data_Auxce_0_1 ;
    wire \uart_drone.data_Auxce_0_0_2 ;
    wire \uart_drone.data_Auxce_0_3 ;
    wire \uart_drone.data_Auxce_0_0_4 ;
    wire \uart_drone.data_Auxce_0_5 ;
    wire \uart_drone.data_Auxce_0_6 ;
    wire \uart_drone.un1_state_2_0 ;
    wire debug_CH0_16A_c;
    wire \uart_drone.N_152 ;
    wire \uart_drone.state_RNIOU0NZ0Z_4 ;
    wire \uart_drone.data_AuxZ0Z_0 ;
    wire \uart_drone.data_AuxZ0Z_1 ;
    wire \uart_drone.data_AuxZ0Z_2 ;
    wire \uart_drone.data_AuxZ0Z_3 ;
    wire \uart_drone.data_AuxZ0Z_4 ;
    wire \uart_drone.data_AuxZ0Z_5 ;
    wire \uart_drone.data_AuxZ0Z_6 ;
    wire \uart_drone.data_AuxZ0Z_7 ;
    wire \uart_drone.data_rdyc_1_0 ;
    wire \uart_drone.timer_Count_RNIES9Q1Z0Z_2 ;
    wire \pid_front.error_cry_2_c_RNIFP8GZ0Z1 ;
    wire \pid_front.m26_2_03_0_m2_ns_1_cascade_ ;
    wire \pid_front.m27_2_03_0_0_cascade_ ;
    wire \pid_front.N_253 ;
    wire \dron_frame_decoder_1.drone_H_disp_front_7 ;
    wire drone_H_disp_front_i_7;
    wire drone_H_disp_front_i_8;
    wire \dron_frame_decoder_1.drone_H_disp_front_9 ;
    wire drone_H_disp_front_i_9;
    wire uart_drone_data_1;
    wire drone_H_disp_side_1;
    wire uart_drone_data_2;
    wire drone_H_disp_side_2;
    wire drone_H_disp_side_3;
    wire \dron_frame_decoder_1.drone_H_disp_side_4 ;
    wire \dron_frame_decoder_1.drone_H_disp_side_5 ;
    wire uart_drone_data_6;
    wire \dron_frame_decoder_1.drone_H_disp_side_6 ;
    wire \dron_frame_decoder_1.N_724_0 ;
    wire \pid_side.error_i_reg_esr_RNO_6Z0Z_12_cascade_ ;
    wire dron_frame_decoder_1_source_H_disp_front_fast_0;
    wire \dron_frame_decoder_1.N_708_0 ;
    wire \pid_front.N_510_cascade_ ;
    wire \pid_front.N_596_cascade_ ;
    wire \pid_front.m9_2_03_3_i_0_o2_1 ;
    wire \pid_front.m9_2_03_3_i_3_cascade_ ;
    wire \pid_front.N_162_cascade_ ;
    wire uart_drone_data_3;
    wire uart_drone_data_4;
    wire uart_drone_data_5;
    wire drone_H_disp_front_13;
    wire uart_drone_data_7;
    wire drone_H_disp_front_15;
    wire uart_drone_data_0;
    wire \dron_frame_decoder_1.drone_H_disp_front_8 ;
    wire \dron_frame_decoder_1.N_700_0 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_21 ;
    wire \pid_alt.N_545 ;
    wire \pid_alt.error_i_acumm7lto13 ;
    wire \pid_alt.error_i_acummZ0Z_13 ;
    wire \pid_alt.N_72_i_0 ;
    wire \pid_alt.un1_reset_1_0_i ;
    wire \pid_front.error_axb_8_l_ofx_0 ;
    wire drone_H_disp_front_11;
    wire front_command_7;
    wire \pid_front.error_axbZ0Z_7 ;
    wire drone_H_disp_front_12;
    wire drone_H_disp_front_i_12;
    wire \pid_front.un1_reset_i_a2_5 ;
    wire \pid_front.source_pid10lt4_0 ;
    wire \pid_front.un1_reset_i_a2_4 ;
    wire \pid_front.state_RNIPKTDZ0Z_0 ;
    wire \pid_front.state_RNIPKTDZ0Z_0_cascade_ ;
    wire bfn_13_23_0_;
    wire \pid_front.un1_pid_prereg_0_cry_0_c_THRU_CO ;
    wire \pid_front.pid_preregZ0Z_1 ;
    wire \pid_front.un1_pid_prereg_0_cry_0 ;
    wire \pid_front.error_d_reg_prev_esr_RNID19M1Z0Z_1 ;
    wire \pid_front.un1_pid_prereg_0_cry_1 ;
    wire \pid_front.un1_pid_prereg_0_cry_2 ;
    wire \pid_front.pid_preregZ0Z_4 ;
    wire \pid_front.un1_pid_prereg_0_cry_3 ;
    wire \pid_front.pid_preregZ0Z_5 ;
    wire \pid_front.un1_pid_prereg_0_cry_4 ;
    wire \pid_front.pid_preregZ0Z_6 ;
    wire \pid_front.un1_pid_prereg_0_cry_5 ;
    wire \pid_front.un1_pid_prereg_0_cry_6 ;
    wire \pid_front.pid_preregZ0Z_7 ;
    wire bfn_13_24_0_;
    wire \pid_front.error_p_reg_esr_RNI3K9L1Z0Z_6 ;
    wire \pid_front.error_p_reg_esr_RNIS0F23Z0Z_7 ;
    wire \pid_front.pid_preregZ0Z_8 ;
    wire \pid_front.un1_pid_prereg_0_cry_7 ;
    wire \pid_front.error_p_reg_esr_RNIV7CQ2Z0Z_8 ;
    wire \pid_front.error_p_reg_esr_RNIPC5D1Z0Z_7 ;
    wire \pid_front.pid_preregZ0Z_9 ;
    wire \pid_front.un1_pid_prereg_0_cry_8 ;
    wire \pid_front.pid_preregZ0Z_10 ;
    wire \pid_front.un1_pid_prereg_0_cry_9 ;
    wire \pid_front.pid_preregZ0Z_11 ;
    wire \pid_front.un1_pid_prereg_0_cry_10 ;
    wire \pid_front.pid_preregZ0Z_12 ;
    wire \pid_front.un1_pid_prereg_0_cry_11 ;
    wire \pid_front.pid_preregZ0Z_13 ;
    wire \pid_front.un1_pid_prereg_0_cry_12 ;
    wire \pid_front.un1_pid_prereg_0_cry_13_THRU_CO ;
    wire \pid_front.un1_pid_prereg_0_cry_13 ;
    wire \pid_front.un1_pid_prereg_0_cry_14 ;
    wire \pid_front.pid_preregZ0Z_15 ;
    wire bfn_13_25_0_;
    wire \pid_front.pid_preregZ0Z_16 ;
    wire \pid_front.un1_pid_prereg_0_cry_15 ;
    wire \pid_front.pid_preregZ0Z_17 ;
    wire \pid_front.un1_pid_prereg_0_cry_16 ;
    wire \pid_front.pid_preregZ0Z_18 ;
    wire \pid_front.un1_pid_prereg_0_cry_17 ;
    wire \pid_front.pid_preregZ0Z_19 ;
    wire \pid_front.un1_pid_prereg_0_cry_18 ;
    wire \pid_front.error_p_reg_esr_RNI80EDDZ0Z_17 ;
    wire \pid_front.pid_preregZ0Z_20 ;
    wire \pid_front.un1_pid_prereg_0_cry_19 ;
    wire \pid_front.error_p_reg_esr_RNIRNJEDZ0Z_18 ;
    wire \pid_front.error_p_reg_esr_RNIQOPM6Z0Z_18 ;
    wire \pid_front.pid_preregZ0Z_21 ;
    wire \pid_front.un1_pid_prereg_0_cry_20 ;
    wire \pid_front.error_p_reg_esr_RNI1VPN6Z0Z_19 ;
    wire \pid_front.pid_preregZ0Z_22 ;
    wire \pid_front.un1_pid_prereg_0_cry_21 ;
    wire \pid_front.un1_pid_prereg_0_cry_22 ;
    wire \pid_front.pid_preregZ0Z_23 ;
    wire bfn_13_26_0_;
    wire \pid_front.pid_preregZ0Z_24 ;
    wire \pid_front.un1_pid_prereg_0_cry_23 ;
    wire \pid_front.pid_preregZ0Z_25 ;
    wire \pid_front.un1_pid_prereg_0_cry_24 ;
    wire \pid_front.pid_preregZ0Z_26 ;
    wire \pid_front.un1_pid_prereg_0_cry_25 ;
    wire \pid_front.pid_preregZ0Z_27 ;
    wire \pid_front.un1_pid_prereg_0_cry_26 ;
    wire \pid_front.pid_preregZ0Z_28 ;
    wire \pid_front.un1_pid_prereg_0_cry_27 ;
    wire \pid_front.pid_preregZ0Z_29 ;
    wire \pid_front.un1_pid_prereg_0_cry_28 ;
    wire \pid_front.un1_pid_prereg_0_cry_29 ;
    wire \pid_front.pid_preregZ0Z_30 ;
    wire \pid_front.N_2358_i_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNI6B6FZ0Z_6 ;
    wire \pid_front.error_p_reg_esr_RNIBG6F_0Z0Z_7 ;
    wire \pid_front.error_p_reg_esr_RNI6B6FZ0Z_6_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNI3K9L1_0Z0Z_6 ;
    wire \pid_front.error_p_reg_esr_RNIMVC9Z0Z_6_cascade_ ;
    wire \pid_front.error_d_reg_prevZ0Z_6 ;
    wire \pid_front.O_0_5 ;
    wire \pid_front.error_p_regZ0Z_1 ;
    wire \pid_front.un1_pid_prereg_9_0_cascade_ ;
    wire \pid_front.error_d_reg_prev_esr_RNIMRLTZ0Z_0 ;
    wire \pid_front.O_4 ;
    wire \pid_front.error_d_reg_prevZ0Z_0 ;
    wire \pid_front.error_d_reg_prev_esr_RNIAHDKZ0Z_0 ;
    wire \pid_front.N_5_0 ;
    wire \pid_front.error_p_reg_esr_RNI6D5L7Z0Z_12_cascade_ ;
    wire \pid_front.un1_pid_prereg_0_axb_14 ;
    wire \pid_front.O_3 ;
    wire \pid_front.error_d_regZ0Z_0 ;
    wire bfn_14_3_0_;
    wire \pid_side.un11lto30_i_a2_0_and ;
    wire \pid_side.un11lto30_i_a2 ;
    wire \pid_side.un11lto30_i_a2_0 ;
    wire \pid_side.un11lto30_i_a2_2_and ;
    wire \pid_side.un11lto30_i_a2_1 ;
    wire \pid_side.un11lto30_i_a2_2 ;
    wire \pid_side.un11lto30_i_a2_3 ;
    wire \pid_side.un11lto30_i_a2_4 ;
    wire \pid_side.un11lto30_i_a2_5 ;
    wire \pid_side.un11lto30_i_a2_6 ;
    wire \pid_side.source_pid_9_i_0_o3_0_11 ;
    wire bfn_14_4_0_;
    wire \pid_side.un1_reset_i_a2_5 ;
    wire \pid_side.N_291 ;
    wire \pid_side.un1_reset_i_o3_0 ;
    wire \pid_side.N_631_cascade_ ;
    wire side_order_4;
    wire \pid_side.un1_reset_i_a2_3_4_cascade_ ;
    wire \pid_side.N_593 ;
    wire \pid_side.N_593_cascade_ ;
    wire side_order_5;
    wire \pid_side.N_11_i ;
    wire \pid_side.N_386 ;
    wire \pid_side.N_631 ;
    wire side_order_0;
    wire \pid_side.state_0_1 ;
    wire \pid_side.un1_reset_0_i_3 ;
    wire \pid_side.N_251 ;
    wire \pid_side.error_i_acumm16lto3 ;
    wire \pid_side.error_i_acumm_preregZ0Z_5 ;
    wire \pid_side.error_i_acumm_preregZ0Z_6 ;
    wire \pid_side.error_i_acumm_preregZ0Z_4 ;
    wire \pid_side.error_i_acumm_13_0_a2_2_2_2_cascade_ ;
    wire \pid_side.N_255 ;
    wire \pid_side.error_i_acumm_13_i_0_tz_7 ;
    wire \pid_side.error_i_acumm_preregZ0Z_1 ;
    wire \pid_side.N_181 ;
    wire \pid_side.N_483_cascade_ ;
    wire \pid_side.error_i_acumm_13_0_a2_2_4_2 ;
    wire \pid_side.error_i_acumm_preregZ0Z_9 ;
    wire \pid_side.error_i_acumm_preregZ0Z_8 ;
    wire \pid_side.N_217 ;
    wire \pid_side.error_i_acumm_preregZ0Z_7 ;
    wire \pid_side.N_488_cascade_ ;
    wire \pid_side.N_601 ;
    wire \pid_side.N_601_cascade_ ;
    wire \pid_side.error_i_acumm_preregZ0Z_0 ;
    wire \pid_side.N_484_cascade_ ;
    wire \pid_side.N_484 ;
    wire \pid_side.error_i_acumm_preregZ0Z_2 ;
    wire \pid_side.error_i_acumm_13_0_tz_0_0 ;
    wire \pid_side.N_634 ;
    wire \pid_side.error_i_acumm_preregZ0Z_10 ;
    wire \pid_side.N_355_cascade_ ;
    wire \pid_side.N_242_cascade_ ;
    wire \pid_side.un10lto12 ;
    wire \pid_side.N_227 ;
    wire \pid_side.N_205 ;
    wire \pid_side.N_285 ;
    wire \pid_side.N_353_cascade_ ;
    wire \pid_side.error_i_acumm_preregZ0Z_11 ;
    wire \pid_front.pid_preregZ0Z_0 ;
    wire front_order_0;
    wire \pid_front.pid_preregZ0Z_2 ;
    wire front_order_2;
    wire \pid_front.N_386 ;
    wire \pid_front.N_631 ;
    wire \pid_front.pid_preregZ0Z_3 ;
    wire front_order_3;
    wire \pid_front.state_0_1 ;
    wire \pid_front.un1_reset_0_i_3 ;
    wire \pid_side.error_d_reg_prev_esr_RNI5RIOZ0Z_14_cascade_ ;
    wire \pid_side.un1_pid_prereg_0_20_cascade_ ;
    wire \pid_side.un1_pid_prereg_0_22_cascade_ ;
    wire \pid_side.un1_pid_prereg_0_20 ;
    wire \pid_side.un1_pid_prereg_0_21 ;
    wire \pid_side.error_i_acumm_preregZ0Z_13 ;
    wire \pid_side.error_i_acumm_13_i_o2_0_10_3 ;
    wire \pid_side.error_i_acumm_preregZ0Z_18 ;
    wire \pid_side.error_i_acumm_preregZ0Z_25 ;
    wire \pid_side.error_i_acumm_preregZ0Z_26 ;
    wire \pid_side.N_338 ;
    wire pid_side_N_382_4_cascade_;
    wire \pid_side.N_382_cascade_ ;
    wire \pid_side.N_64 ;
    wire \pid_side.state_RNIL5IFZ0Z_0_cascade_ ;
    wire \pid_side.state_RNIIIOOZ0Z_0 ;
    wire \pid_side.stateZ0Z_0 ;
    wire \pid_side.stateZ0Z_1 ;
    wire \pid_front.state_ns_0_cascade_ ;
    wire \pid_front.N_536_1 ;
    wire \pid_front.N_297 ;
    wire \pid_front.O_0_22 ;
    wire \pid_front.O_0_8 ;
    wire \pid_front.O_7 ;
    wire drone_H_disp_side_11;
    wire \pid_front.N_581_cascade_ ;
    wire \pid_front.error_i_reg_esr_RNO_0Z0Z_10_cascade_ ;
    wire \pid_front.N_581 ;
    wire \pid_front.error_cry_1_0_c_RNII2EF1Z0Z_0_cascade_ ;
    wire \pid_front.N_228 ;
    wire \pid_front.N_228_cascade_ ;
    wire \pid_front.error_i_reg_9_sn_26 ;
    wire \pid_front.error_cry_1_0_c_RNII2EFZ0Z1 ;
    wire \pid_front.N_182_cascade_ ;
    wire \pid_front.N_597_cascade_ ;
    wire \pid_front.m12_2_03_4_i_0_cascade_ ;
    wire \pid_front.N_583 ;
    wire \pid_front.N_583_cascade_ ;
    wire \pid_front.N_597 ;
    wire \pid_front.error_i_reg_esr_RNO_0Z0Z_8_cascade_ ;
    wire \pid_front.N_598 ;
    wire \pid_front.m28_2_03_0 ;
    wire \pid_front.m28_2_03_0_0 ;
    wire \pid_front.N_302_cascade_ ;
    wire \pid_front.error_i_reg_9_rn_2_25_cascade_ ;
    wire \pid_front.error_i_reg_9_sn_25 ;
    wire \pid_front.m9_2_03_3_i_3 ;
    wire \pid_front.m27_2_03_0 ;
    wire \pid_front.N_154 ;
    wire \pid_front.N_225_cascade_ ;
    wire \pid_front.N_478_cascade_ ;
    wire \pid_front.error_i_reg_9_N_5L8_0_1_cascade_ ;
    wire \pid_front.error_i_reg_esr_RNO_0Z0Z_21 ;
    wire \pid_front.N_45_i_i_0_cascade_ ;
    wire \pid_front.error_cry_1_0_c_RNINF5AZ0Z3_cascade_ ;
    wire \pid_front.un4_error_i_reg_28_ns_1_1_cascade_ ;
    wire \pid_front.error_i_reg_9_1_18 ;
    wire \pid_front.un4_error_i_reg_28_ns_1_cascade_ ;
    wire \pid_front.m6_2_01 ;
    wire \pid_front.un1_pid_prereg_0_11 ;
    wire \pid_front.un1_pid_prereg_0_12_cascade_ ;
    wire \pid_front.un1_pid_prereg_0_10 ;
    wire \pid_front.error_d_reg_prev_esr_RNIV42ACZ0Z_21 ;
    wire \pid_front.error_d_reg_prev_esr_RNIU58I5Z0Z_21 ;
    wire \pid_front.un1_pid_prereg_0_12 ;
    wire \pid_front.un1_pid_prereg_0_14_cascade_ ;
    wire \pid_front.error_d_reg_prev_esr_RNION3U9Z0Z_21 ;
    wire \pid_front.un1_pid_prereg_0_13 ;
    wire \pid_front.un1_pid_prereg_0_15_cascade_ ;
    wire \pid_front.error_d_reg_prev_esr_RNIQHRB4Z0Z_21 ;
    wire \pid_front.error_p_reg_esr_RNID8DF2Z0Z_3 ;
    wire \pid_front.error_p_reg_esr_RNIR7E8Z0Z_3 ;
    wire \pid_front.error_p_reg_esr_RNIR7E8Z0Z_3_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNIRJAF2Z0Z_3 ;
    wire \pid_front.error_p_regZ0Z_4 ;
    wire \pid_front.error_p_reg_esr_RNIUAE8_0Z0Z_4 ;
    wire \pid_front.error_p_reg_esr_RNIPKK71Z0Z_2 ;
    wire \pid_front.error_p_regZ0Z_3 ;
    wire \pid_front.error_d_reg_prevZ0Z_3 ;
    wire \pid_front.error_p_reg_esr_RNIR7E8_0Z0Z_3 ;
    wire \pid_front.error_p_reg_esr_RNIR7E8_0Z0Z_3_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNIQ7CF2Z0Z_2 ;
    wire \pid_front.error_d_reg_prevZ0Z_1 ;
    wire \pid_front.error_d_regZ0Z_1 ;
    wire \pid_front.error_d_reg_prev_esr_RNIFSHOZ0Z_1 ;
    wire \pid_front.error_d_reg_prev_esr_RNI1JN71Z0Z_1 ;
    wire \pid_alt.state_0_0 ;
    wire \pid_front.error_d_reg_prev_esr_RNI1K4E5Z0Z_10 ;
    wire \pid_front.N_2370_i ;
    wire \pid_front.error_p_reg_esr_RNIB9N71Z0Z_5 ;
    wire \pid_front.un1_pid_prereg_0_1_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNIUFCM6Z0Z_14 ;
    wire \pid_front.un1_pid_prereg_0_2_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNICIRCDZ0Z_14 ;
    wire \pid_front.un1_pid_prereg_0_0 ;
    wire \pid_front.un1_pid_prereg_0_1 ;
    wire \pid_front.un1_pid_prereg_0_0_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNIA6C3NZ0Z_14 ;
    wire \pid_front.error_d_reg_prev_esr_RNIQ9AEDZ0Z_10 ;
    wire \pid_front.un1_pid_prereg_0_17_cascade_ ;
    wire \pid_front.error_d_reg_prev_esr_RNIUNTB4Z0Z_21 ;
    wire \pid_front.un1_pid_prereg_0_18_cascade_ ;
    wire \pid_front.error_d_reg_prev_esr_RNI0MTN8Z0Z_21 ;
    wire \pid_front.un1_pid_prereg_0_14 ;
    wire \pid_front.un1_pid_prereg_0_15 ;
    wire \pid_front.un1_pid_prereg_0_17 ;
    wire \pid_front.error_d_reg_prev_esr_RNIO9PN8Z0Z_21 ;
    wire \pid_front.error_p_reg_esr_RNIE2FM6Z0Z_15 ;
    wire \pid_front.un1_pid_prereg_0_19_cascade_ ;
    wire \pid_front.error_d_reg_prev_esr_RNI2UVB4Z0Z_21 ;
    wire \pid_front.error_p_regZ0Z_6 ;
    wire \pid_front.error_p_reg_esr_RNIMVC9_0Z0Z_6 ;
    wire \pid_front.error_p_reg_esr_RNIJ26O1Z0Z_5 ;
    wire \pid_front.error_d_reg_prev_esr_RNISAJOZ0Z_6 ;
    wire \pid_front.un1_pid_prereg_66_0_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNIUBTV2Z0Z_5 ;
    wire \pid_front.error_p_reg_esr_RNIVOSGZ0Z_5 ;
    wire \pid_front.error_d_reg_prevZ0Z_5 ;
    wire \pid_front.error_p_reg_esr_RNIUAE8Z0Z_4 ;
    wire \pid_front.error_p_regZ0Z_5 ;
    wire \pid_front.error_p_reg_esr_RNIVOSG_0Z0Z_5 ;
    wire \pid_front.error_p_reg_esr_RNIVOSG_0Z0Z_5_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNIB9N71_0Z0Z_5 ;
    wire \pid_front.un1_pid_prereg_0_20_cascade_ ;
    wire \pid_front.error_d_reg_prev_esr_RNI642C4Z0Z_21 ;
    wire \pid_front.un1_pid_prereg_0_22_cascade_ ;
    wire \pid_front.error_d_reg_prev_esr_RNIGE6O8Z0Z_21 ;
    wire \pid_front.un1_pid_prereg_0_18 ;
    wire \pid_front.un1_pid_prereg_0_19 ;
    wire \pid_front.un1_pid_prereg_0_20 ;
    wire \pid_front.error_d_reg_prev_esr_RNI822O8Z0Z_21 ;
    wire \pid_front.un1_pid_prereg_0_23_cascade_ ;
    wire \pid_front.error_d_reg_prev_esr_RNIAA4C4Z0Z_21 ;
    wire \pid_front.un1_pid_prereg_0_21 ;
    wire \pid_side.error_i_acumm_preregZ0Z_14 ;
    wire \pid_side.error_i_acumm_13_i_o2_0_10_12 ;
    wire \pid_side.error_i_acumm_13_i_o2_0_8_12 ;
    wire \pid_side.error_i_acumm_13_i_o2_0_9_12_cascade_ ;
    wire \pid_side.error_i_acumm_13_i_o2_0_7_12 ;
    wire \pid_side.N_203 ;
    wire \pid_side.error_i_acumm_preregZ0Z_22 ;
    wire \pid_side.error_i_acumm_preregZ0Z_27 ;
    wire \pid_side.error_i_acumm_13_i_o2_0_8_3 ;
    wire \pid_side.error_i_acumm_preregZ0Z_19 ;
    wire \pid_side.error_i_acumm_preregZ0Z_20 ;
    wire \pid_side.error_i_acumm_preregZ0Z_21 ;
    wire \pid_side.error_i_acumm_preregZ0Z_23 ;
    wire \pid_side.error_i_acumm_preregZ0Z_17 ;
    wire \pid_side.error_i_acumm_13_i_o2_0_9_3 ;
    wire \pid_side.error_i_acumm_preregZ0Z_15 ;
    wire \pid_side.error_i_acumm_preregZ0Z_16 ;
    wire \pid_side.un11lto30_i_a2_5_and ;
    wire \pid_side.un11lto30_i_a2_5_and_cascade_ ;
    wire \pid_side.N_175 ;
    wire \pid_side.N_175_cascade_ ;
    wire \pid_side.pid_preregZ0Z_14 ;
    wire \pid_side.N_277 ;
    wire \pid_side.un11lto30_i_a2_6_and ;
    wire \pid_side.un11lto30_i_a2_3_and ;
    wire \pid_side.un11lto30_i_a2_4_and ;
    wire \pid_side.un1_pid_prereg_0_1_cascade_ ;
    wire \pid_side.un1_pid_prereg_0_2_cascade_ ;
    wire \pid_side.un1_pid_prereg_0_3_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNI5RIOZ0Z_14 ;
    wire \pid_side.un1_pid_prereg_0_0 ;
    wire \pid_side.un1_pid_prereg_0_0_cascade_ ;
    wire \pid_side.un1_pid_prereg_0_1 ;
    wire \pid_side.error_d_reg_prev_esr_RNIB1JOZ0Z_16 ;
    wire \pid_side.error_d_reg_prev_esr_RNIB1JOZ0Z_16_cascade_ ;
    wire \pid_side.un1_pid_prereg_0_2 ;
    wire \pid_side.un1_pid_prereg_0_3 ;
    wire \pid_side.un1_pid_prereg_0_4_cascade_ ;
    wire \pid_side.error_d_reg_prevZ0Z_16 ;
    wire \pid_side.error_d_reg_prev_esr_RNIB1JO_0Z0Z_16 ;
    wire \pid_side.error_d_reg_prev_esr_RNIE4JO_0Z0Z_17 ;
    wire \pid_side.un1_pid_prereg_0_5_cascade_ ;
    wire \pid_side.error_i_acummZ0Z_0 ;
    wire bfn_15_8_0_;
    wire \pid_side.error_i_acummZ0Z_1 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_0 ;
    wire \pid_side.error_i_acummZ0Z_2 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_1 ;
    wire \pid_side.error_i_regZ0Z_3 ;
    wire \pid_side.error_i_acummZ0Z_3 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_2 ;
    wire \pid_side.error_i_acummZ0Z_4 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_3 ;
    wire \pid_side.error_i_acummZ0Z_5 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_4 ;
    wire \pid_side.error_i_acummZ0Z_6 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_5 ;
    wire \pid_side.error_i_acummZ0Z_7 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_6 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_7 ;
    wire \pid_side.error_i_acummZ0Z_8 ;
    wire bfn_15_9_0_;
    wire \pid_side.error_i_acummZ0Z_9 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_8 ;
    wire \pid_side.error_i_acummZ0Z_10 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_9 ;
    wire \pid_side.error_i_acummZ0Z_11 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_10 ;
    wire \pid_side.error_i_acummZ0Z_12 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_11 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_12 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_13 ;
    wire \pid_side.error_i_reg_esr_RNIQ9ORZ0Z_15 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_14 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_15 ;
    wire \pid_side.error_i_reg_esr_RNISCPRZ0Z_16 ;
    wire bfn_15_10_0_;
    wire \pid_side.error_i_reg_esr_RNIUFQRZ0Z_17 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_16 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_17 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_18 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_19 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_20 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_21 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_22 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_23 ;
    wire bfn_15_11_0_;
    wire \pid_side.un1_error_i_acumm_prereg_cry_24 ;
    wire \pid_side.error_i_reg_esr_RNIUHTSZ0Z_26 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_25 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_26 ;
    wire \pid_side.error_i_acummZ0Z_13 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_27 ;
    wire \pid_side.error_i_acumm_preregZ0Z_28 ;
    wire \pid_side.error_i_acumm_preregZ0Z_24 ;
    wire \pid_side.error_i_regZ0Z_1 ;
    wire \pid_side.N_302_cascade_ ;
    wire \pid_side.error_i_regZ0Z_25 ;
    wire \pid_side.error_i_reg_9_rn_0_27_cascade_ ;
    wire \pid_side.N_42_i_i_0 ;
    wire \pid_side.error_i_regZ0Z_27 ;
    wire \pid_side.error_i_regZ0Z_14 ;
    wire \pid_front.error_i_reg_esr_RNO_5Z0Z_21 ;
    wire pid_side_N_174_cascade_;
    wire \pid_front.error_i_reg_esr_RNO_4Z0Z_21 ;
    wire pid_side_N_495_cascade_;
    wire \pid_side.m4_2_01_cascade_ ;
    wire \pid_side.error_i_regZ0Z_0 ;
    wire \pid_side.m4_2_01_1 ;
    wire \pid_side.m64_i_o2_0_cascade_ ;
    wire \pid_side.error_cry_1_c_RNI6K4BZ0Z1_cascade_ ;
    wire \pid_side.N_111 ;
    wire \pid_front.N_161_cascade_ ;
    wire \pid_front.N_398 ;
    wire \pid_front.m78_0_0 ;
    wire \pid_front.m78_0_1_cascade_ ;
    wire \pid_front.N_626 ;
    wire \pid_front.N_626_cascade_ ;
    wire \pid_front.error_i_reg_esr_RNO_0Z0Z_6_cascade_ ;
    wire \pid_front.N_232 ;
    wire \pid_front.m10_2_03_3_i_0_o2_0 ;
    wire \pid_front.N_207 ;
    wire \pid_front.N_556 ;
    wire \pid_front.m10_2_03_3_i_0_o2_0_cascade_ ;
    wire \pid_front.m10_2_03_3_i_3_cascade_ ;
    wire \pid_front.N_301 ;
    wire \pid_front.N_510 ;
    wire \pid_front.N_554_cascade_ ;
    wire \pid_front.N_543 ;
    wire pid_side_m13_2_03_4_i_0_a2_3_0;
    wire \pid_front.m13_2_03_4_i_0_o2_2 ;
    wire \pid_front.m13_2_03_4_i_0_o2_2_cascade_ ;
    wire \pid_front.error_i_reg_esr_RNO_0Z0Z_9_cascade_ ;
    wire \pid_front.m13_2_03_4_i_0_o2_1 ;
    wire \pid_front.N_184_cascade_ ;
    wire \pid_front.N_576 ;
    wire \pid_front.N_575_cascade_ ;
    wire \pid_front.N_229 ;
    wire \pid_front.m11_2_03_3_i_3 ;
    wire \pid_front.m11_2_03_3_i_3_cascade_ ;
    wire \pid_front.un1_pid_prereg_0 ;
    wire bfn_15_19_0_;
    wire \pid_front.un1_error_i_acumm_prereg_cry_0 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_1 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_2 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_3 ;
    wire \pid_front.error_i_regZ0Z_5 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_4 ;
    wire \pid_front.error_i_regZ0Z_6 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_5 ;
    wire \pid_front.error_i_regZ0Z_7 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_6 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_7 ;
    wire \pid_front.error_i_regZ0Z_8 ;
    wire bfn_15_20_0_;
    wire \pid_front.error_i_regZ0Z_9 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_8 ;
    wire \pid_front.error_i_regZ0Z_10 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_9 ;
    wire \pid_front.error_i_regZ0Z_11 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_10 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_11 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_12 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_13 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_14 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_15 ;
    wire bfn_15_21_0_;
    wire \pid_front.un1_error_i_acumm_prereg_cry_16 ;
    wire \pid_front.error_i_regZ0Z_18 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_17 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_18 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_19 ;
    wire \pid_front.error_i_regZ0Z_21 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_20 ;
    wire \pid_front.error_i_regZ0Z_22 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_21 ;
    wire \pid_front.error_i_regZ0Z_23 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_22 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_23 ;
    wire \pid_front.error_i_regZ0Z_24 ;
    wire bfn_15_22_0_;
    wire \pid_front.error_i_regZ0Z_25 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_24 ;
    wire \pid_front.error_i_regZ0Z_26 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_25 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_26 ;
    wire \pid_front.error_i_acummZ0Z_13 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_27 ;
    wire \pid_front.error_p_reg_esr_RNIO4E8_0Z0Z_2 ;
    wire \pid_front.error_p_regZ0Z_2 ;
    wire \pid_front.error_d_reg_prevZ0Z_2 ;
    wire \pid_front.error_p_reg_esr_RNIO4E8Z0Z_2 ;
    wire \pid_front.error_p_regZ0Z_17 ;
    wire \pid_front.error_d_reg_prevZ0Z_17 ;
    wire \pid_front.error_p_reg_esr_RNIKG5U_0Z0Z_10_cascade_ ;
    wire \pid_front.error_d_reg_prev_esr_RNI379B2Z0Z_10_cascade_ ;
    wire \pid_front.error_d_reg_prev_esr_RNI5JRF4_0Z0Z_10 ;
    wire \pid_front.error_p_reg_esr_RNIKG5UZ0Z_10 ;
    wire \pid_front.un1_pid_prereg_153_0 ;
    wire \pid_front.un1_pid_prereg_0_16 ;
    wire \pid_front.error_d_reg_prev_esr_RNI379B2Z0Z_10 ;
    wire \pid_front.error_d_reg_prev_esr_RNI5JRF4Z0Z_10 ;
    wire \pid_front.error_d_reg_prev_esr_RNI5JRF4Z0Z_10_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNIEU1SDZ0Z_12 ;
    wire \pid_front.error_p_reg_esr_RNIUKHM6Z0Z_16 ;
    wire \pid_front.un1_pid_prereg_0_6_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNICS5DDZ0Z_16 ;
    wire \pid_front.error_p_reg_esr_RNIQ9C61_0Z0Z_17 ;
    wire \pid_front.error_p_reg_esr_RNIN6C61Z0Z_16 ;
    wire \pid_front.un1_pid_prereg_0_4 ;
    wire \pid_front.un1_pid_prereg_0_2 ;
    wire \pid_front.un1_pid_prereg_0_3 ;
    wire \pid_front.un1_pid_prereg_0_4_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNICN0DDZ0Z_15 ;
    wire \pid_front.error_p_regZ0Z_16 ;
    wire \pid_front.error_p_reg_esr_RNIN6C61_0Z0Z_16 ;
    wire \pid_front.error_d_reg_prevZ0Z_16 ;
    wire \pid_front.error_i_acumm_preregZ0Z_13 ;
    wire \pid_front.error_i_acumm_preregZ0Z_18 ;
    wire \pid_front.error_i_reg_esr_RNI8KHVZ0Z_25 ;
    wire \pid_front.error_i_acumm_preregZ0Z_25 ;
    wire \pid_front.error_i_reg_esr_RNIANIVZ0Z_26 ;
    wire \pid_front.error_i_acumm_preregZ0Z_26 ;
    wire \pid_front.error_d_reg_prev_esr_RNIL8SR5Z0Z_12 ;
    wire \pid_front.error_p_reg_esr_RNITCC61_0Z0Z_18 ;
    wire \pid_front.error_p_reg_esr_RNIQ9C61Z0Z_17 ;
    wire \pid_front.error_i_reg_esr_RNICOGUZ0Z_18 ;
    wire \pid_front.un1_pid_prereg_0_5 ;
    wire \pid_front.O_16 ;
    wire \pid_front.O_0_17 ;
    wire \pid_front.error_d_reg_prev_esr_RNI8QE61_0Z0Z_20 ;
    wire \pid_front.error_d_reg_prev_esr_RNI8QE61Z0Z_20 ;
    wire \pid_front.O_0_24 ;
    wire \pid_front.error_d_reg_fast_esr_RNISQ181Z0Z_12_cascade_ ;
    wire \pid_front.error_d_reg_esr_RNIETB61_3Z0Z_13 ;
    wire \pid_front.g1_2_1 ;
    wire \pid_front.g0_3_2_cascade_ ;
    wire \pid_front.error_i_reg_esr_RNI29BUZ0Z_13 ;
    wire \pid_front.g1_3_cascade_ ;
    wire \pid_front.error_d_regZ0Z_13 ;
    wire \pid_front.N_2401_0_cascade_ ;
    wire \pid_front.g0_2 ;
    wire \pid_side.source_pid10lt4_0 ;
    wire bfn_16_4_0_;
    wire \pid_side.pid_preregZ0Z_0 ;
    wire \pid_side.un1_pid_prereg_0_cry_0_c_THRU_CO ;
    wire \pid_side.pid_preregZ0Z_1 ;
    wire \pid_side.un1_pid_prereg_0_cry_0 ;
    wire \pid_side.pid_preregZ0Z_2 ;
    wire \pid_side.un1_pid_prereg_0_cry_1 ;
    wire \pid_side.pid_preregZ0Z_3 ;
    wire \pid_side.un1_pid_prereg_0_cry_2 ;
    wire \pid_side.pid_preregZ0Z_4 ;
    wire \pid_side.un1_pid_prereg_0_cry_3 ;
    wire \pid_side.pid_preregZ0Z_5 ;
    wire \pid_side.un1_pid_prereg_0_cry_4 ;
    wire \pid_side.pid_preregZ0Z_6 ;
    wire \pid_side.un1_pid_prereg_0_cry_5 ;
    wire \pid_side.un1_pid_prereg_0_cry_6 ;
    wire \pid_side.pid_preregZ0Z_7 ;
    wire bfn_16_5_0_;
    wire \pid_side.pid_preregZ0Z_8 ;
    wire \pid_side.un1_pid_prereg_0_cry_7 ;
    wire \pid_side.pid_preregZ0Z_9 ;
    wire \pid_side.un1_pid_prereg_0_cry_8 ;
    wire \pid_side.pid_preregZ0Z_10 ;
    wire \pid_side.un1_pid_prereg_0_cry_9 ;
    wire \pid_side.pid_preregZ0Z_11 ;
    wire \pid_side.un1_pid_prereg_0_cry_10 ;
    wire \pid_side.pid_preregZ0Z_12 ;
    wire \pid_side.un1_pid_prereg_0_cry_11 ;
    wire \pid_side.pid_preregZ0Z_13 ;
    wire \pid_side.un1_pid_prereg_0_cry_12 ;
    wire \pid_side.un1_pid_prereg_0_cry_13_THRU_CO ;
    wire \pid_side.un1_pid_prereg_0_cry_13 ;
    wire \pid_side.un1_pid_prereg_0_cry_14 ;
    wire \pid_side.pid_preregZ0Z_15 ;
    wire bfn_16_6_0_;
    wire \pid_side.error_d_reg_prev_esr_RNI2SL2GZ0Z_12 ;
    wire \pid_side.pid_preregZ0Z_16 ;
    wire \pid_side.un1_pid_prereg_0_cry_15 ;
    wire \pid_side.error_d_reg_prev_esr_RNISHTJ9Z0Z_14 ;
    wire \pid_side.error_d_reg_prev_esr_RNIMFTP4Z0Z_14 ;
    wire \pid_side.pid_preregZ0Z_17 ;
    wire \pid_side.un1_pid_prereg_0_cry_16 ;
    wire \pid_side.error_d_reg_prev_esr_RNISM2K9Z0Z_15 ;
    wire \pid_side.error_d_reg_prev_esr_RNI620Q4Z0Z_15 ;
    wire \pid_side.pid_preregZ0Z_18 ;
    wire \pid_side.un1_pid_prereg_0_cry_17 ;
    wire \pid_side.error_d_reg_prev_esr_RNIMK2Q4Z0Z_16 ;
    wire \pid_side.pid_preregZ0Z_19 ;
    wire \pid_side.un1_pid_prereg_0_cry_18 ;
    wire \pid_side.pid_preregZ0Z_20 ;
    wire \pid_side.un1_pid_prereg_0_cry_19 ;
    wire \pid_side.pid_preregZ0Z_21 ;
    wire \pid_side.un1_pid_prereg_0_cry_20 ;
    wire \pid_side.pid_preregZ0Z_22 ;
    wire \pid_side.un1_pid_prereg_0_cry_21 ;
    wire \pid_side.un1_pid_prereg_0_cry_22 ;
    wire \pid_side.pid_preregZ0Z_23 ;
    wire bfn_16_7_0_;
    wire \pid_side.pid_preregZ0Z_24 ;
    wire \pid_side.un1_pid_prereg_0_cry_23 ;
    wire \pid_side.pid_preregZ0Z_25 ;
    wire \pid_side.un1_pid_prereg_0_cry_24 ;
    wire \pid_side.error_d_reg_prev_esr_RNI8N8M6Z0Z_21 ;
    wire \pid_side.pid_preregZ0Z_26 ;
    wire \pid_side.un1_pid_prereg_0_cry_25 ;
    wire \pid_side.error_d_reg_prev_esr_RNIG3DM6Z0Z_21 ;
    wire \pid_side.error_d_reg_prev_esr_RNIME5B3Z0Z_21 ;
    wire \pid_side.pid_preregZ0Z_27 ;
    wire \pid_side.un1_pid_prereg_0_cry_26 ;
    wire \pid_side.error_d_reg_prev_esr_RNIQK7B3Z0Z_21 ;
    wire \pid_side.pid_preregZ0Z_28 ;
    wire \pid_side.un1_pid_prereg_0_cry_27 ;
    wire \pid_side.pid_preregZ0Z_29 ;
    wire \pid_side.un1_pid_prereg_0_cry_28 ;
    wire \pid_side.un1_pid_prereg_0_cry_29 ;
    wire \pid_side.pid_preregZ0Z_30 ;
    wire \pid_side.state_0_g_0 ;
    wire \pid_side.error_d_reg_prev_esr_RNIC7HE7Z0Z_21 ;
    wire \pid_side.un1_pid_prereg_0_11_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNIPUAR4Z0Z_19 ;
    wire \pid_side.error_d_reg_prev_esr_RNIE21B3Z0Z_21 ;
    wire \pid_side.un1_pid_prereg_0_15_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNIASUA3Z0Z_21 ;
    wire \pid_side.error_i_reg_esr_RNIK2OSZ0Z_21 ;
    wire \pid_side.un1_pid_prereg_370_1 ;
    wire \pid_side.error_i_reg_esr_RNIRGURZ0Z_20 ;
    wire \pid_side.un1_pid_prereg_0_9_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNIIOAQ4Z0Z_18 ;
    wire \pid_side.error_i_reg_esr_RNI0JRRZ0Z_18 ;
    wire \pid_side.error_i_reg_esr_RNI2MSRZ0Z_19 ;
    wire \pid_side.un1_pid_prereg_0_7_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNI675Q4Z0Z_17 ;
    wire \pid_side.N_3_i_1_1_cascade_ ;
    wire \pid_side.N_5 ;
    wire \pid_side.N_3_i_1_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNIQTGL4Z0Z_12_cascade_ ;
    wire \pid_side.un1_pid_prereg_0_axb_14 ;
    wire \pid_side.N_5_0 ;
    wire \pid_side.un1_pid_prereg_79_cascade_ ;
    wire \pid_side.N_543 ;
    wire CONSTANT_ONE_NET;
    wire \pid_side.m13_2_03_4_i_0_o2_1_cascade_ ;
    wire \pid_side.m13_2_03_4_i_3 ;
    wire \pid_side.m13_2_03_4_i_3_cascade_ ;
    wire \pid_side.error_i_regZ0Z_9 ;
    wire \pid_side.state_ns_0 ;
    wire \pid_side.error_i_regZ0Z_7 ;
    wire \pid_side.N_163 ;
    wire \pid_side.N_163_cascade_ ;
    wire \pid_side.N_186_cascade_ ;
    wire \pid_side.error_i_reg_9_sn_27 ;
    wire \pid_front.N_394 ;
    wire \pid_front.error_i_reg_9_rn_1_26 ;
    wire pid_side_m10_2_03_3_i_0_a2_1_0_cascade_;
    wire \pid_side.m13_2_03_4_i_0_o2_1_0_cascade_ ;
    wire \pid_side.error_cry_3_0_c_RNIER8NCZ0 ;
    wire \pid_side.m18_2_03_4_o3_1_cascade_ ;
    wire \pid_side.N_263_cascade_ ;
    wire \pid_side.error_i_reg_esr_RNO_1Z0Z_14 ;
    wire \pid_side.m18_2_03_4_o3_1_1 ;
    wire \pid_front.N_629 ;
    wire \pid_side.N_228_0 ;
    wire \pid_side.m16_2_03_4_0_cascade_ ;
    wire \pid_side.N_263 ;
    wire \pid_side.N_189_cascade_ ;
    wire \pid_side.m5_0_03_4_i_i_0 ;
    wire \pid_side.N_6 ;
    wire \pid_side.N_6_cascade_ ;
    wire \pid_side.error_i_reg_esr_RNO_2Z0Z_16_cascade_ ;
    wire \pid_side.error_i_regZ0Z_16 ;
    wire \pid_side.m4_2_01 ;
    wire \pid_side.error_i_reg_esr_RNO_1Z0Z_16 ;
    wire \pid_side.N_259 ;
    wire \pid_side.N_259_cascade_ ;
    wire \pid_side.error_i_reg_esr_RNO_2Z0Z_14 ;
    wire \pid_front.N_156 ;
    wire \pid_front.N_163_cascade_ ;
    wire \pid_front.N_186 ;
    wire \pid_front.N_186_cascade_ ;
    wire \pid_front.N_338 ;
    wire \pid_front.N_339 ;
    wire \pid_front.N_42_i_i_0_cascade_ ;
    wire \pid_front.error_i_reg_9_sn_27 ;
    wire \pid_front.error_i_regZ0Z_27 ;
    wire \pid_front.error_i_reg_9_rn_0_27 ;
    wire \pid_front.N_458 ;
    wire \pid_front.N_314_cascade_ ;
    wire \pid_front.N_225 ;
    wire \pid_front.m24_2_03_0_0_cascade_ ;
    wire \pid_front.m24_2_03_0_1 ;
    wire \pid_front.m24_2_03_0_cascade_ ;
    wire \pid_front.error_i_regZ0Z_20 ;
    wire \pid_front.error_i_regZ0Z_0 ;
    wire \pid_front.error_cry_1_c_RNILQ1FZ0Z2 ;
    wire pid_side_N_607_cascade_;
    wire \pid_front.error_cry_1_0_c_RNINF5AZ0Z3 ;
    wire \pid_front.error_i_regZ0Z_2 ;
    wire \pid_front.error_i_regZ0Z_1 ;
    wire pid_front_N_335_cascade_;
    wire \pid_side.error_i_reg_9_1_rn_sx_16_cascade_ ;
    wire \pid_side.error_i_reg_9_1_sn_16 ;
    wire \pid_side.error_i_reg_9_1_rn_0_16_cascade_ ;
    wire \pid_side.error_i_reg_9_1_16 ;
    wire \pid_front.N_600_cascade_ ;
    wire \pid_front.error_i_acumm_preregZ0Z_0 ;
    wire \pid_front.error_i_acumm_13_0_tz_1_0_cascade_ ;
    wire \pid_front.error_i_acummZ0Z_0 ;
    wire \pid_front.error_i_acummZ0Z_1 ;
    wire \pid_front.error_i_acumm_13_0_tz_1_0 ;
    wire \pid_front.error_i_acummZ0Z_2 ;
    wire \pid_front.error_i_acummZ0Z_6 ;
    wire \pid_front.error_i_acummZ0Z_5 ;
    wire \pid_front.N_633_cascade_ ;
    wire \pid_front.N_530 ;
    wire \pid_front.N_251 ;
    wire \pid_front.N_251_cascade_ ;
    wire \pid_front.error_i_acummZ0Z_4 ;
    wire \pid_front.error_i_acummZ0Z_7 ;
    wire \pid_front.error_i_acummZ0Z_8 ;
    wire \pid_front.N_62_i_1_cascade_ ;
    wire \pid_front.error_i_acummZ0Z_3 ;
    wire \pid_front.N_177 ;
    wire \pid_front.N_177_cascade_ ;
    wire \pid_front.N_158_cascade_ ;
    wire \pid_front.N_601 ;
    wire \pid_front.N_208 ;
    wire \pid_front.N_181 ;
    wire \pid_front.N_483 ;
    wire \pid_front.un1_pid_prereg_0_25_cascade_ ;
    wire \pid_front.error_d_reg_prev_esr_RNIDF6C4Z0Z_21 ;
    wire \pid_front.un1_pid_prereg_0_axb_30 ;
    wire \pid_front.error_d_reg_prev_esr_RNIR0EO8Z0Z_21 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_27_c_RNIDSKV ;
    wire \pid_front.un1_pid_prereg_0_26 ;
    wire \pid_front.un1_pid_prereg_0_24 ;
    wire \pid_front.un1_pid_prereg_0_23 ;
    wire \pid_front.un1_pid_prereg_0_22 ;
    wire \pid_front.un1_pid_prereg_0_24_cascade_ ;
    wire \pid_front.un1_pid_prereg_0_25 ;
    wire \pid_front.error_d_reg_prev_esr_RNINPAO8Z0Z_21 ;
    wire \pid_front.error_p_regZ0Z_20 ;
    wire \pid_front.un1_pid_prereg_370_1 ;
    wire \pid_front.error_d_reg_prevZ0Z_20 ;
    wire \pid_front.error_d_reg_prevZ0Z_21 ;
    wire \pid_front.error_d_regZ0Z_4 ;
    wire \pid_front.error_d_reg_prevZ0Z_4 ;
    wire \pid_front.error_p_reg_esr_RNIGL6FZ0Z_8 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_8_c_RNI1BPE ;
    wire \pid_front.g0_1_0 ;
    wire \pid_front.error_p_reg_esr_RNI8NB61_1Z0Z_11 ;
    wire \pid_front.error_d_reg_prevZ0Z_15 ;
    wire \pid_front.error_p_reg_esr_RNIK3C61Z0Z_15 ;
    wire \pid_front.error_d_reg_fast_esr_RNI5VGKZ0Z_12 ;
    wire \pid_front.error_d_reg_fast_esr_RNID6KB1Z0Z_12_cascade_ ;
    wire \pid_front.error_d_reg_fast_esr_RNIQSG63Z0Z_12_cascade_ ;
    wire \pid_front.error_d_reg_esr_RNIETB61Z0Z_13 ;
    wire \pid_front.error_p_reg_esr_RNIH0C61_0Z0Z_14 ;
    wire \pid_front.error_p_reg_esr_RNIK42C6Z0Z_14_cascade_ ;
    wire \pid_front.un1_pid_prereg_167_0_1_cascade_ ;
    wire \pid_front.un1_pid_prereg_167_0 ;
    wire \pid_front.error_d_reg_fast_esr_RNIR9PO_0Z0Z_13 ;
    wire \pid_front.error_d_reg_fast_esr_RNIQSG63Z0Z_12 ;
    wire \pid_front.error_d_reg_prev_esr_RNIJVGT4Z0Z_12 ;
    wire \pid_front.error_p_reg_esr_RNILTVH2Z0Z_12 ;
    wire \pid_front.N_2394_i ;
    wire \pid_front.N_3_i_1_1_cascade_ ;
    wire \pid_front.N_3_i_1 ;
    wire \pid_front.un1_pid_prereg_79 ;
    wire \pid_front.un1_pid_prereg_135_0 ;
    wire \pid_front.error_d_reg_prev_fastZ0Z_12 ;
    wire \pid_front.O_0_4 ;
    wire \pid_front.error_p_regZ0Z_0 ;
    wire \pid_front.O_0_14 ;
    wire \pid_front.O_0_15 ;
    wire \pid_front.O_0_16 ;
    wire \pid_front.O_0_18 ;
    wire \pid_front.O_0_19 ;
    wire \pid_front.error_p_regZ0Z_15 ;
    wire \pid_front.error_p_regZ0Z_13 ;
    wire \pid_front.error_d_reg_prevZ0Z_13 ;
    wire \pid_front.error_d_reg_fastZ0Z_13 ;
    wire \pid_front.error_p_regZ0Z_14 ;
    wire \pid_front.error_d_reg_prevZ0Z_14 ;
    wire \pid_front.N_2401_0_0_0_cascade_ ;
    wire \pid_front.N_4_1_1_1 ;
    wire \pid_front.g0_2_0_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNIBIFG6Z0Z_12 ;
    wire \pid_side.error_d_reg_prev_esr_RNISKLO_0Z0Z_20 ;
    wire \pid_side.error_d_reg_prevZ0Z_20 ;
    wire \pid_side.error_d_reg_prev_esr_RNISKLOZ0Z_20 ;
    wire \pid_side.error_d_reg_prev_esr_RNIOUJE2Z0Z_6_cascade_ ;
    wire \pid_side.un1_pid_prereg_66_0_cascade_ ;
    wire \pid_side.error_p_reg_esr_RNIRH187Z0Z_5 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_5_c_RNIC5QN ;
    wire \pid_side.error_d_reg_prev_esr_RNIOUJE2Z0Z_6 ;
    wire \pid_side.error_p_reg_esr_RNIBABR4Z0Z_5 ;
    wire \pid_side.error_d_reg_prev_esr_RNI8UIO_0Z0Z_15 ;
    wire \pid_side.error_d_reg_prevZ0Z_15 ;
    wire \pid_side.error_d_reg_prev_esr_RNI8UIOZ0Z_15 ;
    wire \pid_side.error_d_reg_prev_esr_RNIE4JOZ0Z_17 ;
    wire \pid_side.error_d_reg_prevZ0Z_17 ;
    wire \pid_side.error_d_reg_prev_esr_RNIGI4KKZ0Z_12 ;
    wire \pid_side.error_d_reg_prev_esr_RNI73UC2_0Z0Z_14 ;
    wire \pid_side.error_d_reg_prev_esr_RNICCO8BZ0Z_12 ;
    wire \pid_side.error_d_reg_prev_esr_RNIBNLL9Z0Z_18 ;
    wire \pid_side.error_d_reg_prev_esr_RNI2BI34Z0Z_21 ;
    wire \pid_side.error_i_reg_esr_RNIM5PSZ0Z_22 ;
    wire \pid_side.un1_pid_prereg_0_13 ;
    wire \pid_side.un1_pid_prereg_0_10 ;
    wire \pid_side.un1_pid_prereg_0_11 ;
    wire \pid_side.un1_pid_prereg_0_13_cascade_ ;
    wire \pid_side.un1_pid_prereg_0_12 ;
    wire \pid_side.error_d_reg_prev_esr_RNIR9TU8Z0Z_21 ;
    wire \pid_side.un1_pid_prereg_0_axb_30 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_26_c_RNI0LUS ;
    wire \pid_side.un1_pid_prereg_0_22 ;
    wire \pid_side.un1_pid_prereg_0_24_cascade_ ;
    wire \pid_side.un1_pid_prereg_0_23 ;
    wire \pid_side.error_d_reg_prev_esr_RNINEHM6Z0Z_21 ;
    wire \pid_side.error_d_reg_prev_esr_RNIRLKM6Z0Z_21 ;
    wire \pid_side.un1_pid_prereg_0_15 ;
    wire \pid_side.un1_pid_prereg_0_14 ;
    wire \pid_side.un1_pid_prereg_0_17_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNIOUVL6Z0Z_21 ;
    wire \pid_side.error_i_reg_esr_RNIO8QSZ0Z_23 ;
    wire \pid_side.un1_pid_prereg_0_4 ;
    wire \pid_side.un1_pid_prereg_0_5 ;
    wire \pid_side.error_d_reg_prev_esr_RNISR7K9Z0Z_16 ;
    wire \pid_side.error_i_reg_esr_RNIQBRSZ0Z_24 ;
    wire \pid_side.un1_pid_prereg_0_17 ;
    wire \pid_side.un1_pid_prereg_0_16 ;
    wire \pid_side.un1_pid_prereg_0_18_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNI0B4M6Z0Z_21 ;
    wire \pid_side.un1_pid_prereg_0_7 ;
    wire \pid_side.un1_pid_prereg_0_9 ;
    wire \pid_side.un1_pid_prereg_0_6 ;
    wire \pid_side.un1_pid_prereg_0_8 ;
    wire \pid_side.error_d_reg_prev_esr_RNIOVFK9Z0Z_17 ;
    wire \pid_side.un1_pid_prereg_0_18 ;
    wire \pid_side.error_d_reg_prev_esr_RNII83B3Z0Z_21 ;
    wire \pid_side.error_p_reg_esr_RNI4O091_0Z0Z_10_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNIV62K2Z0Z_10_cascade_ ;
    wire \pid_side.error_p_reg_esr_RNI4O091Z0Z_10 ;
    wire \pid_side.un1_pid_prereg_153_0_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNII28CBZ0Z_10 ;
    wire \pid_side.error_d_reg_prev_esr_RNIV62K2Z0Z_10 ;
    wire \pid_side.error_d_reg_prev_esr_RNID3GT3Z0Z_10 ;
    wire \pid_side.error_i_reg_esr_RNIJVKRZ0Z_12 ;
    wire \pid_side.error_d_reg_prev_esr_RNI9LLC4Z0Z_12 ;
    wire \pid_side.error_d_reg_prev_esr_RNID3GT3Z0Z_10_cascade_ ;
    wire \pid_side.error_p_reg_esr_RNIL0VP1Z0Z_12 ;
    wire \pid_side.error_d_reg_prev_esr_RNIUOPVAZ0Z_10 ;
    wire \pid_side.un1_pid_prereg_167_0_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNI59QR8Z0Z_12 ;
    wire \pid_side.un1_pid_prereg_167_0_1 ;
    wire \pid_side.un1_pid_prereg_79 ;
    wire \pid_side.error_d_reg_fast_esr_RNIPEC11Z0Z_12_cascade_ ;
    wire \pid_side.error_d_reg_fast_esr_RNIEIJH2Z0Z_12_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNIJHVG3Z0Z_12 ;
    wire \pid_side.error_d_reg_fast_esr_RNIPHKNZ0Z_12 ;
    wire \pid_side.error_d_reg_esr_RNI2OIOZ0Z_13 ;
    wire \pid_side.error_d_reg_fast_esr_RNIFGGE_0Z0Z_13 ;
    wire \pid_side.error_d_reg_prev_esr_RNI5RIO_0Z0Z_14 ;
    wire \pid_side.error_d_reg_fast_esr_RNIEIJH2Z0Z_12 ;
    wire \pid_side.error_d_reg_prev_esr_RNI4M9H4Z0Z_14 ;
    wire xy_ki_5;
    wire pid_side_N_490_cascade_;
    wire \pid_side.m78_0_a2_sx_cascade_ ;
    wire \pid_side.N_394 ;
    wire pid_side_m78_0_a2_0_0;
    wire \pid_side.m78_0_1 ;
    wire \pid_side.m78_0_0_cascade_ ;
    wire \pid_side.error_i_regZ0Z_11 ;
    wire \pid_side.N_626 ;
    wire \pid_side.N_626_cascade_ ;
    wire \pid_side.N_398 ;
    wire \pid_side.N_161_cascade_ ;
    wire \pid_side.m13_2_03_4_i_0_o2_2_1 ;
    wire \pid_side.N_594 ;
    wire \pid_side.N_594_cascade_ ;
    wire \pid_side.error_i_reg_9_sn_13_cascade_ ;
    wire \pid_side.error_i_regZ0Z_13 ;
    wire \pid_side.error_i_reg_esr_RNO_1_0_17 ;
    wire \pid_side.error_i_regZ0Z_17 ;
    wire \pid_side.m16_2_03_4 ;
    wire \pid_side.m0_2_03_cascade_ ;
    wire \pid_side.error_i_regZ0Z_12 ;
    wire \pid_side.m1_0_03_cascade_ ;
    wire \pid_side.error_i_reg_9_rn_1_13 ;
    wire \pid_side.N_232_cascade_ ;
    wire \pid_side.N_549_cascade_ ;
    wire \pid_side.error_i_reg_esr_RNO_0_0_6_cascade_ ;
    wire \pid_side.error_i_regZ0Z_6 ;
    wire \pid_side.N_580 ;
    wire \pid_side.N_156_cascade_ ;
    wire \pid_side.N_182 ;
    wire pid_side_m10_2_03_3_i_0_a2_1_0;
    wire \pid_side.N_549 ;
    wire \pid_side.N_182_cascade_ ;
    wire \Commands_frame_decoder.source_CH3data_1_sqmuxa ;
    wire \Commands_frame_decoder.N_403 ;
    wire \Commands_frame_decoder.stateZ0Z_5 ;
    wire \dron_frame_decoder_1.state_RNI6P6KZ0Z_4 ;
    wire \dron_frame_decoder_1.N_218 ;
    wire \dron_frame_decoder_1.stateZ0Z_7 ;
    wire debug_CH1_0A_c;
    wire \pid_alt.stateZ0Z_0 ;
    wire \pid_alt.N_72_i ;
    wire \pid_front.error_p_reg_esr_RNICMVCGZ0Z_14 ;
    wire \pid_side.N_2601_i ;
    wire \pid_front.N_429 ;
    wire \pid_front.N_332_cascade_ ;
    wire \pid_front.N_262 ;
    wire \pid_front.error_i_reg_esr_RNO_0Z0Z_17_cascade_ ;
    wire \pid_front.error_i_regZ0Z_17 ;
    wire \pid_front.N_6 ;
    wire \pid_front.m1_0_03 ;
    wire \pid_front.error_i_reg_esr_RNO_1Z0Z_17 ;
    wire \pid_front.m16_2_03_4_0_cascade_ ;
    wire \pid_front.m16_2_03_4_cascade_ ;
    wire \pid_front.error_i_regZ0Z_12 ;
    wire \pid_front.m18_2_03_4_1_cascade_ ;
    wire \pid_front.error_i_regZ0Z_14 ;
    wire \pid_front.N_580 ;
    wire \pid_front.N_187 ;
    wire \pid_front.N_263 ;
    wire \pid_front.N_54_i_1 ;
    wire \pid_front.N_54_i_1_cascade_ ;
    wire \pid_front.error_i_reg_esr_RNO_5Z0Z_16_cascade_ ;
    wire \pid_front.error_i_reg_9_rn_0_16_cascade_ ;
    wire \pid_front.error_i_regZ0Z_16 ;
    wire \pid_front.error_i_reg_9_sn_16 ;
    wire \pid_front.N_188 ;
    wire \pid_front.N_259 ;
    wire \pid_front.N_259_cascade_ ;
    wire \pid_front.N_111 ;
    wire \pid_front.error_i_reg_9_1_14 ;
    wire \pid_front.N_454 ;
    wire \pid_front.N_515_cascade_ ;
    wire \pid_front.N_450_cascade_ ;
    wire \pid_front.N_446_cascade_ ;
    wire \pid_front.m20_2_03_0_2 ;
    wire \pid_front.N_515 ;
    wire \pid_front.N_438_cascade_ ;
    wire \pid_front.error_i_reg_esr_RNI4CCUZ0Z_14 ;
    wire \pid_front.error_i_acumm_preregZ0Z_14 ;
    wire \pid_front.error_i_reg_esr_RNI2BEVZ0Z_22 ;
    wire \pid_front.error_i_acumm_preregZ0Z_22 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_26_c_RNICQJV ;
    wire \pid_front.error_i_acumm_preregZ0Z_27 ;
    wire \pid_front.N_439 ;
    wire \pid_side.N_109 ;
    wire \pid_front.error_d_reg_prevZ0Z_19 ;
    wire \pid_front.error_p_regZ0Z_19 ;
    wire \pid_front.error_p_reg_esr_RNI0GC61Z0Z_19 ;
    wire \pid_front.N_531_cascade_ ;
    wire \pid_front.N_255 ;
    wire \pid_front.error_i_acumm_preregZ0Z_9 ;
    wire \pid_front.N_633 ;
    wire \pid_front.N_255_cascade_ ;
    wire \pid_front.error_i_acummZ0Z_9 ;
    wire \pid_front.N_276 ;
    wire \pid_front.N_276_cascade_ ;
    wire \pid_front.N_632 ;
    wire pid_side_N_382_4;
    wire xy_ki_7;
    wire xy_ki_6;
    wire reset_system;
    wire \pid_front.stateZ0Z_0 ;
    wire \pid_front.N_382_cascade_ ;
    wire \pid_front.stateZ0Z_1 ;
    wire \pid_front.N_217 ;
    wire \pid_front.error_p_regZ0Z_10 ;
    wire \pid_front.N_2382_i_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNIFM3D1Z0Z_10_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNI6R6D1Z0Z_8 ;
    wire \pid_front.error_p_reg_esr_RNIS5CU3Z0Z_9 ;
    wire \pid_front.error_p_reg_esr_RNILQ6FZ0Z_9 ;
    wire \pid_front.error_d_reg_prev_esr_RNI1K4E5_0Z0Z_10 ;
    wire \pid_front.error_p_reg_esr_RNIFM3D1Z0Z_10 ;
    wire \pid_front.error_p_reg_esr_RNINU9V7Z0Z_9 ;
    wire \pid_front.error_d_reg_prevZ0Z_10 ;
    wire \pid_front.error_d_reg_prevZ0Z_9 ;
    wire \pid_front.N_2376_i ;
    wire \pid_front.error_d_reg_prevZ0Z_8 ;
    wire \pid_front.error_p_regZ0Z_9 ;
    wire \pid_front.N_2376_i_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNILQ6F_0Z0Z_9 ;
    wire \pid_front.error_i_acumm_preregZ0Z_15 ;
    wire \pid_front.error_i_reg_esr_RNI8IEUZ0Z_16 ;
    wire \pid_front.error_i_acumm_preregZ0Z_16 ;
    wire \pid_front.error_i_reg_esr_RNIALFUZ0Z_17 ;
    wire \pid_front.error_i_acumm_preregZ0Z_17 ;
    wire \pid_front.error_i_reg_esr_RNI6HGVZ0Z_24 ;
    wire \pid_front.error_i_acumm_preregZ0Z_24 ;
    wire \pid_front.error_p_reg_esr_RNIK3C61_0Z0Z_15 ;
    wire \pid_front.error_p_reg_esr_RNIH0C61Z0Z_14 ;
    wire \pid_front.error_i_reg_esr_RNI6FDUZ0Z_15 ;
    wire \pid_front.error_p_reg_esr_RNIBJ5B3_0Z0Z_14 ;
    wire \pid_front.error_p_reg_esr_RNIOH2JDZ0Z_12 ;
    wire \pid_front.error_p_reg_esr_RNIBJ5B3_0Z0Z_14_cascade_ ;
    wire \pid_front.error_d_reg_prev_esr_RNI13Q1DZ0Z_12 ;
    wire \pid_front.error_p_reg_esr_RNI4820UZ0Z_12 ;
    wire \pid_front.error_i_acumm_13_i_o2_0_9_3 ;
    wire \pid_front.error_i_acumm_13_i_o2_0_10_3 ;
    wire \pid_front.error_i_acumm_13_i_o2_0_7_3 ;
    wire \pid_front.error_i_acumm_13_i_o2_0_9_12 ;
    wire \pid_front.error_i_acumm_13_i_o2_0_10_12 ;
    wire \pid_front.error_i_acumm_13_i_o2_0_7_12 ;
    wire \pid_front.error_i_acumm_13_i_o2_0_8_12 ;
    wire \pid_front.error_i_acumm_preregZ0Z_19 ;
    wire \pid_front.error_i_acumm_13_i_o2_0_8_3 ;
    wire \pid_front.error_i_reg_esr_RNI7MJUZ0Z_20 ;
    wire \pid_front.error_i_acumm_preregZ0Z_20 ;
    wire \pid_front.error_i_reg_esr_RNI08DVZ0Z_21 ;
    wire \pid_front.error_i_acumm_preregZ0Z_21 ;
    wire \pid_front.error_i_reg_esr_RNI4EFVZ0Z_23 ;
    wire \pid_front.error_i_acumm_preregZ0Z_23 ;
    wire \pid_front.error_p_reg_esr_RNI0GC61_0Z0Z_19 ;
    wire \pid_front.error_i_reg_esr_RNIERHUZ0Z_19 ;
    wire \pid_front.un1_pid_prereg_0_7 ;
    wire \pid_front.un1_pid_prereg_0_7_cascade_ ;
    wire \pid_front.un1_pid_prereg_0_6 ;
    wire \pid_front.error_p_reg_esr_RNIE7KM6Z0Z_17 ;
    wire \pid_front.error_d_reg_fastZ0Z_12 ;
    wire \pid_front.error_p_regZ0Z_11 ;
    wire \pid_front.g0_1_0_1_cascade_ ;
    wire \pid_front.error_p_regZ0Z_12 ;
    wire \pid_front.g0_1 ;
    wire \pid_front.N_5 ;
    wire \pid_front.error_d_reg_prevZ0Z_11 ;
    wire \pid_front.N_763_0 ;
    wire \pid_front.state_RNIM14NZ0Z_0 ;
    wire \pid_side.N_2565_i_cascade_ ;
    wire \pid_side.error_p_reg_esr_RNINKTC1_0Z0Z_7 ;
    wire \pid_side.error_p_reg_esr_RNIIFTC1Z0Z_6 ;
    wire \pid_side.error_p_reg_esr_RNINKTC1_0Z0Z_7_cascade_ ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_6_c_RNI6FLJ ;
    wire \pid_side.error_p_reg_esr_RNIFJGD3_0Z0Z_6 ;
    wire \pid_side.error_d_reg_prevZ0Z_6 ;
    wire \pid_side.error_p_reg_esr_RNINKTC1Z0Z_7 ;
    wire \pid_side.error_p_reg_esr_RNIFJGD3Z0Z_6 ;
    wire \pid_side.error_p_reg_esr_RNINKTC1Z0Z_7_cascade_ ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_7_c_RNIIDSN ;
    wire \pid_side.error_p_reg_esr_RNIKF8V6Z0Z_7 ;
    wire \pid_side.error_i_regZ0Z_8 ;
    wire \pid_side.error_p_reg_esr_RNI5SNH3Z0Z_7 ;
    wire \pid_side.error_p_reg_esr_RNISPTC1Z0Z_8_cascade_ ;
    wire \pid_side.error_p_reg_esr_RNIECBV6Z0Z_8 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_8_c_RNICNNJ ;
    wire \pid_side.error_p_reg_esr_RNISPTC1Z0Z_8 ;
    wire \pid_side.error_p_reg_esr_RNI1VTC1_0Z0Z_9 ;
    wire \pid_side.N_2577_i ;
    wire \pid_side.N_2577_i_cascade_ ;
    wire \pid_side.error_p_reg_esr_RNISPTC1_0Z0Z_8 ;
    wire \pid_side.un1_pid_prereg_9_0_cascade_ ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_0_c_RNITGKN ;
    wire \pid_side.error_d_reg_prev_esr_RNIM6H42Z0Z_0 ;
    wire \pid_side.un1_pid_prereg_0_25 ;
    wire \pid_side.un1_pid_prereg_0_25_cascade_ ;
    wire \pid_side.un1_pid_prereg_0_24 ;
    wire \pid_side.error_d_reg_prev_esr_RNITP9B3Z0Z_21 ;
    wire \pid_side.un1_pid_prereg_0 ;
    wire \pid_side.error_d_reg_prev_esr_RNIHEJ01Z0Z_0 ;
    wire \pid_side.error_i_reg_esr_RNISESSZ0Z_25 ;
    wire \pid_side.un1_pid_prereg_0_19 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_27_c_RNI1NVS ;
    wire \pid_side.un1_pid_prereg_0_26 ;
    wire \pid_side.error_i_reg_esr_RNIGRJRZ0Z_11 ;
    wire \pid_side.error_d_reg_prev_esr_RNID3GT3_0Z0Z_10 ;
    wire \pid_side.error_d_reg_prev_esr_RNITU3P4Z0Z_10 ;
    wire \pid_side.N_2571_i ;
    wire \pid_side.error_d_reg_prevZ0Z_7 ;
    wire \pid_side.state_RNIL5IFZ0Z_0 ;
    wire \pid_side.error_d_reg_prevZ0Z_21 ;
    wire \pid_side.error_d_reg_prevZ0Z_8 ;
    wire \pid_side.error_p_reg_esr_RNI9GJD3Z0Z_8 ;
    wire \pid_side.error_p_reg_esr_RNI1VTC1Z0Z_9_cascade_ ;
    wire \pid_side.error_p_reg_esr_RNIBMBO6Z0Z_10 ;
    wire \pid_side.N_2589_i_cascade_ ;
    wire \pid_side.N_2583_i ;
    wire \pid_side.error_p_reg_esr_RNI1VTC1Z0Z_9 ;
    wire \pid_side.error_i_reg_esr_RNI6OOIZ0Z_10 ;
    wire \pid_side.error_d_reg_prev_esr_RNITU3P4_0Z0Z_10 ;
    wire \pid_side.error_p_reg_esr_RNIRE1B1Z0Z_10 ;
    wire \pid_side.error_p_reg_esr_RNIV4S38Z0Z_10 ;
    wire \pid_side.error_d_reg_prevZ0Z_9 ;
    wire \pid_side.error_d_reg_prevZ0Z_10 ;
    wire \pid_side.O_1_13 ;
    wire \pid_side.error_d_regZ0Z_10 ;
    wire \pid_side.O_2_14 ;
    wire \pid_side.error_p_regZ0Z_10 ;
    wire \pid_front.m19_2_03_0_0_1_cascade_ ;
    wire \pid_front.N_161 ;
    wire pid_side_m27_2_03_0_a2_0_0;
    wire \pid_side.N_253_cascade_ ;
    wire \pid_side.m27_2_03_0_cascade_ ;
    wire \pid_side.error_i_regZ0Z_23 ;
    wire \pid_side.N_576 ;
    wire \pid_side.m11_2_03_3_i_3 ;
    wire \pid_side.error_i_reg_esr_RNO_3Z0Z_14 ;
    wire pid_side_N_216_cascade_;
    wire \pid_side.error_i_reg_esr_RNO_6Z0Z_17_cascade_ ;
    wire \pid_side.m21_2_03_0_0 ;
    wire \pid_side.m21_2_03_0_1_cascade_ ;
    wire \pid_side.error_i_reg_esr_RNO_0_0_17 ;
    wire \pid_side.error_i_reg_esr_RNO_5Z0Z_17 ;
    wire xy_ki_fast_fast_3;
    wire pid_side_N_235;
    wire pid_side_N_235_cascade_;
    wire \pid_side.m28_2_03_0_0_cascade_ ;
    wire \pid_side.m28_2_03_0_cascade_ ;
    wire \pid_side.error_i_reg_9_rn_0_24_cascade_ ;
    wire \pid_side.error_i_regZ0Z_24 ;
    wire \pid_side.m56_0_o2_0 ;
    wire \pid_side.m56_0_o2_0_cascade_ ;
    wire \pid_side.error_i_reg_9_sn_24 ;
    wire \pid_front.m78_0_m2_1_ns_1 ;
    wire \pid_side.error_cry_2_0_c_RNI7C2SZ0_cascade_ ;
    wire \pid_side.N_155 ;
    wire \pid_side.error_cry_2_0_c_RNI7A6PZ0Z2_cascade_ ;
    wire \pid_side.N_204 ;
    wire \pid_side.N_204_cascade_ ;
    wire \pid_side.N_186 ;
    wire \pid_side.g0_16_1_cascade_ ;
    wire \pid_side.N_228_cascade_ ;
    wire \pid_side.error_i_reg_9_1_26_cascade_ ;
    wire \pid_side.error_i_regZ0Z_26 ;
    wire \pid_side.m10_2_03_3_i_0_o2_1_1_cascade_ ;
    wire \pid_side.m51_0_o2_0 ;
    wire \pid_side.N_228 ;
    wire \pid_side.error_i_regZ0Z_10 ;
    wire \pid_side.m10_2_03_3_i_3 ;
    wire \pid_side.error_i_regZ0Z_22 ;
    wire \pid_front.N_186_0 ;
    wire \pid_front.error_i_reg_esr_RNO_5_0_12 ;
    wire \pid_side.m10_2_03_3_i_0_o2_0_1_cascade_ ;
    wire \pid_side.N_185_cascade_ ;
    wire \pid_side.m11_2_03_3_i_0_o2_1 ;
    wire \pid_front.error_13 ;
    wire \pid_front.error_9 ;
    wire \pid_side.N_185 ;
    wire \pid_side.N_207 ;
    wire \pid_side.m10_2_03_3_i_0_o2_1 ;
    wire \pid_front.m78_0_a2_sx ;
    wire \pid_front.N_524 ;
    wire \pid_front.error_cry_1_c_RNIJE4MZ0Z2_cascade_ ;
    wire \pid_front.N_182 ;
    wire \pid_front.m8_2_03_3_i_0 ;
    wire \pid_front.m8_2_03_3_i_0_cascade_ ;
    wire \pid_front.error_i_regZ0Z_4 ;
    wire \pid_front.m58_0_o2_N_2LZ0Z1 ;
    wire \pid_front.error_cry_1_0_c_RNI590GZ0Z1_cascade_ ;
    wire \pid_front.N_183 ;
    wire \pid_front.error_cry_1_0_c_RNINTZ0Z963 ;
    wire \pid_front.error_1 ;
    wire \pid_front.N_40_0_i_i_o2_0_cascade_ ;
    wire \pid_front.error_3 ;
    wire \pid_front.error_cry_2_c_RNIKGVOZ0Z2_cascade_ ;
    wire \pid_front.N_245 ;
    wire \pid_front.error_i_reg_9_sn_rn_0_15_cascade_ ;
    wire \pid_front.m19_2_03_0_0 ;
    wire \pid_front.error_i_reg_9_rn_1_15 ;
    wire \pid_front.error_i_reg_9_sn_15_cascade_ ;
    wire \pid_front.m19_2_03_0_1 ;
    wire \pid_front.error_i_regZ0Z_15 ;
    wire \pid_front.N_226_cascade_ ;
    wire \pid_front.m21_2_03_0_0 ;
    wire \pid_front.m22_2_03_0_0 ;
    wire \pid_front.error_11 ;
    wire \pid_front.N_254 ;
    wire \pid_front.N_254_cascade_ ;
    wire \pid_front.error_i_reg_9_N_2L1_1_cascade_ ;
    wire \pid_front.N_226 ;
    wire \pid_front.error_i_reg_esr_RNO_0Z0Z_16 ;
    wire \pid_front.N_594 ;
    wire \pid_front.N_611 ;
    wire \pid_front.error_12 ;
    wire pid_side_N_495;
    wire \pid_front.N_569_cascade_ ;
    wire \pid_front.error_8 ;
    wire \pid_front.error_i_reg_9_sn_13 ;
    wire \pid_front.error_i_reg_9_rn_2_13 ;
    wire \pid_front.N_436_cascade_ ;
    wire \pid_front.error_i_regZ0Z_13 ;
    wire \pid_front.N_184 ;
    wire \pid_front.N_231 ;
    wire \pid_front.N_437 ;
    wire \pid_front.m10_2_03_3_i_0_a2_0 ;
    wire \pid_front.error_i_acumm_13_0_a2_2_2_2 ;
    wire \pid_front.N_603 ;
    wire \pid_front.N_603_cascade_ ;
    wire \pid_front.error_i_acumm_13_0_a2_3_1_2 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_2_c_RNI68OM ;
    wire \pid_front.error_i_acumm16lto3 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_4_c_RNICGQM ;
    wire \pid_front.error_i_acumm_preregZ0Z_5 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_5_c_RNIOULE ;
    wire \pid_front.error_i_acumm_preregZ0Z_6 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_9_c_RNIIPQK ;
    wire \pid_front.error_i_reg_esr_RNIS09UZ0Z_11 ;
    wire \pid_front.error_i_acumm_preregZ0Z_10 ;
    wire \pid_front.N_355_cascade_ ;
    wire \pid_front.error_i_acummZ0Z_10 ;
    wire \pid_front.N_203 ;
    wire \pid_front.error_i_acumm_preregZ0Z_11 ;
    wire \pid_front.N_353_cascade_ ;
    wire \pid_front.error_i_acummZ0Z_11 ;
    wire \pid_front.N_227 ;
    wire \pid_front.error_i_acumm_preregZ0Z_28 ;
    wire \pid_front.N_205 ;
    wire \pid_front.N_242_cascade_ ;
    wire \pid_front.N_285 ;
    wire \pid_front.error_i_acummZ0Z_12 ;
    wire \pid_front.N_64 ;
    wire \pid_front.error_i_reg_esr_RNIV4AUZ0Z_12 ;
    wire \pid_front.un10lto12 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_0_c_RNI9AGE ;
    wire \pid_front.error_i_acumm_preregZ0Z_1 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_1_c_RNICEHE ;
    wire \pid_front.error_i_acumm_preregZ0Z_2 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_3_c_RNI9CPM ;
    wire \pid_front.error_i_acumm_preregZ0Z_4 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_6_c_RNIIOSM ;
    wire \pid_front.error_i_acumm_preregZ0Z_7 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_7_c_RNIU6OE ;
    wire \pid_front.error_i_acumm_preregZ0Z_8 ;
    wire \pid_front.state_0_g_0 ;
    wire \pid_front.error_p_regZ0Z_18 ;
    wire \pid_front.error_d_reg_prevZ0Z_18 ;
    wire \pid_front.error_p_reg_esr_RNITCC61Z0Z_18 ;
    wire \pid_side.error_p_reg_esr_RNI6FM11Z0Z_6 ;
    wire \pid_side.error_p_reg_esr_RNI76TK1Z0Z_5 ;
    wire \pid_side.error_p_reg_esr_RNIIHEQZ0Z_4 ;
    wire \pid_side.error_p_reg_esr_RNIIHEQZ0Z_4_cascade_ ;
    wire \pid_side.error_p_reg_esr_RNI76TK1_0Z0Z_5_cascade_ ;
    wire \pid_side.error_p_reg_esr_RNIG7MC2Z0Z_5 ;
    wire \pid_side.error_p_reg_esr_RNI76TK1_0Z0Z_5 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_4_c_RNI91PN ;
    wire \pid_side.error_p_reg_esr_RNIG7MC2_0Z0Z_5 ;
    wire \pid_side.error_p_reg_esr_RNIG7MC2_0Z0Z_5_cascade_ ;
    wire \pid_side.error_p_reg_esr_RNIN4BP4Z0Z_3 ;
    wire \pid_side.error_d_reg_prevZ0Z_4 ;
    wire \pid_side.error_p_reg_esr_RNIIHEQ_0Z0Z_4 ;
    wire \pid_side.error_p_reg_esr_RNIIHEQ_0Z0Z_4_cascade_ ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_3_c_RNI6TNN ;
    wire \pid_side.error_p_reg_esr_RNISL2L4Z0Z_3 ;
    wire \pid_side.error_d_reg_prev_esr_RNIKAJOZ0Z_19 ;
    wire \pid_side.error_d_reg_prev_esr_RNIKAJO_0Z0Z_19 ;
    wire \pid_side.error_d_reg_prevZ0Z_5 ;
    wire \pid_side.error_p_reg_esr_RNI6FM11_0Z0Z_6 ;
    wire \pid_side.error_d_reg_esr_RNI2OIO_3Z0Z_13 ;
    wire \pid_side.error_d_reg_fast_esr_RNIC6BTZ0Z_12_cascade_ ;
    wire \pid_side.error_d_reg_prev_fastZ0Z_12 ;
    wire \pid_side.g1_2_1 ;
    wire \pid_side.g0_3_2_cascade_ ;
    wire \pid_side.error_i_reg_esr_RNIO6NRZ0Z_14 ;
    wire \pid_side.g1_3_cascade_ ;
    wire \pid_side.error_i_reg_esr_RNIM3MRZ0Z_13 ;
    wire \pid_side.error_p_reg_esr_RNI46CB9Z0Z_12 ;
    wire \pid_side.N_2608_0_cascade_ ;
    wire \pid_side.g0_2 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_1_c_RNI0LLN ;
    wire \pid_side.error_d_reg_prev_esr_RNI905J4Z0Z_1 ;
    wire \pid_side.error_p_reg_esr_RNIIQL11Z0Z_1_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNIBGIE2Z0Z_1 ;
    wire \pid_side.error_d_reg_prev_esr_RNIBGIE2Z0Z_1_cascade_ ;
    wire \pid_side.error_p_reg_esr_RNIIQL11_0Z0Z_1 ;
    wire \pid_side.error_d_reg_prevZ0Z_0 ;
    wire \pid_side.error_p_reg_esr_RNICBEQ_0Z0Z_2 ;
    wire pid_side_error_i_reg_9_sn_rn_1_15;
    wire \pid_side.error_i_reg_9_sn_rn_0_15_cascade_ ;
    wire \pid_side.error_i_reg_9_sn_sn_15 ;
    wire \pid_side.N_161 ;
    wire \pid_side.N_258_cascade_ ;
    wire \pid_side.error_i_reg_9_rn_1_15 ;
    wire \pid_side.m19_2_03_0_0_cascade_ ;
    wire \pid_side.error_i_reg_9_sn_15 ;
    wire \pid_side.error_i_regZ0Z_15 ;
    wire \pid_side.N_245 ;
    wire \pid_side.N_245_cascade_ ;
    wire \pid_side.N_262 ;
    wire pid_side_N_306;
    wire pid_front_N_474_1;
    wire pid_side_N_306_cascade_;
    wire \pid_side.m27_2_03_0_0 ;
    wire pid_side_N_492;
    wire \pid_side.error_i_reg_esr_RNO_5Z0Z_14_cascade_ ;
    wire \pid_side.error_i_reg_esr_RNO_4Z0Z_14 ;
    wire \pid_side.N_160 ;
    wire \pid_side.N_160_cascade_ ;
    wire \pid_side.N_224_cascade_ ;
    wire \pid_side.N_258 ;
    wire \pid_side.m17_2_03_4_0 ;
    wire pid_side_N_491_cascade_;
    wire \pid_front.m21_2_03_0_1_1_cascade_ ;
    wire \pid_front.N_163 ;
    wire \pid_front.m21_2_03_0_1 ;
    wire \pid_side.m78_0_m2_1_ns_1_cascade_ ;
    wire \pid_side.N_184_cascade_ ;
    wire \pid_side.N_229 ;
    wire \pid_side.N_437 ;
    wire dron_frame_decoder_1_source_H_disp_side_fast_0;
    wire \pid_side.error_axb_0 ;
    wire bfn_20_15_0_;
    wire \pid_side.error_axbZ0Z_1 ;
    wire \pid_side.error_cry_0 ;
    wire \pid_side.error_axbZ0Z_2 ;
    wire \pid_side.error_cry_1 ;
    wire \pid_side.error_axbZ0Z_3 ;
    wire \pid_side.error_cry_2 ;
    wire drone_H_disp_side_i_4;
    wire \pid_side.error_4 ;
    wire \pid_side.error_cry_3 ;
    wire drone_H_disp_side_i_5;
    wire \pid_side.error_cry_0_0 ;
    wire drone_H_disp_side_i_6;
    wire \pid_side.error_cry_1_0 ;
    wire drone_H_disp_side_i_7;
    wire \pid_side.error_cry_2_0 ;
    wire \pid_side.error_cry_3_0 ;
    wire drone_H_disp_side_i_8;
    wire bfn_20_16_0_;
    wire drone_H_disp_side_i_9;
    wire \pid_side.error_cry_4 ;
    wire drone_H_disp_side_i_10;
    wire \pid_side.error_cry_5 ;
    wire \pid_side.error_axbZ0Z_7 ;
    wire \pid_side.error_cry_6 ;
    wire \pid_side.error_axb_8_l_ofxZ0 ;
    wire drone_H_disp_side_12;
    wire \pid_side.error_cry_7 ;
    wire drone_H_disp_side_i_12;
    wire drone_H_disp_side_13;
    wire \pid_side.error_cry_8 ;
    wire drone_H_disp_side_i_13;
    wire \pid_side.error_cry_9 ;
    wire drone_H_disp_side_15;
    wire drone_H_disp_side_14;
    wire \pid_side.error_cry_10 ;
    wire \pid_side.N_224 ;
    wire \pid_side.m19_2_03_0_1 ;
    wire \pid_side.error_i_reg_esr_RNO_4Z0Z_22_cascade_ ;
    wire \pid_side.error_i_reg_esr_RNO_3Z0Z_22 ;
    wire \pid_side.N_297_cascade_ ;
    wire \pid_side.N_301 ;
    wire \pid_side.N_252 ;
    wire \pid_side.N_252_cascade_ ;
    wire \pid_side.m1_0_03 ;
    wire \pid_side.N_537_cascade_ ;
    wire \pid_side.N_189 ;
    wire \pid_side.m9_2_03_3_i_0_o2_0_cascade_ ;
    wire xy_ki_fast_3;
    wire \pid_front.error_10 ;
    wire \pid_front.error_i_reg_esr_RNO_6_0_12_cascade_ ;
    wire \pid_front.error_14 ;
    wire \pid_front.N_228_0 ;
    wire \pid_side.un4_error_i_reg_31_bm_sx ;
    wire \pid_front.error_i_reg_esr_RNO_4Z0Z_19 ;
    wire \pid_front.error_i_reg_esr_RNO_0Z0Z_19 ;
    wire \pid_front.error_i_reg_esr_RNO_1_0_19_cascade_ ;
    wire \pid_front.error_i_regZ0Z_19 ;
    wire \pid_front.state_ns_0_0 ;
    wire \pid_front.error_5 ;
    wire \pid_front.error_6 ;
    wire \pid_front.error_7 ;
    wire \pid_front.N_27_0_i_i_0 ;
    wire \pid_front.N_426_cascade_ ;
    wire \pid_front.error_cry_2_c_RNIKGVOZ0Z2 ;
    wire \pid_front.m7_2_01_cascade_ ;
    wire \pid_front.error_i_reg_esr_RNO_5Z0Z_19 ;
    wire \pid_front.error_i_reg_esr_RNO_2_0_19 ;
    wire \pid_front.error_i_reg_esr_RNO_3Z0Z_19 ;
    wire \pid_front.O_11 ;
    wire \pid_front.error_d_regZ0Z_8 ;
    wire \pid_front.O_6 ;
    wire \pid_front.error_d_regZ0Z_3 ;
    wire \pid_front.O_12 ;
    wire \pid_front.error_d_regZ0Z_9 ;
    wire \pid_front.error_d_reg_prevZ0Z_12 ;
    wire \pid_front.N_5_0_0 ;
    wire \pid_side.O_1_8 ;
    wire \pid_side.error_d_regZ0Z_5 ;
    wire \pid_side.O_1_9 ;
    wire \pid_side.error_d_regZ0Z_6 ;
    wire \pid_side.O_1_10 ;
    wire \pid_side.error_d_regZ0Z_7 ;
    wire \pid_side.O_2_7 ;
    wire \pid_side.error_d_reg_prev_esr_RNI9BFR3Z0Z_1 ;
    wire \pid_side.error_p_reg_esr_RNIU3T36Z0Z_2 ;
    wire \pid_side.error_p_reg_esr_RNICBEQZ0Z_2 ;
    wire \pid_side.error_p_reg_esr_RNICBEQZ0Z_2_cascade_ ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_2_c_RNIQUGJ ;
    wire \pid_side.error_p_reg_esr_RNILOD82Z0Z_2 ;
    wire \pid_side.error_p_reg_esr_RNIFEEQ_0Z0Z_3 ;
    wire \pid_side.error_d_reg_prevZ0Z_2 ;
    wire \pid_side.error_d_reg_prevZ0Z_3 ;
    wire \pid_side.error_p_regZ0Z_3 ;
    wire \pid_side.error_p_reg_esr_RNIFEEQZ0Z_3 ;
    wire \pid_side.O_1_12 ;
    wire \pid_side.error_d_regZ0Z_9 ;
    wire \pid_side.O_1_6 ;
    wire \pid_side.error_d_regZ0Z_3 ;
    wire \pid_side.error_d_reg_prevZ0Z_14 ;
    wire \pid_side.N_2608_0_0_0_cascade_ ;
    wire \pid_side.N_5_1 ;
    wire \pid_side.g0_2_0_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNI7PM14Z0Z_12 ;
    wire \pid_side.error_d_reg_prevZ0Z_13 ;
    wire \pid_side.N_4_1_0_1 ;
    wire \pid_side.error_d_reg_prevZ0Z_12 ;
    wire \pid_side.g0_1_0_1_cascade_ ;
    wire \pid_side.g0_1 ;
    wire \pid_side.O_0_3 ;
    wire \pid_side.error_d_regZ0Z_0 ;
    wire \pid_side.O_1_4 ;
    wire \pid_side.O_2_6 ;
    wire \pid_side.error_p_regZ0Z_2 ;
    wire \pid_side.error_d_reg_fastZ0Z_12 ;
    wire \pid_side.O_1_5 ;
    wire \pid_side.error_d_regZ0Z_2 ;
    wire \pid_side.N_232 ;
    wire \pid_side.N_45_i_i_0_cascade_ ;
    wire \pid_side.N_8_cascade_ ;
    wire \pid_side.error_i_reg_esr_RNO_0Z0Z_18_cascade_ ;
    wire \pid_side.error_i_regZ0Z_18 ;
    wire \pid_side.m22_2_03_0_2 ;
    wire \pid_side.error_cry_1_c_RNI6K4BZ0Z1 ;
    wire \pid_side.N_8 ;
    wire \pid_side.error_i_regZ0Z_2 ;
    wire \pid_front.error_i_reg_9_sn_sn_15 ;
    wire \pid_side.N_314_cascade_ ;
    wire \pid_side.m24_2_03_0_0_cascade_ ;
    wire \pid_side.error_i_reg_esr_RNO_6Z0Z_20_cascade_ ;
    wire \pid_side.error_i_reg_esr_RNO_5Z0Z_20 ;
    wire \pid_side.m24_2_03_0_1 ;
    wire \pid_side.N_162_cascade_ ;
    wire \pid_side.N_206 ;
    wire \pid_side.N_206_cascade_ ;
    wire \pid_side.N_629 ;
    wire \pid_side.m9_2_03_3_i_0_o2_0 ;
    wire \pid_side.m9_2_03_3_i_0_o2_2_cascade_ ;
    wire \pid_side.error_i_regZ0Z_5 ;
    wire xy_ki_fast_3_rep1;
    wire pid_side_N_496_cascade_;
    wire \pid_side.N_536 ;
    wire \pid_side.N_186_0 ;
    wire \pid_side.error_i_reg_esr_RNO_5Z0Z_12 ;
    wire \pid_side.error_9 ;
    wire \pid_side.error_13 ;
    wire \pid_side.N_606 ;
    wire \pid_side.N_606_cascade_ ;
    wire \pid_side.error_5 ;
    wire xy_ki_fast_2;
    wire \pid_side.N_188 ;
    wire \pid_side.N_231 ;
    wire \pid_side.N_231_cascade_ ;
    wire \pid_side.N_184 ;
    wire \pid_side.N_339 ;
    wire \pid_front.error_2 ;
    wire \pid_front.error_4 ;
    wire \pid_front.N_525 ;
    wire \pid_side.error_2 ;
    wire \pid_side.error_1 ;
    wire drone_H_disp_side_0;
    wire \pid_side.error_3 ;
    wire \pid_side.N_40_0_i_i_o2_1 ;
    wire \pid_side.N_40_0_i_i_o2_1_cascade_ ;
    wire \pid_side.N_40_0_i_i_o2_0 ;
    wire \pid_side.N_27_0_i_i_0 ;
    wire \pid_side.m7_2_01_ns_1_cascade_ ;
    wire \pid_side.N_162 ;
    wire \pid_side.m7_2_01 ;
    wire \pid_side.m7_2_01_cascade_ ;
    wire \pid_front.error_15 ;
    wire \pid_front.error_i_reg_9_N_5L8_0_sx ;
    wire \pid_side.error_14 ;
    wire \pid_side.error_10 ;
    wire \pid_side.N_225_cascade_ ;
    wire pid_side_N_174;
    wire \pid_side.m25_2_03_0_2_cascade_ ;
    wire \pid_side.un4_error_i_reg_31_am_1 ;
    wire \pid_side.error_i_reg_esr_RNO_0_0_21_cascade_ ;
    wire \pid_side.error_i_reg_esr_RNO_1Z0Z_21 ;
    wire \pid_side.error_i_regZ0Z_21 ;
    wire \pid_side.N_254_cascade_ ;
    wire pid_side_N_491;
    wire \pid_side.m20_2_03_0_0 ;
    wire pid_side_m20_2_03_0_a2_0_0;
    wire \pid_front.m0_0_03 ;
    wire xy_ki_fast_0;
    wire \pid_front.N_574 ;
    wire \pid_front.state_ns_0 ;
    wire pid_side_N_607;
    wire \pid_front.m7_2_01 ;
    wire \pid_front.error_i_regZ0Z_3 ;
    wire \pid_front.O_21 ;
    wire \pid_front.error_d_regZ0Z_18 ;
    wire \pid_front.O_5 ;
    wire \pid_front.error_d_regZ0Z_2 ;
    wire \pid_front.O_13 ;
    wire \pid_front.error_d_regZ0Z_10 ;
    wire \pid_front.O_15 ;
    wire \pid_front.error_d_regZ0Z_12 ;
    wire \pid_front.O_9 ;
    wire \pid_front.error_d_regZ0Z_6 ;
    wire \pid_side.O_1_11 ;
    wire \pid_side.error_d_regZ0Z_8 ;
    wire \pid_side.O_2_8 ;
    wire \pid_side.error_p_regZ0Z_4 ;
    wire \pid_side.error_d_reg_prevZ0Z_1 ;
    wire \pid_side.error_d_regZ0Z_1 ;
    wire \pid_side.error_d_reg_prev_esr_RNIIFEIZ0Z_1 ;
    wire \pid_side.error_d_reg_prev_esr_RNIH7JOZ0Z_18 ;
    wire \pid_side.error_d_reg_prevZ0Z_19 ;
    wire \pid_side.un1_pid_prereg_135_0 ;
    wire \pid_side.g0_1_0 ;
    wire \pid_side.error_d_reg_prevZ0Z_11 ;
    wire \pid_side.error_d_reg_prev_esr_RNISHIO_1Z0Z_11 ;
    wire \pid_side.error_d_reg_fastZ0Z_13 ;
    wire \pid_side.O_1_14 ;
    wire \pid_side.error_d_regZ0Z_11 ;
    wire \pid_side.m24_2_03_0 ;
    wire \pid_side.error_i_regZ0Z_20 ;
    wire \pid_side.N_156 ;
    wire \pid_side.error_7 ;
    wire \pid_side.N_551_cascade_ ;
    wire \pid_side.m8_2_03_3_i_0 ;
    wire \pid_side.N_230 ;
    wire pid_side_N_496;
    wire \pid_side.N_551 ;
    wire \pid_side.error_i_reg_esr_RNO_0Z0Z_4_cascade_ ;
    wire pid_side_N_490;
    wire \pid_side.error_i_regZ0Z_4 ;
    wire xy_ki_fast_1;
    wire xy_ki_0_rep1;
    wire \pid_side.N_183 ;
    wire \pid_side.N_538_cascade_ ;
    wire \pid_side.error_6 ;
    wire \pid_side.m58_0_o2_0 ;
    wire xy_ki_0_rep2;
    wire \pid_side.m58_0_a2_1_sxZ0 ;
    wire pid_side_N_216;
    wire drone_H_disp_front_0;
    wire \pid_front.m0_2_03 ;
    wire xy_ki_4;
    wire \pid_side.error_i_reg_9_sx_18 ;
    wire xy_ki_2;
    wire \Commands_frame_decoder.source_xy_ki_1_sqmuxa_0 ;
    wire side_command_0;
    wire uart_pc_data_1;
    wire side_command_1;
    wire side_command_2;
    wire side_command_3;
    wire side_command_4;
    wire side_command_5;
    wire side_command_6;
    wire side_command_7;
    wire \Commands_frame_decoder.source_CH2data_1_sqmuxa_0 ;
    wire \pid_side.error_8 ;
    wire xy_ki_3_rep2;
    wire \pid_side.error_12 ;
    wire \pid_side.N_226_cascade_ ;
    wire pid_side_N_164;
    wire \pid_side.N_589 ;
    wire \pid_side.N_459_cascade_ ;
    wire \pid_side.error_11 ;
    wire \pid_side.N_225 ;
    wire xy_ki_1;
    wire \pid_side.m23_2_03_0_2_cascade_ ;
    wire \pid_side.un4_error_i_reg_29_ns_sn ;
    wire \pid_side.un4_error_i_reg_29_ns_rn_0 ;
    wire pid_front_N_335;
    wire \pid_side.m23_2_03_0_1 ;
    wire \pid_side.error_i_reg_esr_RNO_2Z0Z_19_cascade_ ;
    wire \pid_side.error_i_reg_esr_RNO_1Z0Z_19 ;
    wire \pid_side.error_i_regZ0Z_19 ;
    wire \pid_side.state_ns_0_0 ;
    wire reset_module_System_reset_iso_g;
    wire \pid_side.error_15 ;
    wire \pid_side.N_622 ;
    wire pid_side_N_493;
    wire \pid_side.N_226 ;
    wire pid_side_m22_2_03_0_a2_0;
    wire \pid_side.N_254 ;
    wire \pid_side.m22_2_03_0_0 ;
    wire xy_ki_0;
    wire xy_ki_2_rep2;
    wire xy_ki_3;
    wire xy_ki_1_rep2;
    wire pid_front_N_463_1;
    wire uart_pc_data_4;
    wire xy_kd_4;
    wire uart_pc_data_5;
    wire xy_kd_5;
    wire uart_pc_data_6;
    wire xy_kd_6;
    wire uart_pc_data_0;
    wire xy_kd_0;
    wire \pid_side.N_834_0 ;
    wire \pid_side.N_2054_g ;
    wire \pid_side.O_1_7 ;
    wire \pid_side.error_d_regZ0Z_4 ;
    wire \pid_side.error_d_reg_prevZ0Z_18 ;
    wire \pid_side.error_d_reg_prev_esr_RNIH7JO_0Z0Z_18 ;
    wire \pid_side.O_2_12 ;
    wire \pid_side.error_p_regZ0Z_8 ;
    wire \pid_side.O_2_5 ;
    wire \pid_side.error_p_regZ0Z_1 ;
    wire xy_ki_1_rep1;
    wire xy_ki_2_rep1;
    wire xy_ki_3_rep1;
    wire pid_side_m24_2_03_0_a2_0;
    wire \pid_side.O_2_20 ;
    wire \pid_side.error_p_regZ0Z_16 ;
    wire \pid_side.O_2_10 ;
    wire \pid_side.error_p_regZ0Z_6 ;
    wire \pid_side.O_2_11 ;
    wire \pid_side.error_p_regZ0Z_7 ;
    wire \pid_side.O_2_13 ;
    wire \pid_side.error_p_regZ0Z_9 ;
    wire \pid_side.O_2_9 ;
    wire \pid_side.error_p_regZ0Z_5 ;
    wire \pid_side.O_2_4 ;
    wire \pid_side.error_p_regZ0Z_0 ;
    wire \pid_side.O_2_23 ;
    wire \pid_side.error_p_regZ0Z_19 ;
    wire \pid_side.O_2_15 ;
    wire \pid_side.error_p_regZ0Z_11 ;
    wire \pid_side.O_2_16 ;
    wire \pid_side.error_p_regZ0Z_12 ;
    wire \pid_side.O_2_17 ;
    wire \pid_side.error_p_regZ0Z_13 ;
    wire \pid_side.O_2_18 ;
    wire \pid_side.error_p_regZ0Z_14 ;
    wire \pid_side.O_2_19 ;
    wire \pid_side.error_p_regZ0Z_15 ;
    wire \pid_side.O_2_21 ;
    wire \pid_side.error_p_regZ0Z_17 ;
    wire \pid_side.O_2_22 ;
    wire \pid_side.error_p_regZ0Z_18 ;
    wire \pid_side.O_2_24 ;
    wire \pid_side.error_p_regZ0Z_20 ;
    wire \pid_side.O_1_18 ;
    wire \pid_side.error_d_regZ0Z_15 ;
    wire \pid_side.O_1_16 ;
    wire \pid_side.error_d_regZ0Z_13 ;
    wire \pid_side.O_1_17 ;
    wire \pid_side.error_d_regZ0Z_14 ;
    wire \pid_side.O_1_24 ;
    wire \pid_side.error_d_regZ0Z_21 ;
    wire \pid_side.O_1_15 ;
    wire \pid_side.error_d_regZ0Z_12 ;
    wire \pid_side.O_1_20 ;
    wire \pid_side.error_d_regZ0Z_17 ;
    wire \pid_side.O_1_22 ;
    wire \pid_side.error_d_regZ0Z_19 ;
    wire \pid_side.O_1_23 ;
    wire \pid_side.error_d_regZ0Z_20 ;
    wire \pid_side.O_1_21 ;
    wire \pid_side.error_d_regZ0Z_18 ;
    wire \pid_side.O_1_19 ;
    wire \pid_side.error_d_regZ0Z_16 ;
    wire \pid_side.N_868_0 ;
    wire uart_pc_data_2;
    wire xy_kd_2;
    wire uart_pc_data_3;
    wire xy_kd_3;
    wire uart_pc_data_7;
    wire xy_kd_7;
    wire \Commands_frame_decoder.state_RNITUI31Z0Z_13 ;
    wire \pid_front.O_23 ;
    wire \pid_front.error_d_regZ0Z_20 ;
    wire \pid_front.O_22 ;
    wire \pid_front.error_d_regZ0Z_19 ;
    wire \pid_front.O_24 ;
    wire \pid_front.error_d_regZ0Z_21 ;
    wire \pid_front.O_8 ;
    wire \pid_front.error_d_regZ0Z_5 ;
    wire \pid_front.O_10 ;
    wire \pid_front.error_d_regZ0Z_7 ;
    wire \pid_front.O_14 ;
    wire \pid_front.error_d_regZ0Z_11 ;
    wire \pid_front.O_17 ;
    wire \pid_front.error_d_regZ0Z_14 ;
    wire \pid_front.O_18 ;
    wire \pid_front.error_d_regZ0Z_15 ;
    wire \pid_front.O_19 ;
    wire \pid_front.error_d_regZ0Z_16 ;
    wire \pid_front.O_20 ;
    wire \pid_front.error_d_regZ0Z_17 ;
    wire _gnd_net_;
    wire clk_system_pll_g;
    wire \pid_front.N_787_0 ;
    wire N_934_g;

    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .TEST_MODE=1'b0;
    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .SHIFTREG_DIV_MODE=2'b00;
    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .PLLOUT_SELECT="GENCLK";
    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .FILTER_RANGE=3'b001;
    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .FEEDBACK_PATH="SIMPLE";
    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .FDA_RELATIVE=4'b0000;
    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .FDA_FEEDBACK=4'b0000;
    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .ENABLE_ICEGATE=1'b0;
    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .DIVR=4'b0000;
    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .DIVQ=3'b110;
    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .DIVF=7'b0111111;
    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    PLL40 \Pc2drone_pll_inst.Pc2drone_pll_inst_pll  (
            .PLLOUTGLOBAL(),
            .SDI(GNDG0),
            .BYPASS(GNDG0),
            .RESETB(N__65955),
            .PLLOUTCORE(\Pc2drone_pll_inst.clk_system_pll ),
            .LOCK(),
            .SDO(),
            .SCLK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .EXTFEEDBACK(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLIN(N__94801));
    defparam \pid_alt.un2_error_mulonly_0_24_0 .A_REG=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .NEG_TRIGGER=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .MODE_8x8=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .D_REG=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .C_REG=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .B_SIGNED=1'b1;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .B_REG=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .A_SIGNED=1'b1;
    SB_MAC16 \pid_alt.un2_error_mulonly_0_24_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__65953),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__65937),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7,dangling_wire_8,dangling_wire_9,dangling_wire_10,dangling_wire_11,dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15}),
            .ADDSUBBOT(),
            .A({N__38171,N__38222,N__38270,N__38318,N__38366,N__38408,N__38453,N__38505,N__38543,N__37806,N__37847,N__37895,N__37946,N__37988,N__38027,N__48384}),
            .C({dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29,dangling_wire_30,dangling_wire_31}),
            .B({dangling_wire_32,dangling_wire_33,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39,N__36307,N__34804,N__36319,N__52081,N__34780,N__40318,N__34792,N__36295}),
            .OHOLDTOP(),
            .O({dangling_wire_40,dangling_wire_41,dangling_wire_42,dangling_wire_43,dangling_wire_44,dangling_wire_45,dangling_wire_46,\pid_alt.O_5_24 ,\pid_alt.O_5_23 ,\pid_alt.O_5_22 ,\pid_alt.O_5_21 ,\pid_alt.O_5_20 ,\pid_alt.O_5_19 ,\pid_alt.O_5_18 ,\pid_alt.O_5_17 ,\pid_alt.O_5_16 ,\pid_alt.O_5_15 ,\pid_alt.O_5_14 ,\pid_alt.O_5_13 ,\pid_alt.O_5_12 ,\pid_alt.O_5_11 ,\pid_alt.O_5_10 ,\pid_alt.O_5_9 ,\pid_alt.O_5_8 ,\pid_alt.O_5_7 ,\pid_alt.O_5_6 ,\pid_alt.O_5_5 ,\pid_alt.O_5_4 ,dangling_wire_47,dangling_wire_48,dangling_wire_49,dangling_wire_50}));
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .A_REG=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .NEG_TRIGGER=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .MODE_8x8=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .D_REG=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .C_REG=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .B_SIGNED=1'b1;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .B_REG=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .A_SIGNED=1'b1;
    SB_MAC16 \pid_alt.un2_error_2_mulonly_0_24_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__65907),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__65845),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_51,dangling_wire_52,dangling_wire_53,dangling_wire_54,dangling_wire_55,dangling_wire_56,dangling_wire_57,dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66}),
            .ADDSUBBOT(),
            .A({N__38179,N__38226,N__38275,N__38323,N__38371,N__38416,N__38461,N__38504,N__38551,N__37810,N__37855,N__37903,N__37951,N__37993,N__38038,N__48400}),
            .C({dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73,dangling_wire_74,dangling_wire_75,dangling_wire_76,dangling_wire_77,dangling_wire_78,dangling_wire_79,dangling_wire_80,dangling_wire_81,dangling_wire_82}),
            .B({dangling_wire_83,dangling_wire_84,dangling_wire_85,dangling_wire_86,dangling_wire_87,dangling_wire_88,dangling_wire_89,dangling_wire_90,N__33739,N__33751,N__33763,N__33775,N__33787,N__33799,N__33811,N__33823}),
            .OHOLDTOP(),
            .O({dangling_wire_91,dangling_wire_92,dangling_wire_93,dangling_wire_94,dangling_wire_95,dangling_wire_96,dangling_wire_97,\pid_alt.O_3_24 ,\pid_alt.O_3_23 ,\pid_alt.O_3_22 ,\pid_alt.O_3_21 ,\pid_alt.O_3_20 ,\pid_alt.O_3_19 ,\pid_alt.O_3_18 ,\pid_alt.O_3_17 ,\pid_alt.O_3_16 ,\pid_alt.O_3_15 ,\pid_alt.O_3_14 ,\pid_alt.O_3_13 ,\pid_alt.O_3_12 ,\pid_alt.O_3_11 ,\pid_alt.O_3_10 ,\pid_alt.O_3_9 ,\pid_alt.O_3_8 ,\pid_alt.O_3_7 ,\pid_alt.O_3_6 ,\pid_alt.O_3_5 ,\pid_alt.O_3_4 ,dangling_wire_98,dangling_wire_99,dangling_wire_100,dangling_wire_101}));
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .A_REG=1'b0;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .NEG_TRIGGER=1'b0;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .MODE_8x8=1'b0;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .D_REG=1'b0;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .C_REG=1'b0;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .B_SIGNED=1'b1;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .B_REG=1'b0;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .A_SIGNED=1'b1;
    SB_MAC16 \pid_side.un2_error_1_mulonly_0_24_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__65917),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__65956),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,dangling_wire_107,dangling_wire_108,dangling_wire_109,dangling_wire_110,dangling_wire_111,dangling_wire_112,dangling_wire_113,dangling_wire_114,dangling_wire_115,dangling_wire_116,dangling_wire_117}),
            .ADDSUBBOT(),
            .A({N__85936,N__81649,N__80418,N__84933,N__87561,N__81533,N__80491,N__85250,N__83640,N__82860,N__80313,N__77232,N__80868,N__81099,N__81022,N__80934}),
            .C({dangling_wire_118,dangling_wire_119,dangling_wire_120,dangling_wire_121,dangling_wire_122,dangling_wire_123,dangling_wire_124,dangling_wire_125,dangling_wire_126,dangling_wire_127,dangling_wire_128,dangling_wire_129,dangling_wire_130,dangling_wire_131,dangling_wire_132,dangling_wire_133}),
            .B({dangling_wire_134,dangling_wire_135,dangling_wire_136,dangling_wire_137,dangling_wire_138,dangling_wire_139,dangling_wire_140,dangling_wire_141,N__91957,N__88348,N__88534,N__88722,N__92152,N__92356,N__46113,N__88144}),
            .OHOLDTOP(),
            .O({dangling_wire_142,dangling_wire_143,dangling_wire_144,dangling_wire_145,dangling_wire_146,dangling_wire_147,dangling_wire_148,\pid_side.O_1_24 ,\pid_side.O_1_23 ,\pid_side.O_1_22 ,\pid_side.O_1_21 ,\pid_side.O_1_20 ,\pid_side.O_1_19 ,\pid_side.O_1_18 ,\pid_side.O_1_17 ,\pid_side.O_1_16 ,\pid_side.O_1_15 ,\pid_side.O_1_14 ,\pid_side.O_1_13 ,\pid_side.O_1_12 ,\pid_side.O_1_11 ,\pid_side.O_1_10 ,\pid_side.O_1_9 ,\pid_side.O_1_8 ,\pid_side.O_1_7 ,\pid_side.O_1_6 ,\pid_side.O_1_5 ,\pid_side.O_1_4 ,\pid_side.O_0_3 ,dangling_wire_149,dangling_wire_150,dangling_wire_151}));
    defparam \pid_side.un2_error_mulonly_0_24_0 .A_REG=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pid_side.un2_error_mulonly_0_24_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pid_side.un2_error_mulonly_0_24_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pid_side.un2_error_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .NEG_TRIGGER=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .MODE_8x8=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .D_REG=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .C_REG=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .B_SIGNED=1'b1;
    defparam \pid_side.un2_error_mulonly_0_24_0 .B_REG=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pid_side.un2_error_mulonly_0_24_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pid_side.un2_error_mulonly_0_24_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pid_side.un2_error_mulonly_0_24_0 .A_SIGNED=1'b1;
    SB_MAC16 \pid_side.un2_error_mulonly_0_24_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__65949),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__65948),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_152,dangling_wire_153,dangling_wire_154,dangling_wire_155,dangling_wire_156,dangling_wire_157,dangling_wire_158,dangling_wire_159,dangling_wire_160,dangling_wire_161,dangling_wire_162,dangling_wire_163,dangling_wire_164,dangling_wire_165,dangling_wire_166,dangling_wire_167}),
            .ADDSUBBOT(),
            .A({N__85937,N__81655,N__80419,N__84932,N__87562,N__81535,N__80490,N__85251,N__83641,N__82861,N__80314,N__77233,N__80869,N__81110,N__81025,N__80950}),
            .C({dangling_wire_168,dangling_wire_169,dangling_wire_170,dangling_wire_171,dangling_wire_172,dangling_wire_173,dangling_wire_174,dangling_wire_175,dangling_wire_176,dangling_wire_177,dangling_wire_178,dangling_wire_179,dangling_wire_180,dangling_wire_181,dangling_wire_182,dangling_wire_183}),
            .B({dangling_wire_184,dangling_wire_185,dangling_wire_186,dangling_wire_187,dangling_wire_188,dangling_wire_189,dangling_wire_190,dangling_wire_191,N__45577,N__45613,N__45645,N__52027,N__45685,N__45307,N__45339,N__45379}),
            .OHOLDTOP(),
            .O({dangling_wire_192,dangling_wire_193,dangling_wire_194,dangling_wire_195,dangling_wire_196,dangling_wire_197,dangling_wire_198,\pid_side.O_2_24 ,\pid_side.O_2_23 ,\pid_side.O_2_22 ,\pid_side.O_2_21 ,\pid_side.O_2_20 ,\pid_side.O_2_19 ,\pid_side.O_2_18 ,\pid_side.O_2_17 ,\pid_side.O_2_16 ,\pid_side.O_2_15 ,\pid_side.O_2_14 ,\pid_side.O_2_13 ,\pid_side.O_2_12 ,\pid_side.O_2_11 ,\pid_side.O_2_10 ,\pid_side.O_2_9 ,\pid_side.O_2_8 ,\pid_side.O_2_7 ,\pid_side.O_2_6 ,\pid_side.O_2_5 ,\pid_side.O_2_4 ,dangling_wire_199,dangling_wire_200,dangling_wire_201,dangling_wire_202}));
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .A_REG=1'b0;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .NEG_TRIGGER=1'b0;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .MODE_8x8=1'b0;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .D_REG=1'b0;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .C_REG=1'b0;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .B_SIGNED=1'b1;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .B_REG=1'b0;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .A_SIGNED=1'b1;
    SB_MAC16 \pid_front.un2_error_1_mulonly_0_24_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__65954),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__65941),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_203,dangling_wire_204,dangling_wire_205,dangling_wire_206,dangling_wire_207,dangling_wire_208,dangling_wire_209,dangling_wire_210,dangling_wire_211,dangling_wire_212,dangling_wire_213,dangling_wire_214,dangling_wire_215,dangling_wire_216,dangling_wire_217,dangling_wire_218}),
            .ADDSUBBOT(),
            .A({N__80704,N__78319,N__73915,N__74320,N__74518,N__78418,N__73801,N__74871,N__77747,N__77872,N__77983,N__79915,N__74086,N__80017,N__74188,N__84662}),
            .C({dangling_wire_219,dangling_wire_220,dangling_wire_221,dangling_wire_222,dangling_wire_223,dangling_wire_224,dangling_wire_225,dangling_wire_226,dangling_wire_227,dangling_wire_228,dangling_wire_229,dangling_wire_230,dangling_wire_231,dangling_wire_232,dangling_wire_233,dangling_wire_234}),
            .B({dangling_wire_235,dangling_wire_236,dangling_wire_237,dangling_wire_238,dangling_wire_239,dangling_wire_240,dangling_wire_241,dangling_wire_242,N__91956,N__88344,N__88530,N__88726,N__92151,N__92355,N__46117,N__88140}),
            .OHOLDTOP(),
            .O({dangling_wire_243,dangling_wire_244,dangling_wire_245,dangling_wire_246,dangling_wire_247,dangling_wire_248,dangling_wire_249,\pid_front.O_24 ,\pid_front.O_23 ,\pid_front.O_22 ,\pid_front.O_21 ,\pid_front.O_20 ,\pid_front.O_19 ,\pid_front.O_18 ,\pid_front.O_17 ,\pid_front.O_16 ,\pid_front.O_15 ,\pid_front.O_14 ,\pid_front.O_13 ,\pid_front.O_12 ,\pid_front.O_11 ,\pid_front.O_10 ,\pid_front.O_9 ,\pid_front.O_8 ,\pid_front.O_7 ,\pid_front.O_6 ,\pid_front.O_5 ,\pid_front.O_4 ,\pid_front.O_3 ,dangling_wire_250,dangling_wire_251,dangling_wire_252}));
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .A_REG=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .NEG_TRIGGER=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .MODE_8x8=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .D_REG=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .C_REG=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .B_SIGNED=1'b1;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .B_REG=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .A_SIGNED=1'b1;
    SB_MAC16 \pid_alt.un2_error_1_mulonly_0_24_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__65874),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__65829),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_253,dangling_wire_254,dangling_wire_255,dangling_wire_256,dangling_wire_257,dangling_wire_258,dangling_wire_259,dangling_wire_260,dangling_wire_261,dangling_wire_262,dangling_wire_263,dangling_wire_264,dangling_wire_265,dangling_wire_266,dangling_wire_267,dangling_wire_268}),
            .ADDSUBBOT(),
            .A({N__38172,N__38227,N__38271,N__38319,N__38367,N__38409,N__38454,N__38506,N__38544,N__37802,N__37848,N__37896,N__37947,N__37989,N__38034,N__48396}),
            .C({dangling_wire_269,dangling_wire_270,dangling_wire_271,dangling_wire_272,dangling_wire_273,dangling_wire_274,dangling_wire_275,dangling_wire_276,dangling_wire_277,dangling_wire_278,dangling_wire_279,dangling_wire_280,dangling_wire_281,dangling_wire_282,dangling_wire_283,dangling_wire_284}),
            .B({dangling_wire_285,dangling_wire_286,dangling_wire_287,dangling_wire_288,dangling_wire_289,dangling_wire_290,dangling_wire_291,dangling_wire_292,N__34858,N__33883,N__33892,N__34873,N__34885,N__34897,N__34909,N__34921}),
            .OHOLDTOP(),
            .O({dangling_wire_293,dangling_wire_294,dangling_wire_295,dangling_wire_296,dangling_wire_297,dangling_wire_298,dangling_wire_299,\pid_alt.O_4_24 ,\pid_alt.O_4_23 ,\pid_alt.O_4_22 ,\pid_alt.O_4_21 ,\pid_alt.O_4_20 ,\pid_alt.O_4_19 ,\pid_alt.O_4_18 ,\pid_alt.O_4_17 ,\pid_alt.O_4_16 ,\pid_alt.O_4_15 ,\pid_alt.O_4_14 ,\pid_alt.O_4_13 ,\pid_alt.O_4_12 ,\pid_alt.O_4_11 ,\pid_alt.O_4_10 ,\pid_alt.O_4_9 ,\pid_alt.O_4_8 ,\pid_alt.O_4_7 ,\pid_alt.O_4_6 ,\pid_alt.O_4_5 ,\pid_alt.O_4_4 ,dangling_wire_300,dangling_wire_301,dangling_wire_302,dangling_wire_303}));
    defparam \pid_front.un2_error_mulonly_0_24_0 .A_REG=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pid_front.un2_error_mulonly_0_24_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pid_front.un2_error_mulonly_0_24_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pid_front.un2_error_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .NEG_TRIGGER=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .MODE_8x8=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .D_REG=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .C_REG=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .B_SIGNED=1'b1;
    defparam \pid_front.un2_error_mulonly_0_24_0 .B_REG=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pid_front.un2_error_mulonly_0_24_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pid_front.un2_error_mulonly_0_24_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pid_front.un2_error_mulonly_0_24_0 .A_SIGNED=1'b1;
    SB_MAC16 \pid_front.un2_error_mulonly_0_24_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__65936),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__65878),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_304,dangling_wire_305,dangling_wire_306,dangling_wire_307,dangling_wire_308,dangling_wire_309,dangling_wire_310,dangling_wire_311,dangling_wire_312,dangling_wire_313,dangling_wire_314,dangling_wire_315,dangling_wire_316,dangling_wire_317,dangling_wire_318,dangling_wire_319}),
            .ADDSUBBOT(),
            .A({N__80697,N__78324,N__73908,N__74313,N__74514,N__78391,N__73797,N__74857,N__77749,N__77867,N__77982,N__79914,N__74066,N__80013,N__74184,N__84661}),
            .C({dangling_wire_320,dangling_wire_321,dangling_wire_322,dangling_wire_323,dangling_wire_324,dangling_wire_325,dangling_wire_326,dangling_wire_327,dangling_wire_328,dangling_wire_329,dangling_wire_330,dangling_wire_331,dangling_wire_332,dangling_wire_333,dangling_wire_334,dangling_wire_335}),
            .B({dangling_wire_336,dangling_wire_337,dangling_wire_338,dangling_wire_339,dangling_wire_340,dangling_wire_341,dangling_wire_342,dangling_wire_343,N__45570,N__45606,N__45646,N__52017,N__45681,N__45297,N__45340,N__45375}),
            .OHOLDTOP(),
            .O({dangling_wire_344,dangling_wire_345,dangling_wire_346,dangling_wire_347,dangling_wire_348,dangling_wire_349,dangling_wire_350,\pid_front.O_0_24 ,\pid_front.O_0_23 ,\pid_front.O_0_22 ,\pid_front.O_0_21 ,\pid_front.O_0_20 ,\pid_front.O_0_19 ,\pid_front.O_0_18 ,\pid_front.O_0_17 ,\pid_front.O_0_16 ,\pid_front.O_0_15 ,\pid_front.O_0_14 ,\pid_front.O_0_13 ,\pid_front.O_0_12 ,\pid_front.O_0_11 ,\pid_front.O_0_10 ,\pid_front.O_0_9 ,\pid_front.O_0_8 ,\pid_front.O_0_7 ,\pid_front.O_0_6 ,\pid_front.O_0_5 ,\pid_front.O_0_4 ,dangling_wire_351,dangling_wire_352,dangling_wire_353,dangling_wire_354}));
    IO_PAD \Pc2drone_pll_inst.Pc2drone_pll_inst_iopad  (
            .OE(VCCG0),
            .DIN(),
            .DOUT(N__94801),
            .PACKAGEPIN(clk_system));
    defparam uart_input_pc_ibuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD uart_input_pc_ibuf_iopad (
            .OE(N__94787),
            .DIN(N__94786),
            .DOUT(N__94785),
            .PACKAGEPIN(uart_input_pc));
    defparam uart_input_pc_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam uart_input_pc_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO uart_input_pc_ibuf_preio (
            .PADOEN(N__94787),
            .PADOUT(N__94786),
            .PADIN(N__94785),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(uart_input_pc_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_CH2_18A_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_CH2_18A_obuf_iopad (
            .OE(N__94778),
            .DIN(N__94777),
            .DOUT(N__94776),
            .PACKAGEPIN(debug_CH2_18A));
    defparam debug_CH2_18A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_CH2_18A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_CH2_18A_obuf_preio (
            .PADOEN(N__94778),
            .PADOUT(N__94777),
            .PADIN(N__94776),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__52249),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ppm_output_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD ppm_output_obuf_iopad (
            .OE(N__94769),
            .DIN(N__94768),
            .DOUT(N__94767),
            .PACKAGEPIN(ppm_output));
    defparam ppm_output_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ppm_output_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ppm_output_obuf_preio (
            .PADOEN(N__94769),
            .PADOUT(N__94768),
            .PADIN(N__94767),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__49822),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_CH3_20A_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_CH3_20A_obuf_iopad (
            .OE(N__94760),
            .DIN(N__94759),
            .DOUT(N__94758),
            .PACKAGEPIN(debug_CH3_20A));
    defparam debug_CH3_20A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_CH3_20A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_CH3_20A_obuf_preio (
            .PADOEN(N__94760),
            .PADOUT(N__94759),
            .PADIN(N__94758),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__48118),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_CH6_5B_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_CH6_5B_obuf_iopad (
            .OE(N__94751),
            .DIN(N__94750),
            .DOUT(N__94749),
            .PACKAGEPIN(debug_CH6_5B));
    defparam debug_CH6_5B_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_CH6_5B_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_CH6_5B_obuf_preio (
            .PADOEN(N__94751),
            .PADOUT(N__94750),
            .PADIN(N__94749),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam uart_input_drone_ibuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD uart_input_drone_ibuf_iopad (
            .OE(N__94742),
            .DIN(N__94741),
            .DOUT(N__94740),
            .PACKAGEPIN(uart_input_drone));
    defparam uart_input_drone_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam uart_input_drone_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO uart_input_drone_ibuf_preio (
            .PADOEN(N__94742),
            .PADOUT(N__94741),
            .PADIN(N__94740),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(uart_input_drone_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_CH0_16A_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_CH0_16A_obuf_iopad (
            .OE(N__94733),
            .DIN(N__94732),
            .DOUT(N__94731),
            .PACKAGEPIN(debug_CH0_16A));
    defparam debug_CH0_16A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_CH0_16A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_CH0_16A_obuf_preio (
            .PADOEN(N__94733),
            .PADOUT(N__94732),
            .PADIN(N__94731),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__56878),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_CH1_0A_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_CH1_0A_obuf_iopad (
            .OE(N__94724),
            .DIN(N__94723),
            .DOUT(N__94722),
            .PACKAGEPIN(debug_CH1_0A));
    defparam debug_CH1_0A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_CH1_0A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_CH1_0A_obuf_preio (
            .PADOEN(N__94724),
            .PADOUT(N__94723),
            .PADIN(N__94722),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__69202),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_CH5_31B_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_CH5_31B_obuf_iopad (
            .OE(N__94715),
            .DIN(N__94714),
            .DOUT(N__94713),
            .PACKAGEPIN(debug_CH5_31B));
    defparam debug_CH5_31B_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_CH5_31B_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_CH5_31B_obuf_preio (
            .PADOEN(N__94715),
            .PADOUT(N__94714),
            .PADIN(N__94713),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_CH4_2A_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_CH4_2A_obuf_iopad (
            .OE(N__94706),
            .DIN(N__94705),
            .DOUT(N__94704),
            .PACKAGEPIN(debug_CH4_2A));
    defparam debug_CH4_2A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_CH4_2A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_CH4_2A_obuf_preio (
            .PADOEN(N__94706),
            .PADOUT(N__94705),
            .PADIN(N__94704),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__23254 (
            .O(N__94687),
            .I(N__94684));
    LocalMux I__23253 (
            .O(N__94684),
            .I(\pid_front.O_8 ));
    CascadeMux I__23252 (
            .O(N__94681),
            .I(N__94675));
    InMux I__23251 (
            .O(N__94680),
            .I(N__94670));
    InMux I__23250 (
            .O(N__94679),
            .I(N__94670));
    InMux I__23249 (
            .O(N__94678),
            .I(N__94665));
    InMux I__23248 (
            .O(N__94675),
            .I(N__94665));
    LocalMux I__23247 (
            .O(N__94670),
            .I(N__94660));
    LocalMux I__23246 (
            .O(N__94665),
            .I(N__94657));
    InMux I__23245 (
            .O(N__94664),
            .I(N__94652));
    InMux I__23244 (
            .O(N__94663),
            .I(N__94652));
    Span4Mux_h I__23243 (
            .O(N__94660),
            .I(N__94649));
    Span4Mux_h I__23242 (
            .O(N__94657),
            .I(N__94646));
    LocalMux I__23241 (
            .O(N__94652),
            .I(N__94643));
    Span4Mux_h I__23240 (
            .O(N__94649),
            .I(N__94640));
    Span4Mux_h I__23239 (
            .O(N__94646),
            .I(N__94637));
    Span12Mux_h I__23238 (
            .O(N__94643),
            .I(N__94634));
    Span4Mux_h I__23237 (
            .O(N__94640),
            .I(N__94629));
    Span4Mux_h I__23236 (
            .O(N__94637),
            .I(N__94629));
    Odrv12 I__23235 (
            .O(N__94634),
            .I(\pid_front.error_d_regZ0Z_5 ));
    Odrv4 I__23234 (
            .O(N__94629),
            .I(\pid_front.error_d_regZ0Z_5 ));
    InMux I__23233 (
            .O(N__94624),
            .I(N__94621));
    LocalMux I__23232 (
            .O(N__94621),
            .I(\pid_front.O_10 ));
    InMux I__23231 (
            .O(N__94618),
            .I(N__94606));
    InMux I__23230 (
            .O(N__94617),
            .I(N__94606));
    InMux I__23229 (
            .O(N__94616),
            .I(N__94606));
    InMux I__23228 (
            .O(N__94615),
            .I(N__94606));
    LocalMux I__23227 (
            .O(N__94606),
            .I(N__94603));
    Span12Mux_h I__23226 (
            .O(N__94603),
            .I(N__94600));
    Odrv12 I__23225 (
            .O(N__94600),
            .I(\pid_front.error_d_regZ0Z_7 ));
    InMux I__23224 (
            .O(N__94597),
            .I(N__94594));
    LocalMux I__23223 (
            .O(N__94594),
            .I(\pid_front.O_14 ));
    InMux I__23222 (
            .O(N__94591),
            .I(N__94582));
    InMux I__23221 (
            .O(N__94590),
            .I(N__94582));
    InMux I__23220 (
            .O(N__94589),
            .I(N__94577));
    InMux I__23219 (
            .O(N__94588),
            .I(N__94577));
    InMux I__23218 (
            .O(N__94587),
            .I(N__94574));
    LocalMux I__23217 (
            .O(N__94582),
            .I(N__94571));
    LocalMux I__23216 (
            .O(N__94577),
            .I(N__94568));
    LocalMux I__23215 (
            .O(N__94574),
            .I(N__94565));
    Span4Mux_h I__23214 (
            .O(N__94571),
            .I(N__94560));
    Span4Mux_v I__23213 (
            .O(N__94568),
            .I(N__94560));
    Span4Mux_h I__23212 (
            .O(N__94565),
            .I(N__94557));
    Span4Mux_h I__23211 (
            .O(N__94560),
            .I(N__94554));
    Span4Mux_h I__23210 (
            .O(N__94557),
            .I(N__94551));
    Odrv4 I__23209 (
            .O(N__94554),
            .I(\pid_front.error_d_regZ0Z_11 ));
    Odrv4 I__23208 (
            .O(N__94551),
            .I(\pid_front.error_d_regZ0Z_11 ));
    InMux I__23207 (
            .O(N__94546),
            .I(N__94543));
    LocalMux I__23206 (
            .O(N__94543),
            .I(\pid_front.O_17 ));
    InMux I__23205 (
            .O(N__94540),
            .I(N__94537));
    LocalMux I__23204 (
            .O(N__94537),
            .I(N__94532));
    InMux I__23203 (
            .O(N__94536),
            .I(N__94529));
    InMux I__23202 (
            .O(N__94535),
            .I(N__94526));
    Span4Mux_v I__23201 (
            .O(N__94532),
            .I(N__94521));
    LocalMux I__23200 (
            .O(N__94529),
            .I(N__94521));
    LocalMux I__23199 (
            .O(N__94526),
            .I(N__94514));
    Sp12to4 I__23198 (
            .O(N__94521),
            .I(N__94514));
    InMux I__23197 (
            .O(N__94520),
            .I(N__94509));
    InMux I__23196 (
            .O(N__94519),
            .I(N__94509));
    Span12Mux_s6_v I__23195 (
            .O(N__94514),
            .I(N__94504));
    LocalMux I__23194 (
            .O(N__94509),
            .I(N__94504));
    Odrv12 I__23193 (
            .O(N__94504),
            .I(\pid_front.error_d_regZ0Z_14 ));
    InMux I__23192 (
            .O(N__94501),
            .I(N__94498));
    LocalMux I__23191 (
            .O(N__94498),
            .I(\pid_front.O_18 ));
    InMux I__23190 (
            .O(N__94495),
            .I(N__94492));
    LocalMux I__23189 (
            .O(N__94492),
            .I(N__94489));
    Span4Mux_v I__23188 (
            .O(N__94489),
            .I(N__94484));
    InMux I__23187 (
            .O(N__94488),
            .I(N__94479));
    InMux I__23186 (
            .O(N__94487),
            .I(N__94479));
    Sp12to4 I__23185 (
            .O(N__94484),
            .I(N__94474));
    LocalMux I__23184 (
            .O(N__94479),
            .I(N__94474));
    Odrv12 I__23183 (
            .O(N__94474),
            .I(\pid_front.error_d_regZ0Z_15 ));
    InMux I__23182 (
            .O(N__94471),
            .I(N__94468));
    LocalMux I__23181 (
            .O(N__94468),
            .I(\pid_front.O_19 ));
    InMux I__23180 (
            .O(N__94465),
            .I(N__94456));
    InMux I__23179 (
            .O(N__94464),
            .I(N__94456));
    InMux I__23178 (
            .O(N__94463),
            .I(N__94456));
    LocalMux I__23177 (
            .O(N__94456),
            .I(N__94453));
    Span4Mux_h I__23176 (
            .O(N__94453),
            .I(N__94450));
    Span4Mux_h I__23175 (
            .O(N__94450),
            .I(N__94447));
    Span4Mux_h I__23174 (
            .O(N__94447),
            .I(N__94444));
    Odrv4 I__23173 (
            .O(N__94444),
            .I(\pid_front.error_d_regZ0Z_16 ));
    InMux I__23172 (
            .O(N__94441),
            .I(N__94438));
    LocalMux I__23171 (
            .O(N__94438),
            .I(\pid_front.O_20 ));
    InMux I__23170 (
            .O(N__94435),
            .I(N__94426));
    InMux I__23169 (
            .O(N__94434),
            .I(N__94426));
    InMux I__23168 (
            .O(N__94433),
            .I(N__94426));
    LocalMux I__23167 (
            .O(N__94426),
            .I(N__94423));
    Span4Mux_h I__23166 (
            .O(N__94423),
            .I(N__94420));
    Span4Mux_h I__23165 (
            .O(N__94420),
            .I(N__94417));
    Span4Mux_h I__23164 (
            .O(N__94417),
            .I(N__94414));
    Odrv4 I__23163 (
            .O(N__94414),
            .I(\pid_front.error_d_regZ0Z_17 ));
    ClkMux I__23162 (
            .O(N__94411),
            .I(N__93415));
    ClkMux I__23161 (
            .O(N__94410),
            .I(N__93415));
    ClkMux I__23160 (
            .O(N__94409),
            .I(N__93415));
    ClkMux I__23159 (
            .O(N__94408),
            .I(N__93415));
    ClkMux I__23158 (
            .O(N__94407),
            .I(N__93415));
    ClkMux I__23157 (
            .O(N__94406),
            .I(N__93415));
    ClkMux I__23156 (
            .O(N__94405),
            .I(N__93415));
    ClkMux I__23155 (
            .O(N__94404),
            .I(N__93415));
    ClkMux I__23154 (
            .O(N__94403),
            .I(N__93415));
    ClkMux I__23153 (
            .O(N__94402),
            .I(N__93415));
    ClkMux I__23152 (
            .O(N__94401),
            .I(N__93415));
    ClkMux I__23151 (
            .O(N__94400),
            .I(N__93415));
    ClkMux I__23150 (
            .O(N__94399),
            .I(N__93415));
    ClkMux I__23149 (
            .O(N__94398),
            .I(N__93415));
    ClkMux I__23148 (
            .O(N__94397),
            .I(N__93415));
    ClkMux I__23147 (
            .O(N__94396),
            .I(N__93415));
    ClkMux I__23146 (
            .O(N__94395),
            .I(N__93415));
    ClkMux I__23145 (
            .O(N__94394),
            .I(N__93415));
    ClkMux I__23144 (
            .O(N__94393),
            .I(N__93415));
    ClkMux I__23143 (
            .O(N__94392),
            .I(N__93415));
    ClkMux I__23142 (
            .O(N__94391),
            .I(N__93415));
    ClkMux I__23141 (
            .O(N__94390),
            .I(N__93415));
    ClkMux I__23140 (
            .O(N__94389),
            .I(N__93415));
    ClkMux I__23139 (
            .O(N__94388),
            .I(N__93415));
    ClkMux I__23138 (
            .O(N__94387),
            .I(N__93415));
    ClkMux I__23137 (
            .O(N__94386),
            .I(N__93415));
    ClkMux I__23136 (
            .O(N__94385),
            .I(N__93415));
    ClkMux I__23135 (
            .O(N__94384),
            .I(N__93415));
    ClkMux I__23134 (
            .O(N__94383),
            .I(N__93415));
    ClkMux I__23133 (
            .O(N__94382),
            .I(N__93415));
    ClkMux I__23132 (
            .O(N__94381),
            .I(N__93415));
    ClkMux I__23131 (
            .O(N__94380),
            .I(N__93415));
    ClkMux I__23130 (
            .O(N__94379),
            .I(N__93415));
    ClkMux I__23129 (
            .O(N__94378),
            .I(N__93415));
    ClkMux I__23128 (
            .O(N__94377),
            .I(N__93415));
    ClkMux I__23127 (
            .O(N__94376),
            .I(N__93415));
    ClkMux I__23126 (
            .O(N__94375),
            .I(N__93415));
    ClkMux I__23125 (
            .O(N__94374),
            .I(N__93415));
    ClkMux I__23124 (
            .O(N__94373),
            .I(N__93415));
    ClkMux I__23123 (
            .O(N__94372),
            .I(N__93415));
    ClkMux I__23122 (
            .O(N__94371),
            .I(N__93415));
    ClkMux I__23121 (
            .O(N__94370),
            .I(N__93415));
    ClkMux I__23120 (
            .O(N__94369),
            .I(N__93415));
    ClkMux I__23119 (
            .O(N__94368),
            .I(N__93415));
    ClkMux I__23118 (
            .O(N__94367),
            .I(N__93415));
    ClkMux I__23117 (
            .O(N__94366),
            .I(N__93415));
    ClkMux I__23116 (
            .O(N__94365),
            .I(N__93415));
    ClkMux I__23115 (
            .O(N__94364),
            .I(N__93415));
    ClkMux I__23114 (
            .O(N__94363),
            .I(N__93415));
    ClkMux I__23113 (
            .O(N__94362),
            .I(N__93415));
    ClkMux I__23112 (
            .O(N__94361),
            .I(N__93415));
    ClkMux I__23111 (
            .O(N__94360),
            .I(N__93415));
    ClkMux I__23110 (
            .O(N__94359),
            .I(N__93415));
    ClkMux I__23109 (
            .O(N__94358),
            .I(N__93415));
    ClkMux I__23108 (
            .O(N__94357),
            .I(N__93415));
    ClkMux I__23107 (
            .O(N__94356),
            .I(N__93415));
    ClkMux I__23106 (
            .O(N__94355),
            .I(N__93415));
    ClkMux I__23105 (
            .O(N__94354),
            .I(N__93415));
    ClkMux I__23104 (
            .O(N__94353),
            .I(N__93415));
    ClkMux I__23103 (
            .O(N__94352),
            .I(N__93415));
    ClkMux I__23102 (
            .O(N__94351),
            .I(N__93415));
    ClkMux I__23101 (
            .O(N__94350),
            .I(N__93415));
    ClkMux I__23100 (
            .O(N__94349),
            .I(N__93415));
    ClkMux I__23099 (
            .O(N__94348),
            .I(N__93415));
    ClkMux I__23098 (
            .O(N__94347),
            .I(N__93415));
    ClkMux I__23097 (
            .O(N__94346),
            .I(N__93415));
    ClkMux I__23096 (
            .O(N__94345),
            .I(N__93415));
    ClkMux I__23095 (
            .O(N__94344),
            .I(N__93415));
    ClkMux I__23094 (
            .O(N__94343),
            .I(N__93415));
    ClkMux I__23093 (
            .O(N__94342),
            .I(N__93415));
    ClkMux I__23092 (
            .O(N__94341),
            .I(N__93415));
    ClkMux I__23091 (
            .O(N__94340),
            .I(N__93415));
    ClkMux I__23090 (
            .O(N__94339),
            .I(N__93415));
    ClkMux I__23089 (
            .O(N__94338),
            .I(N__93415));
    ClkMux I__23088 (
            .O(N__94337),
            .I(N__93415));
    ClkMux I__23087 (
            .O(N__94336),
            .I(N__93415));
    ClkMux I__23086 (
            .O(N__94335),
            .I(N__93415));
    ClkMux I__23085 (
            .O(N__94334),
            .I(N__93415));
    ClkMux I__23084 (
            .O(N__94333),
            .I(N__93415));
    ClkMux I__23083 (
            .O(N__94332),
            .I(N__93415));
    ClkMux I__23082 (
            .O(N__94331),
            .I(N__93415));
    ClkMux I__23081 (
            .O(N__94330),
            .I(N__93415));
    ClkMux I__23080 (
            .O(N__94329),
            .I(N__93415));
    ClkMux I__23079 (
            .O(N__94328),
            .I(N__93415));
    ClkMux I__23078 (
            .O(N__94327),
            .I(N__93415));
    ClkMux I__23077 (
            .O(N__94326),
            .I(N__93415));
    ClkMux I__23076 (
            .O(N__94325),
            .I(N__93415));
    ClkMux I__23075 (
            .O(N__94324),
            .I(N__93415));
    ClkMux I__23074 (
            .O(N__94323),
            .I(N__93415));
    ClkMux I__23073 (
            .O(N__94322),
            .I(N__93415));
    ClkMux I__23072 (
            .O(N__94321),
            .I(N__93415));
    ClkMux I__23071 (
            .O(N__94320),
            .I(N__93415));
    ClkMux I__23070 (
            .O(N__94319),
            .I(N__93415));
    ClkMux I__23069 (
            .O(N__94318),
            .I(N__93415));
    ClkMux I__23068 (
            .O(N__94317),
            .I(N__93415));
    ClkMux I__23067 (
            .O(N__94316),
            .I(N__93415));
    ClkMux I__23066 (
            .O(N__94315),
            .I(N__93415));
    ClkMux I__23065 (
            .O(N__94314),
            .I(N__93415));
    ClkMux I__23064 (
            .O(N__94313),
            .I(N__93415));
    ClkMux I__23063 (
            .O(N__94312),
            .I(N__93415));
    ClkMux I__23062 (
            .O(N__94311),
            .I(N__93415));
    ClkMux I__23061 (
            .O(N__94310),
            .I(N__93415));
    ClkMux I__23060 (
            .O(N__94309),
            .I(N__93415));
    ClkMux I__23059 (
            .O(N__94308),
            .I(N__93415));
    ClkMux I__23058 (
            .O(N__94307),
            .I(N__93415));
    ClkMux I__23057 (
            .O(N__94306),
            .I(N__93415));
    ClkMux I__23056 (
            .O(N__94305),
            .I(N__93415));
    ClkMux I__23055 (
            .O(N__94304),
            .I(N__93415));
    ClkMux I__23054 (
            .O(N__94303),
            .I(N__93415));
    ClkMux I__23053 (
            .O(N__94302),
            .I(N__93415));
    ClkMux I__23052 (
            .O(N__94301),
            .I(N__93415));
    ClkMux I__23051 (
            .O(N__94300),
            .I(N__93415));
    ClkMux I__23050 (
            .O(N__94299),
            .I(N__93415));
    ClkMux I__23049 (
            .O(N__94298),
            .I(N__93415));
    ClkMux I__23048 (
            .O(N__94297),
            .I(N__93415));
    ClkMux I__23047 (
            .O(N__94296),
            .I(N__93415));
    ClkMux I__23046 (
            .O(N__94295),
            .I(N__93415));
    ClkMux I__23045 (
            .O(N__94294),
            .I(N__93415));
    ClkMux I__23044 (
            .O(N__94293),
            .I(N__93415));
    ClkMux I__23043 (
            .O(N__94292),
            .I(N__93415));
    ClkMux I__23042 (
            .O(N__94291),
            .I(N__93415));
    ClkMux I__23041 (
            .O(N__94290),
            .I(N__93415));
    ClkMux I__23040 (
            .O(N__94289),
            .I(N__93415));
    ClkMux I__23039 (
            .O(N__94288),
            .I(N__93415));
    ClkMux I__23038 (
            .O(N__94287),
            .I(N__93415));
    ClkMux I__23037 (
            .O(N__94286),
            .I(N__93415));
    ClkMux I__23036 (
            .O(N__94285),
            .I(N__93415));
    ClkMux I__23035 (
            .O(N__94284),
            .I(N__93415));
    ClkMux I__23034 (
            .O(N__94283),
            .I(N__93415));
    ClkMux I__23033 (
            .O(N__94282),
            .I(N__93415));
    ClkMux I__23032 (
            .O(N__94281),
            .I(N__93415));
    ClkMux I__23031 (
            .O(N__94280),
            .I(N__93415));
    ClkMux I__23030 (
            .O(N__94279),
            .I(N__93415));
    ClkMux I__23029 (
            .O(N__94278),
            .I(N__93415));
    ClkMux I__23028 (
            .O(N__94277),
            .I(N__93415));
    ClkMux I__23027 (
            .O(N__94276),
            .I(N__93415));
    ClkMux I__23026 (
            .O(N__94275),
            .I(N__93415));
    ClkMux I__23025 (
            .O(N__94274),
            .I(N__93415));
    ClkMux I__23024 (
            .O(N__94273),
            .I(N__93415));
    ClkMux I__23023 (
            .O(N__94272),
            .I(N__93415));
    ClkMux I__23022 (
            .O(N__94271),
            .I(N__93415));
    ClkMux I__23021 (
            .O(N__94270),
            .I(N__93415));
    ClkMux I__23020 (
            .O(N__94269),
            .I(N__93415));
    ClkMux I__23019 (
            .O(N__94268),
            .I(N__93415));
    ClkMux I__23018 (
            .O(N__94267),
            .I(N__93415));
    ClkMux I__23017 (
            .O(N__94266),
            .I(N__93415));
    ClkMux I__23016 (
            .O(N__94265),
            .I(N__93415));
    ClkMux I__23015 (
            .O(N__94264),
            .I(N__93415));
    ClkMux I__23014 (
            .O(N__94263),
            .I(N__93415));
    ClkMux I__23013 (
            .O(N__94262),
            .I(N__93415));
    ClkMux I__23012 (
            .O(N__94261),
            .I(N__93415));
    ClkMux I__23011 (
            .O(N__94260),
            .I(N__93415));
    ClkMux I__23010 (
            .O(N__94259),
            .I(N__93415));
    ClkMux I__23009 (
            .O(N__94258),
            .I(N__93415));
    ClkMux I__23008 (
            .O(N__94257),
            .I(N__93415));
    ClkMux I__23007 (
            .O(N__94256),
            .I(N__93415));
    ClkMux I__23006 (
            .O(N__94255),
            .I(N__93415));
    ClkMux I__23005 (
            .O(N__94254),
            .I(N__93415));
    ClkMux I__23004 (
            .O(N__94253),
            .I(N__93415));
    ClkMux I__23003 (
            .O(N__94252),
            .I(N__93415));
    ClkMux I__23002 (
            .O(N__94251),
            .I(N__93415));
    ClkMux I__23001 (
            .O(N__94250),
            .I(N__93415));
    ClkMux I__23000 (
            .O(N__94249),
            .I(N__93415));
    ClkMux I__22999 (
            .O(N__94248),
            .I(N__93415));
    ClkMux I__22998 (
            .O(N__94247),
            .I(N__93415));
    ClkMux I__22997 (
            .O(N__94246),
            .I(N__93415));
    ClkMux I__22996 (
            .O(N__94245),
            .I(N__93415));
    ClkMux I__22995 (
            .O(N__94244),
            .I(N__93415));
    ClkMux I__22994 (
            .O(N__94243),
            .I(N__93415));
    ClkMux I__22993 (
            .O(N__94242),
            .I(N__93415));
    ClkMux I__22992 (
            .O(N__94241),
            .I(N__93415));
    ClkMux I__22991 (
            .O(N__94240),
            .I(N__93415));
    ClkMux I__22990 (
            .O(N__94239),
            .I(N__93415));
    ClkMux I__22989 (
            .O(N__94238),
            .I(N__93415));
    ClkMux I__22988 (
            .O(N__94237),
            .I(N__93415));
    ClkMux I__22987 (
            .O(N__94236),
            .I(N__93415));
    ClkMux I__22986 (
            .O(N__94235),
            .I(N__93415));
    ClkMux I__22985 (
            .O(N__94234),
            .I(N__93415));
    ClkMux I__22984 (
            .O(N__94233),
            .I(N__93415));
    ClkMux I__22983 (
            .O(N__94232),
            .I(N__93415));
    ClkMux I__22982 (
            .O(N__94231),
            .I(N__93415));
    ClkMux I__22981 (
            .O(N__94230),
            .I(N__93415));
    ClkMux I__22980 (
            .O(N__94229),
            .I(N__93415));
    ClkMux I__22979 (
            .O(N__94228),
            .I(N__93415));
    ClkMux I__22978 (
            .O(N__94227),
            .I(N__93415));
    ClkMux I__22977 (
            .O(N__94226),
            .I(N__93415));
    ClkMux I__22976 (
            .O(N__94225),
            .I(N__93415));
    ClkMux I__22975 (
            .O(N__94224),
            .I(N__93415));
    ClkMux I__22974 (
            .O(N__94223),
            .I(N__93415));
    ClkMux I__22973 (
            .O(N__94222),
            .I(N__93415));
    ClkMux I__22972 (
            .O(N__94221),
            .I(N__93415));
    ClkMux I__22971 (
            .O(N__94220),
            .I(N__93415));
    ClkMux I__22970 (
            .O(N__94219),
            .I(N__93415));
    ClkMux I__22969 (
            .O(N__94218),
            .I(N__93415));
    ClkMux I__22968 (
            .O(N__94217),
            .I(N__93415));
    ClkMux I__22967 (
            .O(N__94216),
            .I(N__93415));
    ClkMux I__22966 (
            .O(N__94215),
            .I(N__93415));
    ClkMux I__22965 (
            .O(N__94214),
            .I(N__93415));
    ClkMux I__22964 (
            .O(N__94213),
            .I(N__93415));
    ClkMux I__22963 (
            .O(N__94212),
            .I(N__93415));
    ClkMux I__22962 (
            .O(N__94211),
            .I(N__93415));
    ClkMux I__22961 (
            .O(N__94210),
            .I(N__93415));
    ClkMux I__22960 (
            .O(N__94209),
            .I(N__93415));
    ClkMux I__22959 (
            .O(N__94208),
            .I(N__93415));
    ClkMux I__22958 (
            .O(N__94207),
            .I(N__93415));
    ClkMux I__22957 (
            .O(N__94206),
            .I(N__93415));
    ClkMux I__22956 (
            .O(N__94205),
            .I(N__93415));
    ClkMux I__22955 (
            .O(N__94204),
            .I(N__93415));
    ClkMux I__22954 (
            .O(N__94203),
            .I(N__93415));
    ClkMux I__22953 (
            .O(N__94202),
            .I(N__93415));
    ClkMux I__22952 (
            .O(N__94201),
            .I(N__93415));
    ClkMux I__22951 (
            .O(N__94200),
            .I(N__93415));
    ClkMux I__22950 (
            .O(N__94199),
            .I(N__93415));
    ClkMux I__22949 (
            .O(N__94198),
            .I(N__93415));
    ClkMux I__22948 (
            .O(N__94197),
            .I(N__93415));
    ClkMux I__22947 (
            .O(N__94196),
            .I(N__93415));
    ClkMux I__22946 (
            .O(N__94195),
            .I(N__93415));
    ClkMux I__22945 (
            .O(N__94194),
            .I(N__93415));
    ClkMux I__22944 (
            .O(N__94193),
            .I(N__93415));
    ClkMux I__22943 (
            .O(N__94192),
            .I(N__93415));
    ClkMux I__22942 (
            .O(N__94191),
            .I(N__93415));
    ClkMux I__22941 (
            .O(N__94190),
            .I(N__93415));
    ClkMux I__22940 (
            .O(N__94189),
            .I(N__93415));
    ClkMux I__22939 (
            .O(N__94188),
            .I(N__93415));
    ClkMux I__22938 (
            .O(N__94187),
            .I(N__93415));
    ClkMux I__22937 (
            .O(N__94186),
            .I(N__93415));
    ClkMux I__22936 (
            .O(N__94185),
            .I(N__93415));
    ClkMux I__22935 (
            .O(N__94184),
            .I(N__93415));
    ClkMux I__22934 (
            .O(N__94183),
            .I(N__93415));
    ClkMux I__22933 (
            .O(N__94182),
            .I(N__93415));
    ClkMux I__22932 (
            .O(N__94181),
            .I(N__93415));
    ClkMux I__22931 (
            .O(N__94180),
            .I(N__93415));
    ClkMux I__22930 (
            .O(N__94179),
            .I(N__93415));
    ClkMux I__22929 (
            .O(N__94178),
            .I(N__93415));
    ClkMux I__22928 (
            .O(N__94177),
            .I(N__93415));
    ClkMux I__22927 (
            .O(N__94176),
            .I(N__93415));
    ClkMux I__22926 (
            .O(N__94175),
            .I(N__93415));
    ClkMux I__22925 (
            .O(N__94174),
            .I(N__93415));
    ClkMux I__22924 (
            .O(N__94173),
            .I(N__93415));
    ClkMux I__22923 (
            .O(N__94172),
            .I(N__93415));
    ClkMux I__22922 (
            .O(N__94171),
            .I(N__93415));
    ClkMux I__22921 (
            .O(N__94170),
            .I(N__93415));
    ClkMux I__22920 (
            .O(N__94169),
            .I(N__93415));
    ClkMux I__22919 (
            .O(N__94168),
            .I(N__93415));
    ClkMux I__22918 (
            .O(N__94167),
            .I(N__93415));
    ClkMux I__22917 (
            .O(N__94166),
            .I(N__93415));
    ClkMux I__22916 (
            .O(N__94165),
            .I(N__93415));
    ClkMux I__22915 (
            .O(N__94164),
            .I(N__93415));
    ClkMux I__22914 (
            .O(N__94163),
            .I(N__93415));
    ClkMux I__22913 (
            .O(N__94162),
            .I(N__93415));
    ClkMux I__22912 (
            .O(N__94161),
            .I(N__93415));
    ClkMux I__22911 (
            .O(N__94160),
            .I(N__93415));
    ClkMux I__22910 (
            .O(N__94159),
            .I(N__93415));
    ClkMux I__22909 (
            .O(N__94158),
            .I(N__93415));
    ClkMux I__22908 (
            .O(N__94157),
            .I(N__93415));
    ClkMux I__22907 (
            .O(N__94156),
            .I(N__93415));
    ClkMux I__22906 (
            .O(N__94155),
            .I(N__93415));
    ClkMux I__22905 (
            .O(N__94154),
            .I(N__93415));
    ClkMux I__22904 (
            .O(N__94153),
            .I(N__93415));
    ClkMux I__22903 (
            .O(N__94152),
            .I(N__93415));
    ClkMux I__22902 (
            .O(N__94151),
            .I(N__93415));
    ClkMux I__22901 (
            .O(N__94150),
            .I(N__93415));
    ClkMux I__22900 (
            .O(N__94149),
            .I(N__93415));
    ClkMux I__22899 (
            .O(N__94148),
            .I(N__93415));
    ClkMux I__22898 (
            .O(N__94147),
            .I(N__93415));
    ClkMux I__22897 (
            .O(N__94146),
            .I(N__93415));
    ClkMux I__22896 (
            .O(N__94145),
            .I(N__93415));
    ClkMux I__22895 (
            .O(N__94144),
            .I(N__93415));
    ClkMux I__22894 (
            .O(N__94143),
            .I(N__93415));
    ClkMux I__22893 (
            .O(N__94142),
            .I(N__93415));
    ClkMux I__22892 (
            .O(N__94141),
            .I(N__93415));
    ClkMux I__22891 (
            .O(N__94140),
            .I(N__93415));
    ClkMux I__22890 (
            .O(N__94139),
            .I(N__93415));
    ClkMux I__22889 (
            .O(N__94138),
            .I(N__93415));
    ClkMux I__22888 (
            .O(N__94137),
            .I(N__93415));
    ClkMux I__22887 (
            .O(N__94136),
            .I(N__93415));
    ClkMux I__22886 (
            .O(N__94135),
            .I(N__93415));
    ClkMux I__22885 (
            .O(N__94134),
            .I(N__93415));
    ClkMux I__22884 (
            .O(N__94133),
            .I(N__93415));
    ClkMux I__22883 (
            .O(N__94132),
            .I(N__93415));
    ClkMux I__22882 (
            .O(N__94131),
            .I(N__93415));
    ClkMux I__22881 (
            .O(N__94130),
            .I(N__93415));
    ClkMux I__22880 (
            .O(N__94129),
            .I(N__93415));
    ClkMux I__22879 (
            .O(N__94128),
            .I(N__93415));
    ClkMux I__22878 (
            .O(N__94127),
            .I(N__93415));
    ClkMux I__22877 (
            .O(N__94126),
            .I(N__93415));
    ClkMux I__22876 (
            .O(N__94125),
            .I(N__93415));
    ClkMux I__22875 (
            .O(N__94124),
            .I(N__93415));
    ClkMux I__22874 (
            .O(N__94123),
            .I(N__93415));
    ClkMux I__22873 (
            .O(N__94122),
            .I(N__93415));
    ClkMux I__22872 (
            .O(N__94121),
            .I(N__93415));
    ClkMux I__22871 (
            .O(N__94120),
            .I(N__93415));
    ClkMux I__22870 (
            .O(N__94119),
            .I(N__93415));
    ClkMux I__22869 (
            .O(N__94118),
            .I(N__93415));
    ClkMux I__22868 (
            .O(N__94117),
            .I(N__93415));
    ClkMux I__22867 (
            .O(N__94116),
            .I(N__93415));
    ClkMux I__22866 (
            .O(N__94115),
            .I(N__93415));
    ClkMux I__22865 (
            .O(N__94114),
            .I(N__93415));
    ClkMux I__22864 (
            .O(N__94113),
            .I(N__93415));
    ClkMux I__22863 (
            .O(N__94112),
            .I(N__93415));
    ClkMux I__22862 (
            .O(N__94111),
            .I(N__93415));
    ClkMux I__22861 (
            .O(N__94110),
            .I(N__93415));
    ClkMux I__22860 (
            .O(N__94109),
            .I(N__93415));
    ClkMux I__22859 (
            .O(N__94108),
            .I(N__93415));
    ClkMux I__22858 (
            .O(N__94107),
            .I(N__93415));
    ClkMux I__22857 (
            .O(N__94106),
            .I(N__93415));
    ClkMux I__22856 (
            .O(N__94105),
            .I(N__93415));
    ClkMux I__22855 (
            .O(N__94104),
            .I(N__93415));
    ClkMux I__22854 (
            .O(N__94103),
            .I(N__93415));
    ClkMux I__22853 (
            .O(N__94102),
            .I(N__93415));
    ClkMux I__22852 (
            .O(N__94101),
            .I(N__93415));
    ClkMux I__22851 (
            .O(N__94100),
            .I(N__93415));
    ClkMux I__22850 (
            .O(N__94099),
            .I(N__93415));
    ClkMux I__22849 (
            .O(N__94098),
            .I(N__93415));
    ClkMux I__22848 (
            .O(N__94097),
            .I(N__93415));
    ClkMux I__22847 (
            .O(N__94096),
            .I(N__93415));
    ClkMux I__22846 (
            .O(N__94095),
            .I(N__93415));
    ClkMux I__22845 (
            .O(N__94094),
            .I(N__93415));
    ClkMux I__22844 (
            .O(N__94093),
            .I(N__93415));
    ClkMux I__22843 (
            .O(N__94092),
            .I(N__93415));
    ClkMux I__22842 (
            .O(N__94091),
            .I(N__93415));
    ClkMux I__22841 (
            .O(N__94090),
            .I(N__93415));
    ClkMux I__22840 (
            .O(N__94089),
            .I(N__93415));
    ClkMux I__22839 (
            .O(N__94088),
            .I(N__93415));
    ClkMux I__22838 (
            .O(N__94087),
            .I(N__93415));
    ClkMux I__22837 (
            .O(N__94086),
            .I(N__93415));
    ClkMux I__22836 (
            .O(N__94085),
            .I(N__93415));
    ClkMux I__22835 (
            .O(N__94084),
            .I(N__93415));
    ClkMux I__22834 (
            .O(N__94083),
            .I(N__93415));
    ClkMux I__22833 (
            .O(N__94082),
            .I(N__93415));
    ClkMux I__22832 (
            .O(N__94081),
            .I(N__93415));
    ClkMux I__22831 (
            .O(N__94080),
            .I(N__93415));
    GlobalMux I__22830 (
            .O(N__93415),
            .I(N__93412));
    gio2CtrlBuf I__22829 (
            .O(N__93412),
            .I(clk_system_pll_g));
    CEMux I__22828 (
            .O(N__93409),
            .I(N__93403));
    CEMux I__22827 (
            .O(N__93408),
            .I(N__93400));
    CEMux I__22826 (
            .O(N__93407),
            .I(N__93396));
    CEMux I__22825 (
            .O(N__93406),
            .I(N__93391));
    LocalMux I__22824 (
            .O(N__93403),
            .I(N__93387));
    LocalMux I__22823 (
            .O(N__93400),
            .I(N__93383));
    CEMux I__22822 (
            .O(N__93399),
            .I(N__93380));
    LocalMux I__22821 (
            .O(N__93396),
            .I(N__93377));
    CEMux I__22820 (
            .O(N__93395),
            .I(N__93374));
    CEMux I__22819 (
            .O(N__93394),
            .I(N__93371));
    LocalMux I__22818 (
            .O(N__93391),
            .I(N__93363));
    CEMux I__22817 (
            .O(N__93390),
            .I(N__93360));
    Span4Mux_v I__22816 (
            .O(N__93387),
            .I(N__93357));
    CEMux I__22815 (
            .O(N__93386),
            .I(N__93352));
    Span4Mux_v I__22814 (
            .O(N__93383),
            .I(N__93347));
    LocalMux I__22813 (
            .O(N__93380),
            .I(N__93347));
    Span4Mux_s1_h I__22812 (
            .O(N__93377),
            .I(N__93342));
    LocalMux I__22811 (
            .O(N__93374),
            .I(N__93342));
    LocalMux I__22810 (
            .O(N__93371),
            .I(N__93339));
    CEMux I__22809 (
            .O(N__93370),
            .I(N__93336));
    CEMux I__22808 (
            .O(N__93369),
            .I(N__93333));
    CEMux I__22807 (
            .O(N__93368),
            .I(N__93329));
    CEMux I__22806 (
            .O(N__93367),
            .I(N__93326));
    CEMux I__22805 (
            .O(N__93366),
            .I(N__93323));
    Span4Mux_h I__22804 (
            .O(N__93363),
            .I(N__93318));
    LocalMux I__22803 (
            .O(N__93360),
            .I(N__93318));
    Span4Mux_h I__22802 (
            .O(N__93357),
            .I(N__93312));
    CEMux I__22801 (
            .O(N__93356),
            .I(N__93309));
    CEMux I__22800 (
            .O(N__93355),
            .I(N__93306));
    LocalMux I__22799 (
            .O(N__93352),
            .I(N__93303));
    Span4Mux_h I__22798 (
            .O(N__93347),
            .I(N__93298));
    Span4Mux_h I__22797 (
            .O(N__93342),
            .I(N__93298));
    Span4Mux_h I__22796 (
            .O(N__93339),
            .I(N__93293));
    LocalMux I__22795 (
            .O(N__93336),
            .I(N__93293));
    LocalMux I__22794 (
            .O(N__93333),
            .I(N__93290));
    CEMux I__22793 (
            .O(N__93332),
            .I(N__93287));
    LocalMux I__22792 (
            .O(N__93329),
            .I(N__93282));
    LocalMux I__22791 (
            .O(N__93326),
            .I(N__93282));
    LocalMux I__22790 (
            .O(N__93323),
            .I(N__93279));
    Span4Mux_v I__22789 (
            .O(N__93318),
            .I(N__93276));
    CEMux I__22788 (
            .O(N__93317),
            .I(N__93273));
    CEMux I__22787 (
            .O(N__93316),
            .I(N__93270));
    CEMux I__22786 (
            .O(N__93315),
            .I(N__93267));
    Span4Mux_h I__22785 (
            .O(N__93312),
            .I(N__93262));
    LocalMux I__22784 (
            .O(N__93309),
            .I(N__93262));
    LocalMux I__22783 (
            .O(N__93306),
            .I(N__93259));
    Span4Mux_h I__22782 (
            .O(N__93303),
            .I(N__93255));
    Span4Mux_h I__22781 (
            .O(N__93298),
            .I(N__93252));
    Span4Mux_h I__22780 (
            .O(N__93293),
            .I(N__93249));
    Span4Mux_v I__22779 (
            .O(N__93290),
            .I(N__93246));
    LocalMux I__22778 (
            .O(N__93287),
            .I(N__93241));
    Span4Mux_v I__22777 (
            .O(N__93282),
            .I(N__93241));
    Span4Mux_v I__22776 (
            .O(N__93279),
            .I(N__93238));
    Span4Mux_v I__22775 (
            .O(N__93276),
            .I(N__93235));
    LocalMux I__22774 (
            .O(N__93273),
            .I(N__93232));
    LocalMux I__22773 (
            .O(N__93270),
            .I(N__93227));
    LocalMux I__22772 (
            .O(N__93267),
            .I(N__93227));
    Span4Mux_v I__22771 (
            .O(N__93262),
            .I(N__93224));
    Span4Mux_v I__22770 (
            .O(N__93259),
            .I(N__93221));
    CEMux I__22769 (
            .O(N__93258),
            .I(N__93218));
    Span4Mux_h I__22768 (
            .O(N__93255),
            .I(N__93211));
    Span4Mux_h I__22767 (
            .O(N__93252),
            .I(N__93211));
    Span4Mux_v I__22766 (
            .O(N__93249),
            .I(N__93211));
    Sp12to4 I__22765 (
            .O(N__93246),
            .I(N__93202));
    Sp12to4 I__22764 (
            .O(N__93241),
            .I(N__93202));
    Sp12to4 I__22763 (
            .O(N__93238),
            .I(N__93202));
    Sp12to4 I__22762 (
            .O(N__93235),
            .I(N__93202));
    Sp12to4 I__22761 (
            .O(N__93232),
            .I(N__93199));
    Span4Mux_h I__22760 (
            .O(N__93227),
            .I(N__93196));
    Span4Mux_v I__22759 (
            .O(N__93224),
            .I(N__93193));
    Span4Mux_h I__22758 (
            .O(N__93221),
            .I(N__93190));
    LocalMux I__22757 (
            .O(N__93218),
            .I(N__93187));
    Sp12to4 I__22756 (
            .O(N__93211),
            .I(N__93180));
    Span12Mux_h I__22755 (
            .O(N__93202),
            .I(N__93180));
    Span12Mux_s8_v I__22754 (
            .O(N__93199),
            .I(N__93180));
    Span4Mux_h I__22753 (
            .O(N__93196),
            .I(N__93177));
    Span4Mux_v I__22752 (
            .O(N__93193),
            .I(N__93170));
    Span4Mux_h I__22751 (
            .O(N__93190),
            .I(N__93170));
    Span4Mux_v I__22750 (
            .O(N__93187),
            .I(N__93170));
    Odrv12 I__22749 (
            .O(N__93180),
            .I(\pid_front.N_787_0 ));
    Odrv4 I__22748 (
            .O(N__93177),
            .I(\pid_front.N_787_0 ));
    Odrv4 I__22747 (
            .O(N__93170),
            .I(\pid_front.N_787_0 ));
    InMux I__22746 (
            .O(N__93163),
            .I(N__93114));
    InMux I__22745 (
            .O(N__93162),
            .I(N__93114));
    InMux I__22744 (
            .O(N__93161),
            .I(N__93114));
    InMux I__22743 (
            .O(N__93160),
            .I(N__93109));
    InMux I__22742 (
            .O(N__93159),
            .I(N__93109));
    InMux I__22741 (
            .O(N__93158),
            .I(N__93106));
    InMux I__22740 (
            .O(N__93157),
            .I(N__93103));
    InMux I__22739 (
            .O(N__93156),
            .I(N__93098));
    InMux I__22738 (
            .O(N__93155),
            .I(N__93098));
    InMux I__22737 (
            .O(N__93154),
            .I(N__93095));
    InMux I__22736 (
            .O(N__93153),
            .I(N__93092));
    InMux I__22735 (
            .O(N__93152),
            .I(N__93087));
    InMux I__22734 (
            .O(N__93151),
            .I(N__93087));
    InMux I__22733 (
            .O(N__93150),
            .I(N__93084));
    InMux I__22732 (
            .O(N__93149),
            .I(N__93081));
    InMux I__22731 (
            .O(N__93148),
            .I(N__93066));
    InMux I__22730 (
            .O(N__93147),
            .I(N__93066));
    InMux I__22729 (
            .O(N__93146),
            .I(N__93066));
    InMux I__22728 (
            .O(N__93145),
            .I(N__93066));
    InMux I__22727 (
            .O(N__93144),
            .I(N__93066));
    InMux I__22726 (
            .O(N__93143),
            .I(N__93066));
    InMux I__22725 (
            .O(N__93142),
            .I(N__93066));
    InMux I__22724 (
            .O(N__93141),
            .I(N__93061));
    InMux I__22723 (
            .O(N__93140),
            .I(N__93061));
    InMux I__22722 (
            .O(N__93139),
            .I(N__93048));
    InMux I__22721 (
            .O(N__93138),
            .I(N__93048));
    InMux I__22720 (
            .O(N__93137),
            .I(N__93048));
    InMux I__22719 (
            .O(N__93136),
            .I(N__93048));
    InMux I__22718 (
            .O(N__93135),
            .I(N__93048));
    InMux I__22717 (
            .O(N__93134),
            .I(N__93048));
    InMux I__22716 (
            .O(N__93133),
            .I(N__93031));
    InMux I__22715 (
            .O(N__93132),
            .I(N__93031));
    InMux I__22714 (
            .O(N__93131),
            .I(N__93031));
    InMux I__22713 (
            .O(N__93130),
            .I(N__93031));
    InMux I__22712 (
            .O(N__93129),
            .I(N__93031));
    InMux I__22711 (
            .O(N__93128),
            .I(N__93031));
    InMux I__22710 (
            .O(N__93127),
            .I(N__93031));
    InMux I__22709 (
            .O(N__93126),
            .I(N__93031));
    InMux I__22708 (
            .O(N__93125),
            .I(N__93026));
    InMux I__22707 (
            .O(N__93124),
            .I(N__93026));
    InMux I__22706 (
            .O(N__93123),
            .I(N__93023));
    InMux I__22705 (
            .O(N__93122),
            .I(N__93020));
    InMux I__22704 (
            .O(N__93121),
            .I(N__93017));
    LocalMux I__22703 (
            .O(N__93114),
            .I(N__92962));
    LocalMux I__22702 (
            .O(N__93109),
            .I(N__92959));
    LocalMux I__22701 (
            .O(N__93106),
            .I(N__92956));
    LocalMux I__22700 (
            .O(N__93103),
            .I(N__92953));
    LocalMux I__22699 (
            .O(N__93098),
            .I(N__92950));
    LocalMux I__22698 (
            .O(N__93095),
            .I(N__92947));
    LocalMux I__22697 (
            .O(N__93092),
            .I(N__92944));
    LocalMux I__22696 (
            .O(N__93087),
            .I(N__92941));
    LocalMux I__22695 (
            .O(N__93084),
            .I(N__92938));
    LocalMux I__22694 (
            .O(N__93081),
            .I(N__92935));
    LocalMux I__22693 (
            .O(N__93066),
            .I(N__92932));
    LocalMux I__22692 (
            .O(N__93061),
            .I(N__92929));
    LocalMux I__22691 (
            .O(N__93048),
            .I(N__92926));
    LocalMux I__22690 (
            .O(N__93031),
            .I(N__92923));
    LocalMux I__22689 (
            .O(N__93026),
            .I(N__92920));
    LocalMux I__22688 (
            .O(N__93023),
            .I(N__92917));
    LocalMux I__22687 (
            .O(N__93020),
            .I(N__92914));
    LocalMux I__22686 (
            .O(N__93017),
            .I(N__92911));
    SRMux I__22685 (
            .O(N__93016),
            .I(N__92770));
    SRMux I__22684 (
            .O(N__93015),
            .I(N__92770));
    SRMux I__22683 (
            .O(N__93014),
            .I(N__92770));
    SRMux I__22682 (
            .O(N__93013),
            .I(N__92770));
    SRMux I__22681 (
            .O(N__93012),
            .I(N__92770));
    SRMux I__22680 (
            .O(N__93011),
            .I(N__92770));
    SRMux I__22679 (
            .O(N__93010),
            .I(N__92770));
    SRMux I__22678 (
            .O(N__93009),
            .I(N__92770));
    SRMux I__22677 (
            .O(N__93008),
            .I(N__92770));
    SRMux I__22676 (
            .O(N__93007),
            .I(N__92770));
    SRMux I__22675 (
            .O(N__93006),
            .I(N__92770));
    SRMux I__22674 (
            .O(N__93005),
            .I(N__92770));
    SRMux I__22673 (
            .O(N__93004),
            .I(N__92770));
    SRMux I__22672 (
            .O(N__93003),
            .I(N__92770));
    SRMux I__22671 (
            .O(N__93002),
            .I(N__92770));
    SRMux I__22670 (
            .O(N__93001),
            .I(N__92770));
    SRMux I__22669 (
            .O(N__93000),
            .I(N__92770));
    SRMux I__22668 (
            .O(N__92999),
            .I(N__92770));
    SRMux I__22667 (
            .O(N__92998),
            .I(N__92770));
    SRMux I__22666 (
            .O(N__92997),
            .I(N__92770));
    SRMux I__22665 (
            .O(N__92996),
            .I(N__92770));
    SRMux I__22664 (
            .O(N__92995),
            .I(N__92770));
    SRMux I__22663 (
            .O(N__92994),
            .I(N__92770));
    SRMux I__22662 (
            .O(N__92993),
            .I(N__92770));
    SRMux I__22661 (
            .O(N__92992),
            .I(N__92770));
    SRMux I__22660 (
            .O(N__92991),
            .I(N__92770));
    SRMux I__22659 (
            .O(N__92990),
            .I(N__92770));
    SRMux I__22658 (
            .O(N__92989),
            .I(N__92770));
    SRMux I__22657 (
            .O(N__92988),
            .I(N__92770));
    SRMux I__22656 (
            .O(N__92987),
            .I(N__92770));
    SRMux I__22655 (
            .O(N__92986),
            .I(N__92770));
    SRMux I__22654 (
            .O(N__92985),
            .I(N__92770));
    SRMux I__22653 (
            .O(N__92984),
            .I(N__92770));
    SRMux I__22652 (
            .O(N__92983),
            .I(N__92770));
    SRMux I__22651 (
            .O(N__92982),
            .I(N__92770));
    SRMux I__22650 (
            .O(N__92981),
            .I(N__92770));
    SRMux I__22649 (
            .O(N__92980),
            .I(N__92770));
    SRMux I__22648 (
            .O(N__92979),
            .I(N__92770));
    SRMux I__22647 (
            .O(N__92978),
            .I(N__92770));
    SRMux I__22646 (
            .O(N__92977),
            .I(N__92770));
    SRMux I__22645 (
            .O(N__92976),
            .I(N__92770));
    SRMux I__22644 (
            .O(N__92975),
            .I(N__92770));
    SRMux I__22643 (
            .O(N__92974),
            .I(N__92770));
    SRMux I__22642 (
            .O(N__92973),
            .I(N__92770));
    SRMux I__22641 (
            .O(N__92972),
            .I(N__92770));
    SRMux I__22640 (
            .O(N__92971),
            .I(N__92770));
    SRMux I__22639 (
            .O(N__92970),
            .I(N__92770));
    SRMux I__22638 (
            .O(N__92969),
            .I(N__92770));
    SRMux I__22637 (
            .O(N__92968),
            .I(N__92770));
    SRMux I__22636 (
            .O(N__92967),
            .I(N__92770));
    SRMux I__22635 (
            .O(N__92966),
            .I(N__92770));
    SRMux I__22634 (
            .O(N__92965),
            .I(N__92770));
    Glb2LocalMux I__22633 (
            .O(N__92962),
            .I(N__92770));
    Glb2LocalMux I__22632 (
            .O(N__92959),
            .I(N__92770));
    Glb2LocalMux I__22631 (
            .O(N__92956),
            .I(N__92770));
    Glb2LocalMux I__22630 (
            .O(N__92953),
            .I(N__92770));
    Glb2LocalMux I__22629 (
            .O(N__92950),
            .I(N__92770));
    Glb2LocalMux I__22628 (
            .O(N__92947),
            .I(N__92770));
    Glb2LocalMux I__22627 (
            .O(N__92944),
            .I(N__92770));
    Glb2LocalMux I__22626 (
            .O(N__92941),
            .I(N__92770));
    Glb2LocalMux I__22625 (
            .O(N__92938),
            .I(N__92770));
    Glb2LocalMux I__22624 (
            .O(N__92935),
            .I(N__92770));
    Glb2LocalMux I__22623 (
            .O(N__92932),
            .I(N__92770));
    Glb2LocalMux I__22622 (
            .O(N__92929),
            .I(N__92770));
    Glb2LocalMux I__22621 (
            .O(N__92926),
            .I(N__92770));
    Glb2LocalMux I__22620 (
            .O(N__92923),
            .I(N__92770));
    Glb2LocalMux I__22619 (
            .O(N__92920),
            .I(N__92770));
    Glb2LocalMux I__22618 (
            .O(N__92917),
            .I(N__92770));
    Glb2LocalMux I__22617 (
            .O(N__92914),
            .I(N__92770));
    Glb2LocalMux I__22616 (
            .O(N__92911),
            .I(N__92770));
    GlobalMux I__22615 (
            .O(N__92770),
            .I(N__92767));
    gio2CtrlBuf I__22614 (
            .O(N__92767),
            .I(N_934_g));
    InMux I__22613 (
            .O(N__92764),
            .I(N__92761));
    LocalMux I__22612 (
            .O(N__92761),
            .I(N__92758));
    Odrv4 I__22611 (
            .O(N__92758),
            .I(\pid_side.O_1_21 ));
    InMux I__22610 (
            .O(N__92755),
            .I(N__92751));
    InMux I__22609 (
            .O(N__92754),
            .I(N__92748));
    LocalMux I__22608 (
            .O(N__92751),
            .I(N__92744));
    LocalMux I__22607 (
            .O(N__92748),
            .I(N__92741));
    InMux I__22606 (
            .O(N__92747),
            .I(N__92738));
    Span4Mux_v I__22605 (
            .O(N__92744),
            .I(N__92733));
    Span4Mux_h I__22604 (
            .O(N__92741),
            .I(N__92733));
    LocalMux I__22603 (
            .O(N__92738),
            .I(N__92730));
    Span4Mux_v I__22602 (
            .O(N__92733),
            .I(N__92727));
    Span4Mux_v I__22601 (
            .O(N__92730),
            .I(N__92724));
    Odrv4 I__22600 (
            .O(N__92727),
            .I(\pid_side.error_d_regZ0Z_18 ));
    Odrv4 I__22599 (
            .O(N__92724),
            .I(\pid_side.error_d_regZ0Z_18 ));
    InMux I__22598 (
            .O(N__92719),
            .I(N__92716));
    LocalMux I__22597 (
            .O(N__92716),
            .I(N__92713));
    Odrv4 I__22596 (
            .O(N__92713),
            .I(\pid_side.O_1_19 ));
    InMux I__22595 (
            .O(N__92710),
            .I(N__92701));
    InMux I__22594 (
            .O(N__92709),
            .I(N__92701));
    InMux I__22593 (
            .O(N__92708),
            .I(N__92701));
    LocalMux I__22592 (
            .O(N__92701),
            .I(N__92698));
    Span4Mux_h I__22591 (
            .O(N__92698),
            .I(N__92695));
    Span4Mux_v I__22590 (
            .O(N__92695),
            .I(N__92692));
    Span4Mux_v I__22589 (
            .O(N__92692),
            .I(N__92689));
    Span4Mux_h I__22588 (
            .O(N__92689),
            .I(N__92686));
    Odrv4 I__22587 (
            .O(N__92686),
            .I(\pid_side.error_d_regZ0Z_16 ));
    CEMux I__22586 (
            .O(N__92683),
            .I(N__92679));
    CEMux I__22585 (
            .O(N__92682),
            .I(N__92673));
    LocalMux I__22584 (
            .O(N__92679),
            .I(N__92669));
    CEMux I__22583 (
            .O(N__92678),
            .I(N__92666));
    CEMux I__22582 (
            .O(N__92677),
            .I(N__92662));
    CEMux I__22581 (
            .O(N__92676),
            .I(N__92658));
    LocalMux I__22580 (
            .O(N__92673),
            .I(N__92652));
    CEMux I__22579 (
            .O(N__92672),
            .I(N__92646));
    Span4Mux_s3_h I__22578 (
            .O(N__92669),
            .I(N__92641));
    LocalMux I__22577 (
            .O(N__92666),
            .I(N__92641));
    CEMux I__22576 (
            .O(N__92665),
            .I(N__92638));
    LocalMux I__22575 (
            .O(N__92662),
            .I(N__92635));
    CEMux I__22574 (
            .O(N__92661),
            .I(N__92632));
    LocalMux I__22573 (
            .O(N__92658),
            .I(N__92629));
    CEMux I__22572 (
            .O(N__92657),
            .I(N__92626));
    CEMux I__22571 (
            .O(N__92656),
            .I(N__92623));
    CEMux I__22570 (
            .O(N__92655),
            .I(N__92620));
    Span4Mux_s3_h I__22569 (
            .O(N__92652),
            .I(N__92616));
    CEMux I__22568 (
            .O(N__92651),
            .I(N__92613));
    CEMux I__22567 (
            .O(N__92650),
            .I(N__92610));
    CEMux I__22566 (
            .O(N__92649),
            .I(N__92607));
    LocalMux I__22565 (
            .O(N__92646),
            .I(N__92604));
    Span4Mux_v I__22564 (
            .O(N__92641),
            .I(N__92601));
    LocalMux I__22563 (
            .O(N__92638),
            .I(N__92598));
    Span4Mux_v I__22562 (
            .O(N__92635),
            .I(N__92591));
    LocalMux I__22561 (
            .O(N__92632),
            .I(N__92591));
    Span4Mux_v I__22560 (
            .O(N__92629),
            .I(N__92591));
    LocalMux I__22559 (
            .O(N__92626),
            .I(N__92586));
    LocalMux I__22558 (
            .O(N__92623),
            .I(N__92586));
    LocalMux I__22557 (
            .O(N__92620),
            .I(N__92583));
    CEMux I__22556 (
            .O(N__92619),
            .I(N__92580));
    Span4Mux_h I__22555 (
            .O(N__92616),
            .I(N__92577));
    LocalMux I__22554 (
            .O(N__92613),
            .I(N__92574));
    LocalMux I__22553 (
            .O(N__92610),
            .I(N__92567));
    LocalMux I__22552 (
            .O(N__92607),
            .I(N__92567));
    Sp12to4 I__22551 (
            .O(N__92604),
            .I(N__92567));
    Span4Mux_s3_h I__22550 (
            .O(N__92601),
            .I(N__92564));
    Span4Mux_s3_h I__22549 (
            .O(N__92598),
            .I(N__92561));
    Span4Mux_h I__22548 (
            .O(N__92591),
            .I(N__92552));
    Span4Mux_v I__22547 (
            .O(N__92586),
            .I(N__92552));
    Span4Mux_v I__22546 (
            .O(N__92583),
            .I(N__92552));
    LocalMux I__22545 (
            .O(N__92580),
            .I(N__92552));
    Sp12to4 I__22544 (
            .O(N__92577),
            .I(N__92545));
    Sp12to4 I__22543 (
            .O(N__92574),
            .I(N__92545));
    Span12Mux_v I__22542 (
            .O(N__92567),
            .I(N__92545));
    Span4Mux_h I__22541 (
            .O(N__92564),
            .I(N__92540));
    Span4Mux_h I__22540 (
            .O(N__92561),
            .I(N__92540));
    Span4Mux_h I__22539 (
            .O(N__92552),
            .I(N__92537));
    Span12Mux_h I__22538 (
            .O(N__92545),
            .I(N__92534));
    Span4Mux_h I__22537 (
            .O(N__92540),
            .I(N__92531));
    Span4Mux_h I__22536 (
            .O(N__92537),
            .I(N__92528));
    Odrv12 I__22535 (
            .O(N__92534),
            .I(\pid_side.N_868_0 ));
    Odrv4 I__22534 (
            .O(N__92531),
            .I(\pid_side.N_868_0 ));
    Odrv4 I__22533 (
            .O(N__92528),
            .I(\pid_side.N_868_0 ));
    InMux I__22532 (
            .O(N__92521),
            .I(N__92510));
    InMux I__22531 (
            .O(N__92520),
            .I(N__92506));
    InMux I__22530 (
            .O(N__92519),
            .I(N__92503));
    InMux I__22529 (
            .O(N__92518),
            .I(N__92500));
    InMux I__22528 (
            .O(N__92517),
            .I(N__92495));
    InMux I__22527 (
            .O(N__92516),
            .I(N__92495));
    InMux I__22526 (
            .O(N__92515),
            .I(N__92491));
    InMux I__22525 (
            .O(N__92514),
            .I(N__92488));
    InMux I__22524 (
            .O(N__92513),
            .I(N__92485));
    LocalMux I__22523 (
            .O(N__92510),
            .I(N__92482));
    InMux I__22522 (
            .O(N__92509),
            .I(N__92479));
    LocalMux I__22521 (
            .O(N__92506),
            .I(N__92476));
    LocalMux I__22520 (
            .O(N__92503),
            .I(N__92471));
    LocalMux I__22519 (
            .O(N__92500),
            .I(N__92466));
    LocalMux I__22518 (
            .O(N__92495),
            .I(N__92466));
    InMux I__22517 (
            .O(N__92494),
            .I(N__92462));
    LocalMux I__22516 (
            .O(N__92491),
            .I(N__92459));
    LocalMux I__22515 (
            .O(N__92488),
            .I(N__92454));
    LocalMux I__22514 (
            .O(N__92485),
            .I(N__92454));
    Span4Mux_h I__22513 (
            .O(N__92482),
            .I(N__92451));
    LocalMux I__22512 (
            .O(N__92479),
            .I(N__92448));
    Span4Mux_v I__22511 (
            .O(N__92476),
            .I(N__92445));
    InMux I__22510 (
            .O(N__92475),
            .I(N__92442));
    InMux I__22509 (
            .O(N__92474),
            .I(N__92439));
    Span4Mux_v I__22508 (
            .O(N__92471),
            .I(N__92436));
    Span4Mux_v I__22507 (
            .O(N__92466),
            .I(N__92433));
    InMux I__22506 (
            .O(N__92465),
            .I(N__92427));
    LocalMux I__22505 (
            .O(N__92462),
            .I(N__92420));
    Span4Mux_v I__22504 (
            .O(N__92459),
            .I(N__92420));
    Span4Mux_h I__22503 (
            .O(N__92454),
            .I(N__92420));
    Span4Mux_v I__22502 (
            .O(N__92451),
            .I(N__92417));
    Span4Mux_v I__22501 (
            .O(N__92448),
            .I(N__92414));
    Span4Mux_v I__22500 (
            .O(N__92445),
            .I(N__92411));
    LocalMux I__22499 (
            .O(N__92442),
            .I(N__92408));
    LocalMux I__22498 (
            .O(N__92439),
            .I(N__92405));
    Sp12to4 I__22497 (
            .O(N__92436),
            .I(N__92400));
    Sp12to4 I__22496 (
            .O(N__92433),
            .I(N__92400));
    InMux I__22495 (
            .O(N__92432),
            .I(N__92393));
    InMux I__22494 (
            .O(N__92431),
            .I(N__92393));
    InMux I__22493 (
            .O(N__92430),
            .I(N__92393));
    LocalMux I__22492 (
            .O(N__92427),
            .I(N__92384));
    Span4Mux_h I__22491 (
            .O(N__92420),
            .I(N__92384));
    Span4Mux_h I__22490 (
            .O(N__92417),
            .I(N__92384));
    Span4Mux_v I__22489 (
            .O(N__92414),
            .I(N__92377));
    Span4Mux_h I__22488 (
            .O(N__92411),
            .I(N__92377));
    Span4Mux_v I__22487 (
            .O(N__92408),
            .I(N__92377));
    Span12Mux_v I__22486 (
            .O(N__92405),
            .I(N__92370));
    Span12Mux_s8_h I__22485 (
            .O(N__92400),
            .I(N__92370));
    LocalMux I__22484 (
            .O(N__92393),
            .I(N__92370));
    InMux I__22483 (
            .O(N__92392),
            .I(N__92365));
    InMux I__22482 (
            .O(N__92391),
            .I(N__92365));
    Odrv4 I__22481 (
            .O(N__92384),
            .I(uart_pc_data_2));
    Odrv4 I__22480 (
            .O(N__92377),
            .I(uart_pc_data_2));
    Odrv12 I__22479 (
            .O(N__92370),
            .I(uart_pc_data_2));
    LocalMux I__22478 (
            .O(N__92365),
            .I(uart_pc_data_2));
    InMux I__22477 (
            .O(N__92356),
            .I(N__92352));
    InMux I__22476 (
            .O(N__92355),
            .I(N__92349));
    LocalMux I__22475 (
            .O(N__92352),
            .I(N__92346));
    LocalMux I__22474 (
            .O(N__92349),
            .I(N__92343));
    Span4Mux_s1_h I__22473 (
            .O(N__92346),
            .I(N__92340));
    Span4Mux_v I__22472 (
            .O(N__92343),
            .I(N__92337));
    Odrv4 I__22471 (
            .O(N__92340),
            .I(xy_kd_2));
    Odrv4 I__22470 (
            .O(N__92337),
            .I(xy_kd_2));
    InMux I__22469 (
            .O(N__92332),
            .I(N__92323));
    InMux I__22468 (
            .O(N__92331),
            .I(N__92316));
    InMux I__22467 (
            .O(N__92330),
            .I(N__92313));
    InMux I__22466 (
            .O(N__92329),
            .I(N__92308));
    InMux I__22465 (
            .O(N__92328),
            .I(N__92308));
    InMux I__22464 (
            .O(N__92327),
            .I(N__92305));
    InMux I__22463 (
            .O(N__92326),
            .I(N__92302));
    LocalMux I__22462 (
            .O(N__92323),
            .I(N__92298));
    InMux I__22461 (
            .O(N__92322),
            .I(N__92295));
    InMux I__22460 (
            .O(N__92321),
            .I(N__92288));
    InMux I__22459 (
            .O(N__92320),
            .I(N__92288));
    InMux I__22458 (
            .O(N__92319),
            .I(N__92288));
    LocalMux I__22457 (
            .O(N__92316),
            .I(N__92284));
    LocalMux I__22456 (
            .O(N__92313),
            .I(N__92280));
    LocalMux I__22455 (
            .O(N__92308),
            .I(N__92276));
    LocalMux I__22454 (
            .O(N__92305),
            .I(N__92273));
    LocalMux I__22453 (
            .O(N__92302),
            .I(N__92270));
    InMux I__22452 (
            .O(N__92301),
            .I(N__92267));
    Span4Mux_h I__22451 (
            .O(N__92298),
            .I(N__92264));
    LocalMux I__22450 (
            .O(N__92295),
            .I(N__92259));
    LocalMux I__22449 (
            .O(N__92288),
            .I(N__92259));
    InMux I__22448 (
            .O(N__92287),
            .I(N__92256));
    Span4Mux_h I__22447 (
            .O(N__92284),
            .I(N__92253));
    InMux I__22446 (
            .O(N__92283),
            .I(N__92250));
    Span4Mux_h I__22445 (
            .O(N__92280),
            .I(N__92247));
    InMux I__22444 (
            .O(N__92279),
            .I(N__92244));
    Span4Mux_v I__22443 (
            .O(N__92276),
            .I(N__92239));
    Span4Mux_h I__22442 (
            .O(N__92273),
            .I(N__92239));
    Span4Mux_h I__22441 (
            .O(N__92270),
            .I(N__92236));
    LocalMux I__22440 (
            .O(N__92267),
            .I(N__92231));
    Sp12to4 I__22439 (
            .O(N__92264),
            .I(N__92228));
    Span4Mux_v I__22438 (
            .O(N__92259),
            .I(N__92225));
    LocalMux I__22437 (
            .O(N__92256),
            .I(N__92222));
    Span4Mux_h I__22436 (
            .O(N__92253),
            .I(N__92219));
    LocalMux I__22435 (
            .O(N__92250),
            .I(N__92216));
    Span4Mux_v I__22434 (
            .O(N__92247),
            .I(N__92213));
    LocalMux I__22433 (
            .O(N__92244),
            .I(N__92208));
    Span4Mux_h I__22432 (
            .O(N__92239),
            .I(N__92208));
    Span4Mux_v I__22431 (
            .O(N__92236),
            .I(N__92205));
    InMux I__22430 (
            .O(N__92235),
            .I(N__92200));
    InMux I__22429 (
            .O(N__92234),
            .I(N__92200));
    Span12Mux_v I__22428 (
            .O(N__92231),
            .I(N__92193));
    Span12Mux_v I__22427 (
            .O(N__92228),
            .I(N__92193));
    Sp12to4 I__22426 (
            .O(N__92225),
            .I(N__92193));
    Span4Mux_h I__22425 (
            .O(N__92222),
            .I(N__92188));
    Sp12to4 I__22424 (
            .O(N__92219),
            .I(N__92183));
    Span12Mux_s11_v I__22423 (
            .O(N__92216),
            .I(N__92183));
    Span4Mux_h I__22422 (
            .O(N__92213),
            .I(N__92178));
    Span4Mux_h I__22421 (
            .O(N__92208),
            .I(N__92178));
    Span4Mux_v I__22420 (
            .O(N__92205),
            .I(N__92173));
    LocalMux I__22419 (
            .O(N__92200),
            .I(N__92173));
    Span12Mux_h I__22418 (
            .O(N__92193),
            .I(N__92170));
    InMux I__22417 (
            .O(N__92192),
            .I(N__92165));
    InMux I__22416 (
            .O(N__92191),
            .I(N__92165));
    Odrv4 I__22415 (
            .O(N__92188),
            .I(uart_pc_data_3));
    Odrv12 I__22414 (
            .O(N__92183),
            .I(uart_pc_data_3));
    Odrv4 I__22413 (
            .O(N__92178),
            .I(uart_pc_data_3));
    Odrv4 I__22412 (
            .O(N__92173),
            .I(uart_pc_data_3));
    Odrv12 I__22411 (
            .O(N__92170),
            .I(uart_pc_data_3));
    LocalMux I__22410 (
            .O(N__92165),
            .I(uart_pc_data_3));
    InMux I__22409 (
            .O(N__92152),
            .I(N__92148));
    InMux I__22408 (
            .O(N__92151),
            .I(N__92145));
    LocalMux I__22407 (
            .O(N__92148),
            .I(N__92142));
    LocalMux I__22406 (
            .O(N__92145),
            .I(N__92139));
    Span4Mux_v I__22405 (
            .O(N__92142),
            .I(N__92134));
    Span4Mux_v I__22404 (
            .O(N__92139),
            .I(N__92134));
    Odrv4 I__22403 (
            .O(N__92134),
            .I(xy_kd_3));
    InMux I__22402 (
            .O(N__92131),
            .I(N__92128));
    LocalMux I__22401 (
            .O(N__92128),
            .I(N__92119));
    InMux I__22400 (
            .O(N__92127),
            .I(N__92116));
    InMux I__22399 (
            .O(N__92126),
            .I(N__92113));
    InMux I__22398 (
            .O(N__92125),
            .I(N__92110));
    InMux I__22397 (
            .O(N__92124),
            .I(N__92107));
    InMux I__22396 (
            .O(N__92123),
            .I(N__92104));
    InMux I__22395 (
            .O(N__92122),
            .I(N__92098));
    Span4Mux_v I__22394 (
            .O(N__92119),
            .I(N__92093));
    LocalMux I__22393 (
            .O(N__92116),
            .I(N__92093));
    LocalMux I__22392 (
            .O(N__92113),
            .I(N__92090));
    LocalMux I__22391 (
            .O(N__92110),
            .I(N__92087));
    LocalMux I__22390 (
            .O(N__92107),
            .I(N__92084));
    LocalMux I__22389 (
            .O(N__92104),
            .I(N__92081));
    InMux I__22388 (
            .O(N__92103),
            .I(N__92078));
    CascadeMux I__22387 (
            .O(N__92102),
            .I(N__92075));
    CascadeMux I__22386 (
            .O(N__92101),
            .I(N__92072));
    LocalMux I__22385 (
            .O(N__92098),
            .I(N__92067));
    Span4Mux_h I__22384 (
            .O(N__92093),
            .I(N__92062));
    Span4Mux_v I__22383 (
            .O(N__92090),
            .I(N__92059));
    Span4Mux_v I__22382 (
            .O(N__92087),
            .I(N__92056));
    Span4Mux_h I__22381 (
            .O(N__92084),
            .I(N__92053));
    Span4Mux_v I__22380 (
            .O(N__92081),
            .I(N__92047));
    LocalMux I__22379 (
            .O(N__92078),
            .I(N__92047));
    InMux I__22378 (
            .O(N__92075),
            .I(N__92042));
    InMux I__22377 (
            .O(N__92072),
            .I(N__92042));
    InMux I__22376 (
            .O(N__92071),
            .I(N__92038));
    InMux I__22375 (
            .O(N__92070),
            .I(N__92035));
    Span4Mux_v I__22374 (
            .O(N__92067),
            .I(N__92032));
    InMux I__22373 (
            .O(N__92066),
            .I(N__92029));
    InMux I__22372 (
            .O(N__92065),
            .I(N__92026));
    Sp12to4 I__22371 (
            .O(N__92062),
            .I(N__92023));
    Sp12to4 I__22370 (
            .O(N__92059),
            .I(N__92018));
    Sp12to4 I__22369 (
            .O(N__92056),
            .I(N__92018));
    Sp12to4 I__22368 (
            .O(N__92053),
            .I(N__92015));
    InMux I__22367 (
            .O(N__92052),
            .I(N__92012));
    Span4Mux_h I__22366 (
            .O(N__92047),
            .I(N__92009));
    LocalMux I__22365 (
            .O(N__92042),
            .I(N__92006));
    InMux I__22364 (
            .O(N__92041),
            .I(N__92003));
    LocalMux I__22363 (
            .O(N__92038),
            .I(N__92000));
    LocalMux I__22362 (
            .O(N__92035),
            .I(N__91997));
    Span4Mux_h I__22361 (
            .O(N__92032),
            .I(N__91992));
    LocalMux I__22360 (
            .O(N__92029),
            .I(N__91992));
    LocalMux I__22359 (
            .O(N__92026),
            .I(N__91989));
    Span12Mux_v I__22358 (
            .O(N__92023),
            .I(N__91982));
    Span12Mux_s9_h I__22357 (
            .O(N__92018),
            .I(N__91982));
    Span12Mux_v I__22356 (
            .O(N__92015),
            .I(N__91982));
    LocalMux I__22355 (
            .O(N__92012),
            .I(N__91973));
    Span4Mux_v I__22354 (
            .O(N__92009),
            .I(N__91973));
    Span4Mux_h I__22353 (
            .O(N__92006),
            .I(N__91973));
    LocalMux I__22352 (
            .O(N__92003),
            .I(N__91973));
    Span4Mux_v I__22351 (
            .O(N__92000),
            .I(N__91966));
    Span4Mux_h I__22350 (
            .O(N__91997),
            .I(N__91966));
    Span4Mux_v I__22349 (
            .O(N__91992),
            .I(N__91966));
    Odrv12 I__22348 (
            .O(N__91989),
            .I(uart_pc_data_7));
    Odrv12 I__22347 (
            .O(N__91982),
            .I(uart_pc_data_7));
    Odrv4 I__22346 (
            .O(N__91973),
            .I(uart_pc_data_7));
    Odrv4 I__22345 (
            .O(N__91966),
            .I(uart_pc_data_7));
    InMux I__22344 (
            .O(N__91957),
            .I(N__91953));
    InMux I__22343 (
            .O(N__91956),
            .I(N__91950));
    LocalMux I__22342 (
            .O(N__91953),
            .I(N__91947));
    LocalMux I__22341 (
            .O(N__91950),
            .I(N__91944));
    Span4Mux_v I__22340 (
            .O(N__91947),
            .I(N__91939));
    Span4Mux_v I__22339 (
            .O(N__91944),
            .I(N__91939));
    Odrv4 I__22338 (
            .O(N__91939),
            .I(xy_kd_7));
    CEMux I__22337 (
            .O(N__91936),
            .I(N__91933));
    LocalMux I__22336 (
            .O(N__91933),
            .I(N__91929));
    CEMux I__22335 (
            .O(N__91932),
            .I(N__91925));
    Span4Mux_v I__22334 (
            .O(N__91929),
            .I(N__91921));
    CEMux I__22333 (
            .O(N__91928),
            .I(N__91918));
    LocalMux I__22332 (
            .O(N__91925),
            .I(N__91914));
    CEMux I__22331 (
            .O(N__91924),
            .I(N__91911));
    Span4Mux_h I__22330 (
            .O(N__91921),
            .I(N__91908));
    LocalMux I__22329 (
            .O(N__91918),
            .I(N__91905));
    CEMux I__22328 (
            .O(N__91917),
            .I(N__91902));
    Span4Mux_s2_h I__22327 (
            .O(N__91914),
            .I(N__91897));
    LocalMux I__22326 (
            .O(N__91911),
            .I(N__91897));
    Span4Mux_h I__22325 (
            .O(N__91908),
            .I(N__91892));
    Span4Mux_h I__22324 (
            .O(N__91905),
            .I(N__91892));
    LocalMux I__22323 (
            .O(N__91902),
            .I(N__91889));
    Span4Mux_h I__22322 (
            .O(N__91897),
            .I(N__91886));
    Span4Mux_h I__22321 (
            .O(N__91892),
            .I(N__91883));
    Span12Mux_v I__22320 (
            .O(N__91889),
            .I(N__91878));
    Sp12to4 I__22319 (
            .O(N__91886),
            .I(N__91878));
    Span4Mux_h I__22318 (
            .O(N__91883),
            .I(N__91875));
    Odrv12 I__22317 (
            .O(N__91878),
            .I(\Commands_frame_decoder.state_RNITUI31Z0Z_13 ));
    Odrv4 I__22316 (
            .O(N__91875),
            .I(\Commands_frame_decoder.state_RNITUI31Z0Z_13 ));
    InMux I__22315 (
            .O(N__91870),
            .I(N__91867));
    LocalMux I__22314 (
            .O(N__91867),
            .I(N__91864));
    Span4Mux_h I__22313 (
            .O(N__91864),
            .I(N__91861));
    Odrv4 I__22312 (
            .O(N__91861),
            .I(\pid_front.O_23 ));
    InMux I__22311 (
            .O(N__91858),
            .I(N__91853));
    InMux I__22310 (
            .O(N__91857),
            .I(N__91848));
    InMux I__22309 (
            .O(N__91856),
            .I(N__91848));
    LocalMux I__22308 (
            .O(N__91853),
            .I(N__91845));
    LocalMux I__22307 (
            .O(N__91848),
            .I(N__91842));
    Span4Mux_v I__22306 (
            .O(N__91845),
            .I(N__91837));
    Span4Mux_v I__22305 (
            .O(N__91842),
            .I(N__91837));
    Span4Mux_h I__22304 (
            .O(N__91837),
            .I(N__91834));
    Span4Mux_h I__22303 (
            .O(N__91834),
            .I(N__91831));
    Odrv4 I__22302 (
            .O(N__91831),
            .I(\pid_front.error_d_regZ0Z_20 ));
    InMux I__22301 (
            .O(N__91828),
            .I(N__91825));
    LocalMux I__22300 (
            .O(N__91825),
            .I(N__91822));
    Span4Mux_v I__22299 (
            .O(N__91822),
            .I(N__91819));
    Odrv4 I__22298 (
            .O(N__91819),
            .I(\pid_front.O_22 ));
    InMux I__22297 (
            .O(N__91816),
            .I(N__91813));
    LocalMux I__22296 (
            .O(N__91813),
            .I(N__91808));
    InMux I__22295 (
            .O(N__91812),
            .I(N__91803));
    InMux I__22294 (
            .O(N__91811),
            .I(N__91803));
    Span4Mux_v I__22293 (
            .O(N__91808),
            .I(N__91798));
    LocalMux I__22292 (
            .O(N__91803),
            .I(N__91798));
    Span4Mux_h I__22291 (
            .O(N__91798),
            .I(N__91795));
    Span4Mux_h I__22290 (
            .O(N__91795),
            .I(N__91792));
    Odrv4 I__22289 (
            .O(N__91792),
            .I(\pid_front.error_d_regZ0Z_19 ));
    InMux I__22288 (
            .O(N__91789),
            .I(N__91786));
    LocalMux I__22287 (
            .O(N__91786),
            .I(N__91783));
    Odrv4 I__22286 (
            .O(N__91783),
            .I(\pid_front.O_24 ));
    CascadeMux I__22285 (
            .O(N__91780),
            .I(N__91776));
    InMux I__22284 (
            .O(N__91779),
            .I(N__91766));
    InMux I__22283 (
            .O(N__91776),
            .I(N__91766));
    InMux I__22282 (
            .O(N__91775),
            .I(N__91766));
    InMux I__22281 (
            .O(N__91774),
            .I(N__91763));
    CascadeMux I__22280 (
            .O(N__91773),
            .I(N__91760));
    LocalMux I__22279 (
            .O(N__91766),
            .I(N__91751));
    LocalMux I__22278 (
            .O(N__91763),
            .I(N__91748));
    InMux I__22277 (
            .O(N__91760),
            .I(N__91741));
    InMux I__22276 (
            .O(N__91759),
            .I(N__91741));
    InMux I__22275 (
            .O(N__91758),
            .I(N__91741));
    InMux I__22274 (
            .O(N__91757),
            .I(N__91737));
    CascadeMux I__22273 (
            .O(N__91756),
            .I(N__91734));
    CascadeMux I__22272 (
            .O(N__91755),
            .I(N__91731));
    InMux I__22271 (
            .O(N__91754),
            .I(N__91727));
    Span4Mux_h I__22270 (
            .O(N__91751),
            .I(N__91720));
    Span4Mux_s3_v I__22269 (
            .O(N__91748),
            .I(N__91720));
    LocalMux I__22268 (
            .O(N__91741),
            .I(N__91720));
    InMux I__22267 (
            .O(N__91740),
            .I(N__91714));
    LocalMux I__22266 (
            .O(N__91737),
            .I(N__91711));
    InMux I__22265 (
            .O(N__91734),
            .I(N__91704));
    InMux I__22264 (
            .O(N__91731),
            .I(N__91704));
    InMux I__22263 (
            .O(N__91730),
            .I(N__91704));
    LocalMux I__22262 (
            .O(N__91727),
            .I(N__91699));
    Span4Mux_v I__22261 (
            .O(N__91720),
            .I(N__91699));
    InMux I__22260 (
            .O(N__91719),
            .I(N__91692));
    InMux I__22259 (
            .O(N__91718),
            .I(N__91692));
    InMux I__22258 (
            .O(N__91717),
            .I(N__91692));
    LocalMux I__22257 (
            .O(N__91714),
            .I(N__91685));
    Span4Mux_v I__22256 (
            .O(N__91711),
            .I(N__91685));
    LocalMux I__22255 (
            .O(N__91704),
            .I(N__91685));
    Span4Mux_h I__22254 (
            .O(N__91699),
            .I(N__91682));
    LocalMux I__22253 (
            .O(N__91692),
            .I(N__91679));
    Span4Mux_h I__22252 (
            .O(N__91685),
            .I(N__91676));
    Span4Mux_h I__22251 (
            .O(N__91682),
            .I(N__91673));
    Span12Mux_h I__22250 (
            .O(N__91679),
            .I(N__91670));
    Span4Mux_h I__22249 (
            .O(N__91676),
            .I(N__91667));
    Odrv4 I__22248 (
            .O(N__91673),
            .I(\pid_front.error_d_regZ0Z_21 ));
    Odrv12 I__22247 (
            .O(N__91670),
            .I(\pid_front.error_d_regZ0Z_21 ));
    Odrv4 I__22246 (
            .O(N__91667),
            .I(\pid_front.error_d_regZ0Z_21 ));
    InMux I__22245 (
            .O(N__91660),
            .I(N__91657));
    LocalMux I__22244 (
            .O(N__91657),
            .I(N__91654));
    Odrv4 I__22243 (
            .O(N__91654),
            .I(\pid_side.O_2_24 ));
    InMux I__22242 (
            .O(N__91651),
            .I(N__91632));
    InMux I__22241 (
            .O(N__91650),
            .I(N__91632));
    InMux I__22240 (
            .O(N__91649),
            .I(N__91632));
    InMux I__22239 (
            .O(N__91648),
            .I(N__91627));
    InMux I__22238 (
            .O(N__91647),
            .I(N__91627));
    InMux I__22237 (
            .O(N__91646),
            .I(N__91622));
    InMux I__22236 (
            .O(N__91645),
            .I(N__91613));
    InMux I__22235 (
            .O(N__91644),
            .I(N__91613));
    InMux I__22234 (
            .O(N__91643),
            .I(N__91613));
    InMux I__22233 (
            .O(N__91642),
            .I(N__91613));
    InMux I__22232 (
            .O(N__91641),
            .I(N__91606));
    InMux I__22231 (
            .O(N__91640),
            .I(N__91606));
    InMux I__22230 (
            .O(N__91639),
            .I(N__91606));
    LocalMux I__22229 (
            .O(N__91632),
            .I(N__91601));
    LocalMux I__22228 (
            .O(N__91627),
            .I(N__91601));
    InMux I__22227 (
            .O(N__91626),
            .I(N__91596));
    InMux I__22226 (
            .O(N__91625),
            .I(N__91596));
    LocalMux I__22225 (
            .O(N__91622),
            .I(N__91591));
    LocalMux I__22224 (
            .O(N__91613),
            .I(N__91588));
    LocalMux I__22223 (
            .O(N__91606),
            .I(N__91581));
    Span4Mux_h I__22222 (
            .O(N__91601),
            .I(N__91581));
    LocalMux I__22221 (
            .O(N__91596),
            .I(N__91581));
    InMux I__22220 (
            .O(N__91595),
            .I(N__91576));
    InMux I__22219 (
            .O(N__91594),
            .I(N__91576));
    Span4Mux_v I__22218 (
            .O(N__91591),
            .I(N__91571));
    Span4Mux_h I__22217 (
            .O(N__91588),
            .I(N__91571));
    Span4Mux_v I__22216 (
            .O(N__91581),
            .I(N__91568));
    LocalMux I__22215 (
            .O(N__91576),
            .I(N__91565));
    Span4Mux_h I__22214 (
            .O(N__91571),
            .I(N__91560));
    Span4Mux_h I__22213 (
            .O(N__91568),
            .I(N__91560));
    Span12Mux_h I__22212 (
            .O(N__91565),
            .I(N__91557));
    Odrv4 I__22211 (
            .O(N__91560),
            .I(\pid_side.error_p_regZ0Z_20 ));
    Odrv12 I__22210 (
            .O(N__91557),
            .I(\pid_side.error_p_regZ0Z_20 ));
    InMux I__22209 (
            .O(N__91552),
            .I(N__91549));
    LocalMux I__22208 (
            .O(N__91549),
            .I(N__91546));
    Span4Mux_h I__22207 (
            .O(N__91546),
            .I(N__91543));
    Odrv4 I__22206 (
            .O(N__91543),
            .I(\pid_side.O_1_18 ));
    InMux I__22205 (
            .O(N__91540),
            .I(N__91531));
    InMux I__22204 (
            .O(N__91539),
            .I(N__91531));
    InMux I__22203 (
            .O(N__91538),
            .I(N__91531));
    LocalMux I__22202 (
            .O(N__91531),
            .I(N__91528));
    Span12Mux_v I__22201 (
            .O(N__91528),
            .I(N__91525));
    Odrv12 I__22200 (
            .O(N__91525),
            .I(\pid_side.error_d_regZ0Z_15 ));
    InMux I__22199 (
            .O(N__91522),
            .I(N__91519));
    LocalMux I__22198 (
            .O(N__91519),
            .I(N__91515));
    InMux I__22197 (
            .O(N__91518),
            .I(N__91512));
    Span4Mux_h I__22196 (
            .O(N__91515),
            .I(N__91509));
    LocalMux I__22195 (
            .O(N__91512),
            .I(N__91506));
    Span4Mux_v I__22194 (
            .O(N__91509),
            .I(N__91503));
    Span4Mux_h I__22193 (
            .O(N__91506),
            .I(N__91500));
    Odrv4 I__22192 (
            .O(N__91503),
            .I(\pid_side.O_1_16 ));
    Odrv4 I__22191 (
            .O(N__91500),
            .I(\pid_side.O_1_16 ));
    InMux I__22190 (
            .O(N__91495),
            .I(N__91489));
    InMux I__22189 (
            .O(N__91494),
            .I(N__91489));
    LocalMux I__22188 (
            .O(N__91489),
            .I(N__91485));
    InMux I__22187 (
            .O(N__91488),
            .I(N__91478));
    Span4Mux_h I__22186 (
            .O(N__91485),
            .I(N__91475));
    InMux I__22185 (
            .O(N__91484),
            .I(N__91466));
    InMux I__22184 (
            .O(N__91483),
            .I(N__91466));
    InMux I__22183 (
            .O(N__91482),
            .I(N__91466));
    InMux I__22182 (
            .O(N__91481),
            .I(N__91466));
    LocalMux I__22181 (
            .O(N__91478),
            .I(N__91459));
    Span4Mux_h I__22180 (
            .O(N__91475),
            .I(N__91459));
    LocalMux I__22179 (
            .O(N__91466),
            .I(N__91459));
    Span4Mux_h I__22178 (
            .O(N__91459),
            .I(N__91456));
    Odrv4 I__22177 (
            .O(N__91456),
            .I(\pid_side.error_d_regZ0Z_13 ));
    InMux I__22176 (
            .O(N__91453),
            .I(N__91450));
    LocalMux I__22175 (
            .O(N__91450),
            .I(N__91447));
    Span4Mux_h I__22174 (
            .O(N__91447),
            .I(N__91444));
    Odrv4 I__22173 (
            .O(N__91444),
            .I(\pid_side.O_1_17 ));
    InMux I__22172 (
            .O(N__91441),
            .I(N__91438));
    LocalMux I__22171 (
            .O(N__91438),
            .I(N__91433));
    InMux I__22170 (
            .O(N__91437),
            .I(N__91428));
    InMux I__22169 (
            .O(N__91436),
            .I(N__91425));
    Span4Mux_v I__22168 (
            .O(N__91433),
            .I(N__91422));
    InMux I__22167 (
            .O(N__91432),
            .I(N__91417));
    InMux I__22166 (
            .O(N__91431),
            .I(N__91417));
    LocalMux I__22165 (
            .O(N__91428),
            .I(N__91412));
    LocalMux I__22164 (
            .O(N__91425),
            .I(N__91412));
    Sp12to4 I__22163 (
            .O(N__91422),
            .I(N__91407));
    LocalMux I__22162 (
            .O(N__91417),
            .I(N__91407));
    Span4Mux_h I__22161 (
            .O(N__91412),
            .I(N__91404));
    Span12Mux_h I__22160 (
            .O(N__91407),
            .I(N__91401));
    Odrv4 I__22159 (
            .O(N__91404),
            .I(\pid_side.error_d_regZ0Z_14 ));
    Odrv12 I__22158 (
            .O(N__91401),
            .I(\pid_side.error_d_regZ0Z_14 ));
    InMux I__22157 (
            .O(N__91396),
            .I(N__91393));
    LocalMux I__22156 (
            .O(N__91393),
            .I(N__91390));
    Span4Mux_h I__22155 (
            .O(N__91390),
            .I(N__91387));
    Odrv4 I__22154 (
            .O(N__91387),
            .I(\pid_side.O_1_24 ));
    CascadeMux I__22153 (
            .O(N__91384),
            .I(N__91371));
    InMux I__22152 (
            .O(N__91383),
            .I(N__91363));
    InMux I__22151 (
            .O(N__91382),
            .I(N__91363));
    InMux I__22150 (
            .O(N__91381),
            .I(N__91363));
    InMux I__22149 (
            .O(N__91380),
            .I(N__91358));
    InMux I__22148 (
            .O(N__91379),
            .I(N__91358));
    InMux I__22147 (
            .O(N__91378),
            .I(N__91354));
    InMux I__22146 (
            .O(N__91377),
            .I(N__91347));
    InMux I__22145 (
            .O(N__91376),
            .I(N__91347));
    InMux I__22144 (
            .O(N__91375),
            .I(N__91347));
    InMux I__22143 (
            .O(N__91374),
            .I(N__91344));
    InMux I__22142 (
            .O(N__91371),
            .I(N__91339));
    InMux I__22141 (
            .O(N__91370),
            .I(N__91339));
    LocalMux I__22140 (
            .O(N__91363),
            .I(N__91334));
    LocalMux I__22139 (
            .O(N__91358),
            .I(N__91334));
    CascadeMux I__22138 (
            .O(N__91357),
            .I(N__91331));
    LocalMux I__22137 (
            .O(N__91354),
            .I(N__91325));
    LocalMux I__22136 (
            .O(N__91347),
            .I(N__91320));
    LocalMux I__22135 (
            .O(N__91344),
            .I(N__91320));
    LocalMux I__22134 (
            .O(N__91339),
            .I(N__91317));
    Span4Mux_h I__22133 (
            .O(N__91334),
            .I(N__91314));
    InMux I__22132 (
            .O(N__91331),
            .I(N__91305));
    InMux I__22131 (
            .O(N__91330),
            .I(N__91305));
    InMux I__22130 (
            .O(N__91329),
            .I(N__91305));
    InMux I__22129 (
            .O(N__91328),
            .I(N__91305));
    Span4Mux_h I__22128 (
            .O(N__91325),
            .I(N__91300));
    Span4Mux_h I__22127 (
            .O(N__91320),
            .I(N__91300));
    Span4Mux_v I__22126 (
            .O(N__91317),
            .I(N__91297));
    Span4Mux_v I__22125 (
            .O(N__91314),
            .I(N__91294));
    LocalMux I__22124 (
            .O(N__91305),
            .I(N__91291));
    Span4Mux_v I__22123 (
            .O(N__91300),
            .I(N__91286));
    Span4Mux_h I__22122 (
            .O(N__91297),
            .I(N__91286));
    Span4Mux_h I__22121 (
            .O(N__91294),
            .I(N__91283));
    Span12Mux_h I__22120 (
            .O(N__91291),
            .I(N__91280));
    Span4Mux_h I__22119 (
            .O(N__91286),
            .I(N__91277));
    Odrv4 I__22118 (
            .O(N__91283),
            .I(\pid_side.error_d_regZ0Z_21 ));
    Odrv12 I__22117 (
            .O(N__91280),
            .I(\pid_side.error_d_regZ0Z_21 ));
    Odrv4 I__22116 (
            .O(N__91277),
            .I(\pid_side.error_d_regZ0Z_21 ));
    InMux I__22115 (
            .O(N__91270),
            .I(N__91267));
    LocalMux I__22114 (
            .O(N__91267),
            .I(N__91264));
    Span4Mux_v I__22113 (
            .O(N__91264),
            .I(N__91260));
    InMux I__22112 (
            .O(N__91263),
            .I(N__91257));
    Span4Mux_h I__22111 (
            .O(N__91260),
            .I(N__91252));
    LocalMux I__22110 (
            .O(N__91257),
            .I(N__91252));
    Odrv4 I__22109 (
            .O(N__91252),
            .I(\pid_side.O_1_15 ));
    InMux I__22108 (
            .O(N__91249),
            .I(N__91240));
    InMux I__22107 (
            .O(N__91248),
            .I(N__91233));
    InMux I__22106 (
            .O(N__91247),
            .I(N__91233));
    InMux I__22105 (
            .O(N__91246),
            .I(N__91226));
    InMux I__22104 (
            .O(N__91245),
            .I(N__91226));
    InMux I__22103 (
            .O(N__91244),
            .I(N__91226));
    InMux I__22102 (
            .O(N__91243),
            .I(N__91223));
    LocalMux I__22101 (
            .O(N__91240),
            .I(N__91220));
    InMux I__22100 (
            .O(N__91239),
            .I(N__91215));
    InMux I__22099 (
            .O(N__91238),
            .I(N__91215));
    LocalMux I__22098 (
            .O(N__91233),
            .I(N__91210));
    LocalMux I__22097 (
            .O(N__91226),
            .I(N__91210));
    LocalMux I__22096 (
            .O(N__91223),
            .I(N__91207));
    Span4Mux_h I__22095 (
            .O(N__91220),
            .I(N__91204));
    LocalMux I__22094 (
            .O(N__91215),
            .I(N__91199));
    Span4Mux_h I__22093 (
            .O(N__91210),
            .I(N__91199));
    Span12Mux_v I__22092 (
            .O(N__91207),
            .I(N__91196));
    Span4Mux_h I__22091 (
            .O(N__91204),
            .I(N__91193));
    Span4Mux_h I__22090 (
            .O(N__91199),
            .I(N__91190));
    Odrv12 I__22089 (
            .O(N__91196),
            .I(\pid_side.error_d_regZ0Z_12 ));
    Odrv4 I__22088 (
            .O(N__91193),
            .I(\pid_side.error_d_regZ0Z_12 ));
    Odrv4 I__22087 (
            .O(N__91190),
            .I(\pid_side.error_d_regZ0Z_12 ));
    InMux I__22086 (
            .O(N__91183),
            .I(N__91180));
    LocalMux I__22085 (
            .O(N__91180),
            .I(N__91177));
    Odrv4 I__22084 (
            .O(N__91177),
            .I(\pid_side.O_1_20 ));
    InMux I__22083 (
            .O(N__91174),
            .I(N__91171));
    LocalMux I__22082 (
            .O(N__91171),
            .I(N__91166));
    InMux I__22081 (
            .O(N__91170),
            .I(N__91161));
    InMux I__22080 (
            .O(N__91169),
            .I(N__91161));
    Span4Mux_v I__22079 (
            .O(N__91166),
            .I(N__91158));
    LocalMux I__22078 (
            .O(N__91161),
            .I(N__91155));
    Span4Mux_h I__22077 (
            .O(N__91158),
            .I(N__91152));
    Span12Mux_v I__22076 (
            .O(N__91155),
            .I(N__91149));
    Span4Mux_h I__22075 (
            .O(N__91152),
            .I(N__91146));
    Odrv12 I__22074 (
            .O(N__91149),
            .I(\pid_side.error_d_regZ0Z_17 ));
    Odrv4 I__22073 (
            .O(N__91146),
            .I(\pid_side.error_d_regZ0Z_17 ));
    InMux I__22072 (
            .O(N__91141),
            .I(N__91138));
    LocalMux I__22071 (
            .O(N__91138),
            .I(N__91135));
    Span4Mux_h I__22070 (
            .O(N__91135),
            .I(N__91132));
    Odrv4 I__22069 (
            .O(N__91132),
            .I(\pid_side.O_1_22 ));
    InMux I__22068 (
            .O(N__91129),
            .I(N__91122));
    InMux I__22067 (
            .O(N__91128),
            .I(N__91122));
    InMux I__22066 (
            .O(N__91127),
            .I(N__91119));
    LocalMux I__22065 (
            .O(N__91122),
            .I(N__91116));
    LocalMux I__22064 (
            .O(N__91119),
            .I(N__91113));
    Span4Mux_h I__22063 (
            .O(N__91116),
            .I(N__91110));
    Span4Mux_h I__22062 (
            .O(N__91113),
            .I(N__91107));
    Span4Mux_v I__22061 (
            .O(N__91110),
            .I(N__91104));
    Odrv4 I__22060 (
            .O(N__91107),
            .I(\pid_side.error_d_regZ0Z_19 ));
    Odrv4 I__22059 (
            .O(N__91104),
            .I(\pid_side.error_d_regZ0Z_19 ));
    InMux I__22058 (
            .O(N__91099),
            .I(N__91096));
    LocalMux I__22057 (
            .O(N__91096),
            .I(N__91093));
    Span4Mux_v I__22056 (
            .O(N__91093),
            .I(N__91090));
    Odrv4 I__22055 (
            .O(N__91090),
            .I(\pid_side.O_1_23 ));
    InMux I__22054 (
            .O(N__91087),
            .I(N__91078));
    InMux I__22053 (
            .O(N__91086),
            .I(N__91078));
    InMux I__22052 (
            .O(N__91085),
            .I(N__91078));
    LocalMux I__22051 (
            .O(N__91078),
            .I(N__91075));
    Span4Mux_h I__22050 (
            .O(N__91075),
            .I(N__91072));
    Span4Mux_v I__22049 (
            .O(N__91072),
            .I(N__91069));
    Span4Mux_h I__22048 (
            .O(N__91069),
            .I(N__91066));
    Span4Mux_v I__22047 (
            .O(N__91066),
            .I(N__91063));
    Odrv4 I__22046 (
            .O(N__91063),
            .I(\pid_side.error_d_regZ0Z_20 ));
    InMux I__22045 (
            .O(N__91060),
            .I(N__91057));
    LocalMux I__22044 (
            .O(N__91057),
            .I(N__91054));
    Odrv4 I__22043 (
            .O(N__91054),
            .I(\pid_side.O_2_23 ));
    InMux I__22042 (
            .O(N__91051),
            .I(N__91045));
    InMux I__22041 (
            .O(N__91050),
            .I(N__91045));
    LocalMux I__22040 (
            .O(N__91045),
            .I(N__91042));
    Span4Mux_v I__22039 (
            .O(N__91042),
            .I(N__91039));
    Span4Mux_h I__22038 (
            .O(N__91039),
            .I(N__91036));
    Odrv4 I__22037 (
            .O(N__91036),
            .I(\pid_side.error_p_regZ0Z_19 ));
    InMux I__22036 (
            .O(N__91033),
            .I(N__91030));
    LocalMux I__22035 (
            .O(N__91030),
            .I(\pid_side.O_2_15 ));
    CascadeMux I__22034 (
            .O(N__91027),
            .I(N__91022));
    InMux I__22033 (
            .O(N__91026),
            .I(N__91017));
    InMux I__22032 (
            .O(N__91025),
            .I(N__91014));
    InMux I__22031 (
            .O(N__91022),
            .I(N__91007));
    InMux I__22030 (
            .O(N__91021),
            .I(N__91007));
    InMux I__22029 (
            .O(N__91020),
            .I(N__91007));
    LocalMux I__22028 (
            .O(N__91017),
            .I(N__91004));
    LocalMux I__22027 (
            .O(N__91014),
            .I(N__90997));
    LocalMux I__22026 (
            .O(N__91007),
            .I(N__90997));
    Span4Mux_h I__22025 (
            .O(N__91004),
            .I(N__90997));
    Span4Mux_h I__22024 (
            .O(N__90997),
            .I(N__90994));
    Odrv4 I__22023 (
            .O(N__90994),
            .I(\pid_side.error_p_regZ0Z_11 ));
    InMux I__22022 (
            .O(N__90991),
            .I(N__90988));
    LocalMux I__22021 (
            .O(N__90988),
            .I(N__90985));
    Odrv4 I__22020 (
            .O(N__90985),
            .I(\pid_side.O_2_16 ));
    InMux I__22019 (
            .O(N__90982),
            .I(N__90979));
    LocalMux I__22018 (
            .O(N__90979),
            .I(N__90975));
    CascadeMux I__22017 (
            .O(N__90978),
            .I(N__90969));
    Span4Mux_h I__22016 (
            .O(N__90975),
            .I(N__90964));
    InMux I__22015 (
            .O(N__90974),
            .I(N__90961));
    InMux I__22014 (
            .O(N__90973),
            .I(N__90958));
    InMux I__22013 (
            .O(N__90972),
            .I(N__90955));
    InMux I__22012 (
            .O(N__90969),
            .I(N__90948));
    InMux I__22011 (
            .O(N__90968),
            .I(N__90948));
    InMux I__22010 (
            .O(N__90967),
            .I(N__90948));
    Span4Mux_h I__22009 (
            .O(N__90964),
            .I(N__90945));
    LocalMux I__22008 (
            .O(N__90961),
            .I(N__90936));
    LocalMux I__22007 (
            .O(N__90958),
            .I(N__90936));
    LocalMux I__22006 (
            .O(N__90955),
            .I(N__90936));
    LocalMux I__22005 (
            .O(N__90948),
            .I(N__90936));
    Odrv4 I__22004 (
            .O(N__90945),
            .I(\pid_side.error_p_regZ0Z_12 ));
    Odrv12 I__22003 (
            .O(N__90936),
            .I(\pid_side.error_p_regZ0Z_12 ));
    InMux I__22002 (
            .O(N__90931),
            .I(N__90928));
    LocalMux I__22001 (
            .O(N__90928),
            .I(N__90925));
    Odrv4 I__22000 (
            .O(N__90925),
            .I(\pid_side.O_2_17 ));
    CascadeMux I__21999 (
            .O(N__90922),
            .I(N__90919));
    InMux I__21998 (
            .O(N__90919),
            .I(N__90912));
    InMux I__21997 (
            .O(N__90918),
            .I(N__90912));
    CascadeMux I__21996 (
            .O(N__90917),
            .I(N__90908));
    LocalMux I__21995 (
            .O(N__90912),
            .I(N__90904));
    InMux I__21994 (
            .O(N__90911),
            .I(N__90901));
    InMux I__21993 (
            .O(N__90908),
            .I(N__90893));
    InMux I__21992 (
            .O(N__90907),
            .I(N__90893));
    Span4Mux_h I__21991 (
            .O(N__90904),
            .I(N__90890));
    LocalMux I__21990 (
            .O(N__90901),
            .I(N__90887));
    InMux I__21989 (
            .O(N__90900),
            .I(N__90880));
    InMux I__21988 (
            .O(N__90899),
            .I(N__90880));
    InMux I__21987 (
            .O(N__90898),
            .I(N__90880));
    LocalMux I__21986 (
            .O(N__90893),
            .I(N__90877));
    Sp12to4 I__21985 (
            .O(N__90890),
            .I(N__90870));
    Span12Mux_h I__21984 (
            .O(N__90887),
            .I(N__90870));
    LocalMux I__21983 (
            .O(N__90880),
            .I(N__90870));
    Odrv4 I__21982 (
            .O(N__90877),
            .I(\pid_side.error_p_regZ0Z_13 ));
    Odrv12 I__21981 (
            .O(N__90870),
            .I(\pid_side.error_p_regZ0Z_13 ));
    InMux I__21980 (
            .O(N__90865),
            .I(N__90862));
    LocalMux I__21979 (
            .O(N__90862),
            .I(N__90859));
    Odrv4 I__21978 (
            .O(N__90859),
            .I(\pid_side.O_2_18 ));
    InMux I__21977 (
            .O(N__90856),
            .I(N__90852));
    CascadeMux I__21976 (
            .O(N__90855),
            .I(N__90848));
    LocalMux I__21975 (
            .O(N__90852),
            .I(N__90844));
    InMux I__21974 (
            .O(N__90851),
            .I(N__90841));
    InMux I__21973 (
            .O(N__90848),
            .I(N__90836));
    InMux I__21972 (
            .O(N__90847),
            .I(N__90836));
    Span4Mux_h I__21971 (
            .O(N__90844),
            .I(N__90833));
    LocalMux I__21970 (
            .O(N__90841),
            .I(N__90828));
    LocalMux I__21969 (
            .O(N__90836),
            .I(N__90828));
    Odrv4 I__21968 (
            .O(N__90833),
            .I(\pid_side.error_p_regZ0Z_14 ));
    Odrv12 I__21967 (
            .O(N__90828),
            .I(\pid_side.error_p_regZ0Z_14 ));
    InMux I__21966 (
            .O(N__90823),
            .I(N__90820));
    LocalMux I__21965 (
            .O(N__90820),
            .I(N__90817));
    Odrv4 I__21964 (
            .O(N__90817),
            .I(\pid_side.O_2_19 ));
    InMux I__21963 (
            .O(N__90814),
            .I(N__90808));
    InMux I__21962 (
            .O(N__90813),
            .I(N__90808));
    LocalMux I__21961 (
            .O(N__90808),
            .I(N__90805));
    Span4Mux_h I__21960 (
            .O(N__90805),
            .I(N__90802));
    Span4Mux_v I__21959 (
            .O(N__90802),
            .I(N__90799));
    Odrv4 I__21958 (
            .O(N__90799),
            .I(\pid_side.error_p_regZ0Z_15 ));
    InMux I__21957 (
            .O(N__90796),
            .I(N__90793));
    LocalMux I__21956 (
            .O(N__90793),
            .I(\pid_side.O_2_21 ));
    InMux I__21955 (
            .O(N__90790),
            .I(N__90786));
    InMux I__21954 (
            .O(N__90789),
            .I(N__90783));
    LocalMux I__21953 (
            .O(N__90786),
            .I(N__90780));
    LocalMux I__21952 (
            .O(N__90783),
            .I(N__90777));
    Span4Mux_v I__21951 (
            .O(N__90780),
            .I(N__90774));
    Span4Mux_h I__21950 (
            .O(N__90777),
            .I(N__90771));
    Span4Mux_h I__21949 (
            .O(N__90774),
            .I(N__90768));
    Span4Mux_h I__21948 (
            .O(N__90771),
            .I(N__90765));
    Span4Mux_h I__21947 (
            .O(N__90768),
            .I(N__90762));
    Span4Mux_h I__21946 (
            .O(N__90765),
            .I(N__90759));
    Odrv4 I__21945 (
            .O(N__90762),
            .I(\pid_side.error_p_regZ0Z_17 ));
    Odrv4 I__21944 (
            .O(N__90759),
            .I(\pid_side.error_p_regZ0Z_17 ));
    InMux I__21943 (
            .O(N__90754),
            .I(N__90751));
    LocalMux I__21942 (
            .O(N__90751),
            .I(\pid_side.O_2_22 ));
    InMux I__21941 (
            .O(N__90748),
            .I(N__90745));
    LocalMux I__21940 (
            .O(N__90745),
            .I(N__90741));
    InMux I__21939 (
            .O(N__90744),
            .I(N__90738));
    Span4Mux_h I__21938 (
            .O(N__90741),
            .I(N__90735));
    LocalMux I__21937 (
            .O(N__90738),
            .I(N__90732));
    Odrv4 I__21936 (
            .O(N__90735),
            .I(\pid_side.error_p_regZ0Z_18 ));
    Odrv4 I__21935 (
            .O(N__90732),
            .I(\pid_side.error_p_regZ0Z_18 ));
    InMux I__21934 (
            .O(N__90727),
            .I(N__90724));
    LocalMux I__21933 (
            .O(N__90724),
            .I(N__90721));
    Span4Mux_v I__21932 (
            .O(N__90721),
            .I(N__90718));
    Odrv4 I__21931 (
            .O(N__90718),
            .I(\pid_side.O_2_5 ));
    InMux I__21930 (
            .O(N__90715),
            .I(N__90710));
    CascadeMux I__21929 (
            .O(N__90714),
            .I(N__90707));
    CascadeMux I__21928 (
            .O(N__90713),
            .I(N__90704));
    LocalMux I__21927 (
            .O(N__90710),
            .I(N__90701));
    InMux I__21926 (
            .O(N__90707),
            .I(N__90696));
    InMux I__21925 (
            .O(N__90704),
            .I(N__90696));
    Span12Mux_h I__21924 (
            .O(N__90701),
            .I(N__90693));
    LocalMux I__21923 (
            .O(N__90696),
            .I(N__90690));
    Odrv12 I__21922 (
            .O(N__90693),
            .I(\pid_side.error_p_regZ0Z_1 ));
    Odrv12 I__21921 (
            .O(N__90690),
            .I(\pid_side.error_p_regZ0Z_1 ));
    CascadeMux I__21920 (
            .O(N__90685),
            .I(N__90682));
    InMux I__21919 (
            .O(N__90682),
            .I(N__90678));
    CascadeMux I__21918 (
            .O(N__90681),
            .I(N__90672));
    LocalMux I__21917 (
            .O(N__90678),
            .I(N__90664));
    CascadeMux I__21916 (
            .O(N__90677),
            .I(N__90659));
    CascadeMux I__21915 (
            .O(N__90676),
            .I(N__90654));
    InMux I__21914 (
            .O(N__90675),
            .I(N__90650));
    InMux I__21913 (
            .O(N__90672),
            .I(N__90642));
    InMux I__21912 (
            .O(N__90671),
            .I(N__90639));
    InMux I__21911 (
            .O(N__90670),
            .I(N__90636));
    InMux I__21910 (
            .O(N__90669),
            .I(N__90629));
    InMux I__21909 (
            .O(N__90668),
            .I(N__90629));
    InMux I__21908 (
            .O(N__90667),
            .I(N__90629));
    Span4Mux_v I__21907 (
            .O(N__90664),
            .I(N__90626));
    InMux I__21906 (
            .O(N__90663),
            .I(N__90623));
    InMux I__21905 (
            .O(N__90662),
            .I(N__90620));
    InMux I__21904 (
            .O(N__90659),
            .I(N__90617));
    CascadeMux I__21903 (
            .O(N__90658),
            .I(N__90614));
    CascadeMux I__21902 (
            .O(N__90657),
            .I(N__90610));
    InMux I__21901 (
            .O(N__90654),
            .I(N__90607));
    CascadeMux I__21900 (
            .O(N__90653),
            .I(N__90604));
    LocalMux I__21899 (
            .O(N__90650),
            .I(N__90601));
    CascadeMux I__21898 (
            .O(N__90649),
            .I(N__90597));
    InMux I__21897 (
            .O(N__90648),
            .I(N__90594));
    CascadeMux I__21896 (
            .O(N__90647),
            .I(N__90591));
    InMux I__21895 (
            .O(N__90646),
            .I(N__90588));
    CascadeMux I__21894 (
            .O(N__90645),
            .I(N__90585));
    LocalMux I__21893 (
            .O(N__90642),
            .I(N__90582));
    LocalMux I__21892 (
            .O(N__90639),
            .I(N__90579));
    LocalMux I__21891 (
            .O(N__90636),
            .I(N__90574));
    LocalMux I__21890 (
            .O(N__90629),
            .I(N__90574));
    Span4Mux_v I__21889 (
            .O(N__90626),
            .I(N__90567));
    LocalMux I__21888 (
            .O(N__90623),
            .I(N__90567));
    LocalMux I__21887 (
            .O(N__90620),
            .I(N__90567));
    LocalMux I__21886 (
            .O(N__90617),
            .I(N__90564));
    InMux I__21885 (
            .O(N__90614),
            .I(N__90561));
    CascadeMux I__21884 (
            .O(N__90613),
            .I(N__90558));
    InMux I__21883 (
            .O(N__90610),
            .I(N__90555));
    LocalMux I__21882 (
            .O(N__90607),
            .I(N__90552));
    InMux I__21881 (
            .O(N__90604),
            .I(N__90549));
    Span4Mux_v I__21880 (
            .O(N__90601),
            .I(N__90546));
    InMux I__21879 (
            .O(N__90600),
            .I(N__90539));
    InMux I__21878 (
            .O(N__90597),
            .I(N__90539));
    LocalMux I__21877 (
            .O(N__90594),
            .I(N__90536));
    InMux I__21876 (
            .O(N__90591),
            .I(N__90533));
    LocalMux I__21875 (
            .O(N__90588),
            .I(N__90530));
    InMux I__21874 (
            .O(N__90585),
            .I(N__90527));
    Span4Mux_v I__21873 (
            .O(N__90582),
            .I(N__90518));
    Span4Mux_v I__21872 (
            .O(N__90579),
            .I(N__90518));
    Span4Mux_v I__21871 (
            .O(N__90574),
            .I(N__90518));
    Span4Mux_h I__21870 (
            .O(N__90567),
            .I(N__90518));
    Span4Mux_v I__21869 (
            .O(N__90564),
            .I(N__90515));
    LocalMux I__21868 (
            .O(N__90561),
            .I(N__90512));
    InMux I__21867 (
            .O(N__90558),
            .I(N__90509));
    LocalMux I__21866 (
            .O(N__90555),
            .I(N__90506));
    Span4Mux_v I__21865 (
            .O(N__90552),
            .I(N__90499));
    LocalMux I__21864 (
            .O(N__90549),
            .I(N__90499));
    Span4Mux_h I__21863 (
            .O(N__90546),
            .I(N__90499));
    CascadeMux I__21862 (
            .O(N__90545),
            .I(N__90495));
    InMux I__21861 (
            .O(N__90544),
            .I(N__90492));
    LocalMux I__21860 (
            .O(N__90539),
            .I(N__90489));
    Span4Mux_v I__21859 (
            .O(N__90536),
            .I(N__90486));
    LocalMux I__21858 (
            .O(N__90533),
            .I(N__90477));
    Span4Mux_v I__21857 (
            .O(N__90530),
            .I(N__90477));
    LocalMux I__21856 (
            .O(N__90527),
            .I(N__90477));
    Span4Mux_h I__21855 (
            .O(N__90518),
            .I(N__90477));
    Span4Mux_h I__21854 (
            .O(N__90515),
            .I(N__90468));
    Span4Mux_v I__21853 (
            .O(N__90512),
            .I(N__90468));
    LocalMux I__21852 (
            .O(N__90509),
            .I(N__90468));
    Span4Mux_h I__21851 (
            .O(N__90506),
            .I(N__90468));
    Span4Mux_v I__21850 (
            .O(N__90499),
            .I(N__90465));
    InMux I__21849 (
            .O(N__90498),
            .I(N__90460));
    InMux I__21848 (
            .O(N__90495),
            .I(N__90460));
    LocalMux I__21847 (
            .O(N__90492),
            .I(N__90451));
    Span4Mux_v I__21846 (
            .O(N__90489),
            .I(N__90451));
    Span4Mux_h I__21845 (
            .O(N__90486),
            .I(N__90451));
    Span4Mux_h I__21844 (
            .O(N__90477),
            .I(N__90451));
    Odrv4 I__21843 (
            .O(N__90468),
            .I(xy_ki_1_rep1));
    Odrv4 I__21842 (
            .O(N__90465),
            .I(xy_ki_1_rep1));
    LocalMux I__21841 (
            .O(N__90460),
            .I(xy_ki_1_rep1));
    Odrv4 I__21840 (
            .O(N__90451),
            .I(xy_ki_1_rep1));
    CascadeMux I__21839 (
            .O(N__90442),
            .I(N__90438));
    CascadeMux I__21838 (
            .O(N__90441),
            .I(N__90428));
    InMux I__21837 (
            .O(N__90438),
            .I(N__90420));
    InMux I__21836 (
            .O(N__90437),
            .I(N__90420));
    InMux I__21835 (
            .O(N__90436),
            .I(N__90420));
    CascadeMux I__21834 (
            .O(N__90435),
            .I(N__90416));
    InMux I__21833 (
            .O(N__90434),
            .I(N__90413));
    InMux I__21832 (
            .O(N__90433),
            .I(N__90409));
    InMux I__21831 (
            .O(N__90432),
            .I(N__90405));
    InMux I__21830 (
            .O(N__90431),
            .I(N__90401));
    InMux I__21829 (
            .O(N__90428),
            .I(N__90398));
    InMux I__21828 (
            .O(N__90427),
            .I(N__90392));
    LocalMux I__21827 (
            .O(N__90420),
            .I(N__90389));
    InMux I__21826 (
            .O(N__90419),
            .I(N__90386));
    InMux I__21825 (
            .O(N__90416),
            .I(N__90383));
    LocalMux I__21824 (
            .O(N__90413),
            .I(N__90380));
    InMux I__21823 (
            .O(N__90412),
            .I(N__90373));
    LocalMux I__21822 (
            .O(N__90409),
            .I(N__90370));
    CascadeMux I__21821 (
            .O(N__90408),
            .I(N__90367));
    LocalMux I__21820 (
            .O(N__90405),
            .I(N__90364));
    InMux I__21819 (
            .O(N__90404),
            .I(N__90361));
    LocalMux I__21818 (
            .O(N__90401),
            .I(N__90356));
    LocalMux I__21817 (
            .O(N__90398),
            .I(N__90356));
    InMux I__21816 (
            .O(N__90397),
            .I(N__90351));
    InMux I__21815 (
            .O(N__90396),
            .I(N__90351));
    InMux I__21814 (
            .O(N__90395),
            .I(N__90348));
    LocalMux I__21813 (
            .O(N__90392),
            .I(N__90344));
    Span4Mux_h I__21812 (
            .O(N__90389),
            .I(N__90336));
    LocalMux I__21811 (
            .O(N__90386),
            .I(N__90336));
    LocalMux I__21810 (
            .O(N__90383),
            .I(N__90336));
    Span4Mux_h I__21809 (
            .O(N__90380),
            .I(N__90333));
    InMux I__21808 (
            .O(N__90379),
            .I(N__90324));
    InMux I__21807 (
            .O(N__90378),
            .I(N__90324));
    InMux I__21806 (
            .O(N__90377),
            .I(N__90324));
    InMux I__21805 (
            .O(N__90376),
            .I(N__90324));
    LocalMux I__21804 (
            .O(N__90373),
            .I(N__90321));
    Span4Mux_v I__21803 (
            .O(N__90370),
            .I(N__90318));
    InMux I__21802 (
            .O(N__90367),
            .I(N__90315));
    Span4Mux_v I__21801 (
            .O(N__90364),
            .I(N__90310));
    LocalMux I__21800 (
            .O(N__90361),
            .I(N__90310));
    Span4Mux_v I__21799 (
            .O(N__90356),
            .I(N__90303));
    LocalMux I__21798 (
            .O(N__90351),
            .I(N__90303));
    LocalMux I__21797 (
            .O(N__90348),
            .I(N__90303));
    CascadeMux I__21796 (
            .O(N__90347),
            .I(N__90299));
    Span4Mux_h I__21795 (
            .O(N__90344),
            .I(N__90296));
    InMux I__21794 (
            .O(N__90343),
            .I(N__90293));
    Span4Mux_v I__21793 (
            .O(N__90336),
            .I(N__90288));
    Span4Mux_h I__21792 (
            .O(N__90333),
            .I(N__90288));
    LocalMux I__21791 (
            .O(N__90324),
            .I(N__90283));
    Span12Mux_v I__21790 (
            .O(N__90321),
            .I(N__90283));
    Span4Mux_h I__21789 (
            .O(N__90318),
            .I(N__90274));
    LocalMux I__21788 (
            .O(N__90315),
            .I(N__90274));
    Span4Mux_v I__21787 (
            .O(N__90310),
            .I(N__90274));
    Span4Mux_v I__21786 (
            .O(N__90303),
            .I(N__90274));
    InMux I__21785 (
            .O(N__90302),
            .I(N__90269));
    InMux I__21784 (
            .O(N__90299),
            .I(N__90269));
    Odrv4 I__21783 (
            .O(N__90296),
            .I(xy_ki_2_rep1));
    LocalMux I__21782 (
            .O(N__90293),
            .I(xy_ki_2_rep1));
    Odrv4 I__21781 (
            .O(N__90288),
            .I(xy_ki_2_rep1));
    Odrv12 I__21780 (
            .O(N__90283),
            .I(xy_ki_2_rep1));
    Odrv4 I__21779 (
            .O(N__90274),
            .I(xy_ki_2_rep1));
    LocalMux I__21778 (
            .O(N__90269),
            .I(xy_ki_2_rep1));
    CascadeMux I__21777 (
            .O(N__90256),
            .I(N__90248));
    CascadeMux I__21776 (
            .O(N__90255),
            .I(N__90244));
    CascadeMux I__21775 (
            .O(N__90254),
            .I(N__90241));
    CascadeMux I__21774 (
            .O(N__90253),
            .I(N__90236));
    InMux I__21773 (
            .O(N__90252),
            .I(N__90231));
    InMux I__21772 (
            .O(N__90251),
            .I(N__90224));
    InMux I__21771 (
            .O(N__90248),
            .I(N__90224));
    InMux I__21770 (
            .O(N__90247),
            .I(N__90224));
    InMux I__21769 (
            .O(N__90244),
            .I(N__90217));
    InMux I__21768 (
            .O(N__90241),
            .I(N__90212));
    InMux I__21767 (
            .O(N__90240),
            .I(N__90212));
    CascadeMux I__21766 (
            .O(N__90239),
            .I(N__90208));
    InMux I__21765 (
            .O(N__90236),
            .I(N__90204));
    InMux I__21764 (
            .O(N__90235),
            .I(N__90201));
    InMux I__21763 (
            .O(N__90234),
            .I(N__90198));
    LocalMux I__21762 (
            .O(N__90231),
            .I(N__90193));
    LocalMux I__21761 (
            .O(N__90224),
            .I(N__90193));
    InMux I__21760 (
            .O(N__90223),
            .I(N__90190));
    InMux I__21759 (
            .O(N__90222),
            .I(N__90185));
    InMux I__21758 (
            .O(N__90221),
            .I(N__90185));
    CascadeMux I__21757 (
            .O(N__90220),
            .I(N__90182));
    LocalMux I__21756 (
            .O(N__90217),
            .I(N__90178));
    LocalMux I__21755 (
            .O(N__90212),
            .I(N__90175));
    InMux I__21754 (
            .O(N__90211),
            .I(N__90168));
    InMux I__21753 (
            .O(N__90208),
            .I(N__90168));
    InMux I__21752 (
            .O(N__90207),
            .I(N__90168));
    LocalMux I__21751 (
            .O(N__90204),
            .I(N__90163));
    LocalMux I__21750 (
            .O(N__90201),
            .I(N__90163));
    LocalMux I__21749 (
            .O(N__90198),
            .I(N__90160));
    Span4Mux_v I__21748 (
            .O(N__90193),
            .I(N__90157));
    LocalMux I__21747 (
            .O(N__90190),
            .I(N__90151));
    LocalMux I__21746 (
            .O(N__90185),
            .I(N__90151));
    InMux I__21745 (
            .O(N__90182),
            .I(N__90146));
    InMux I__21744 (
            .O(N__90181),
            .I(N__90146));
    Span4Mux_v I__21743 (
            .O(N__90178),
            .I(N__90139));
    Span4Mux_v I__21742 (
            .O(N__90175),
            .I(N__90139));
    LocalMux I__21741 (
            .O(N__90168),
            .I(N__90139));
    Span4Mux_v I__21740 (
            .O(N__90163),
            .I(N__90132));
    Span4Mux_v I__21739 (
            .O(N__90160),
            .I(N__90132));
    Span4Mux_h I__21738 (
            .O(N__90157),
            .I(N__90132));
    InMux I__21737 (
            .O(N__90156),
            .I(N__90127));
    Span4Mux_v I__21736 (
            .O(N__90151),
            .I(N__90123));
    LocalMux I__21735 (
            .O(N__90146),
            .I(N__90120));
    Span4Mux_h I__21734 (
            .O(N__90139),
            .I(N__90117));
    Span4Mux_h I__21733 (
            .O(N__90132),
            .I(N__90114));
    InMux I__21732 (
            .O(N__90131),
            .I(N__90109));
    InMux I__21731 (
            .O(N__90130),
            .I(N__90109));
    LocalMux I__21730 (
            .O(N__90127),
            .I(N__90106));
    InMux I__21729 (
            .O(N__90126),
            .I(N__90103));
    Span4Mux_h I__21728 (
            .O(N__90123),
            .I(N__90094));
    Span4Mux_v I__21727 (
            .O(N__90120),
            .I(N__90094));
    Span4Mux_h I__21726 (
            .O(N__90117),
            .I(N__90094));
    Span4Mux_s3_h I__21725 (
            .O(N__90114),
            .I(N__90094));
    LocalMux I__21724 (
            .O(N__90109),
            .I(N__90089));
    Span12Mux_h I__21723 (
            .O(N__90106),
            .I(N__90089));
    LocalMux I__21722 (
            .O(N__90103),
            .I(xy_ki_3_rep1));
    Odrv4 I__21721 (
            .O(N__90094),
            .I(xy_ki_3_rep1));
    Odrv12 I__21720 (
            .O(N__90089),
            .I(xy_ki_3_rep1));
    InMux I__21719 (
            .O(N__90082),
            .I(N__90079));
    LocalMux I__21718 (
            .O(N__90079),
            .I(N__90075));
    InMux I__21717 (
            .O(N__90078),
            .I(N__90072));
    Span4Mux_h I__21716 (
            .O(N__90075),
            .I(N__90069));
    LocalMux I__21715 (
            .O(N__90072),
            .I(N__90066));
    Span4Mux_h I__21714 (
            .O(N__90069),
            .I(N__90063));
    Span4Mux_v I__21713 (
            .O(N__90066),
            .I(N__90060));
    Odrv4 I__21712 (
            .O(N__90063),
            .I(pid_side_m24_2_03_0_a2_0));
    Odrv4 I__21711 (
            .O(N__90060),
            .I(pid_side_m24_2_03_0_a2_0));
    InMux I__21710 (
            .O(N__90055),
            .I(N__90052));
    LocalMux I__21709 (
            .O(N__90052),
            .I(N__90049));
    Odrv4 I__21708 (
            .O(N__90049),
            .I(\pid_side.O_2_20 ));
    InMux I__21707 (
            .O(N__90046),
            .I(N__90040));
    InMux I__21706 (
            .O(N__90045),
            .I(N__90040));
    LocalMux I__21705 (
            .O(N__90040),
            .I(N__90037));
    Span4Mux_h I__21704 (
            .O(N__90037),
            .I(N__90034));
    Span4Mux_h I__21703 (
            .O(N__90034),
            .I(N__90031));
    Span4Mux_h I__21702 (
            .O(N__90031),
            .I(N__90028));
    Odrv4 I__21701 (
            .O(N__90028),
            .I(\pid_side.error_p_regZ0Z_16 ));
    InMux I__21700 (
            .O(N__90025),
            .I(N__90022));
    LocalMux I__21699 (
            .O(N__90022),
            .I(N__90019));
    Odrv4 I__21698 (
            .O(N__90019),
            .I(\pid_side.O_2_10 ));
    CascadeMux I__21697 (
            .O(N__90016),
            .I(N__90011));
    InMux I__21696 (
            .O(N__90015),
            .I(N__90008));
    CascadeMux I__21695 (
            .O(N__90014),
            .I(N__90005));
    InMux I__21694 (
            .O(N__90011),
            .I(N__90002));
    LocalMux I__21693 (
            .O(N__90008),
            .I(N__89999));
    InMux I__21692 (
            .O(N__90005),
            .I(N__89996));
    LocalMux I__21691 (
            .O(N__90002),
            .I(N__89993));
    Span4Mux_h I__21690 (
            .O(N__89999),
            .I(N__89988));
    LocalMux I__21689 (
            .O(N__89996),
            .I(N__89988));
    Span4Mux_h I__21688 (
            .O(N__89993),
            .I(N__89983));
    Span4Mux_h I__21687 (
            .O(N__89988),
            .I(N__89983));
    Odrv4 I__21686 (
            .O(N__89983),
            .I(\pid_side.error_p_regZ0Z_6 ));
    InMux I__21685 (
            .O(N__89980),
            .I(N__89977));
    LocalMux I__21684 (
            .O(N__89977),
            .I(N__89974));
    Odrv4 I__21683 (
            .O(N__89974),
            .I(\pid_side.O_2_11 ));
    CascadeMux I__21682 (
            .O(N__89971),
            .I(N__89967));
    InMux I__21681 (
            .O(N__89970),
            .I(N__89962));
    InMux I__21680 (
            .O(N__89967),
            .I(N__89962));
    LocalMux I__21679 (
            .O(N__89962),
            .I(N__89959));
    Span4Mux_h I__21678 (
            .O(N__89959),
            .I(N__89956));
    Span4Mux_h I__21677 (
            .O(N__89956),
            .I(N__89953));
    Odrv4 I__21676 (
            .O(N__89953),
            .I(\pid_side.error_p_regZ0Z_7 ));
    InMux I__21675 (
            .O(N__89950),
            .I(N__89947));
    LocalMux I__21674 (
            .O(N__89947),
            .I(N__89944));
    Odrv4 I__21673 (
            .O(N__89944),
            .I(\pid_side.O_2_13 ));
    CascadeMux I__21672 (
            .O(N__89941),
            .I(N__89937));
    InMux I__21671 (
            .O(N__89940),
            .I(N__89934));
    InMux I__21670 (
            .O(N__89937),
            .I(N__89931));
    LocalMux I__21669 (
            .O(N__89934),
            .I(N__89928));
    LocalMux I__21668 (
            .O(N__89931),
            .I(N__89923));
    Span4Mux_v I__21667 (
            .O(N__89928),
            .I(N__89923));
    Span4Mux_h I__21666 (
            .O(N__89923),
            .I(N__89920));
    Odrv4 I__21665 (
            .O(N__89920),
            .I(\pid_side.error_p_regZ0Z_9 ));
    InMux I__21664 (
            .O(N__89917),
            .I(N__89914));
    LocalMux I__21663 (
            .O(N__89914),
            .I(N__89911));
    Odrv4 I__21662 (
            .O(N__89911),
            .I(\pid_side.O_2_9 ));
    CascadeMux I__21661 (
            .O(N__89908),
            .I(N__89905));
    InMux I__21660 (
            .O(N__89905),
            .I(N__89902));
    LocalMux I__21659 (
            .O(N__89902),
            .I(N__89898));
    InMux I__21658 (
            .O(N__89901),
            .I(N__89895));
    Span4Mux_v I__21657 (
            .O(N__89898),
            .I(N__89890));
    LocalMux I__21656 (
            .O(N__89895),
            .I(N__89890));
    Span4Mux_h I__21655 (
            .O(N__89890),
            .I(N__89887));
    Odrv4 I__21654 (
            .O(N__89887),
            .I(\pid_side.error_p_regZ0Z_5 ));
    InMux I__21653 (
            .O(N__89884),
            .I(N__89881));
    LocalMux I__21652 (
            .O(N__89881),
            .I(\pid_side.O_2_4 ));
    CascadeMux I__21651 (
            .O(N__89878),
            .I(N__89875));
    InMux I__21650 (
            .O(N__89875),
            .I(N__89871));
    InMux I__21649 (
            .O(N__89874),
            .I(N__89868));
    LocalMux I__21648 (
            .O(N__89871),
            .I(N__89863));
    LocalMux I__21647 (
            .O(N__89868),
            .I(N__89863));
    Span4Mux_h I__21646 (
            .O(N__89863),
            .I(N__89860));
    Span4Mux_v I__21645 (
            .O(N__89860),
            .I(N__89857));
    Span4Mux_h I__21644 (
            .O(N__89857),
            .I(N__89854));
    Odrv4 I__21643 (
            .O(N__89854),
            .I(\pid_side.error_p_regZ0Z_0 ));
    InMux I__21642 (
            .O(N__89851),
            .I(N__89846));
    CascadeMux I__21641 (
            .O(N__89850),
            .I(N__89843));
    CascadeMux I__21640 (
            .O(N__89849),
            .I(N__89839));
    LocalMux I__21639 (
            .O(N__89846),
            .I(N__89834));
    InMux I__21638 (
            .O(N__89843),
            .I(N__89829));
    InMux I__21637 (
            .O(N__89842),
            .I(N__89829));
    InMux I__21636 (
            .O(N__89839),
            .I(N__89823));
    InMux I__21635 (
            .O(N__89838),
            .I(N__89823));
    InMux I__21634 (
            .O(N__89837),
            .I(N__89812));
    Span4Mux_v I__21633 (
            .O(N__89834),
            .I(N__89807));
    LocalMux I__21632 (
            .O(N__89829),
            .I(N__89807));
    InMux I__21631 (
            .O(N__89828),
            .I(N__89804));
    LocalMux I__21630 (
            .O(N__89823),
            .I(N__89801));
    CascadeMux I__21629 (
            .O(N__89822),
            .I(N__89798));
    CascadeMux I__21628 (
            .O(N__89821),
            .I(N__89795));
    InMux I__21627 (
            .O(N__89820),
            .I(N__89790));
    InMux I__21626 (
            .O(N__89819),
            .I(N__89784));
    InMux I__21625 (
            .O(N__89818),
            .I(N__89781));
    InMux I__21624 (
            .O(N__89817),
            .I(N__89778));
    InMux I__21623 (
            .O(N__89816),
            .I(N__89775));
    CascadeMux I__21622 (
            .O(N__89815),
            .I(N__89772));
    LocalMux I__21621 (
            .O(N__89812),
            .I(N__89767));
    Span4Mux_h I__21620 (
            .O(N__89807),
            .I(N__89767));
    LocalMux I__21619 (
            .O(N__89804),
            .I(N__89762));
    Span4Mux_v I__21618 (
            .O(N__89801),
            .I(N__89762));
    InMux I__21617 (
            .O(N__89798),
            .I(N__89759));
    InMux I__21616 (
            .O(N__89795),
            .I(N__89756));
    InMux I__21615 (
            .O(N__89794),
            .I(N__89752));
    InMux I__21614 (
            .O(N__89793),
            .I(N__89749));
    LocalMux I__21613 (
            .O(N__89790),
            .I(N__89743));
    InMux I__21612 (
            .O(N__89789),
            .I(N__89740));
    InMux I__21611 (
            .O(N__89788),
            .I(N__89737));
    InMux I__21610 (
            .O(N__89787),
            .I(N__89734));
    LocalMux I__21609 (
            .O(N__89784),
            .I(N__89731));
    LocalMux I__21608 (
            .O(N__89781),
            .I(N__89727));
    LocalMux I__21607 (
            .O(N__89778),
            .I(N__89724));
    LocalMux I__21606 (
            .O(N__89775),
            .I(N__89721));
    InMux I__21605 (
            .O(N__89772),
            .I(N__89718));
    Span4Mux_v I__21604 (
            .O(N__89767),
            .I(N__89711));
    Span4Mux_h I__21603 (
            .O(N__89762),
            .I(N__89711));
    LocalMux I__21602 (
            .O(N__89759),
            .I(N__89711));
    LocalMux I__21601 (
            .O(N__89756),
            .I(N__89708));
    InMux I__21600 (
            .O(N__89755),
            .I(N__89705));
    LocalMux I__21599 (
            .O(N__89752),
            .I(N__89700));
    LocalMux I__21598 (
            .O(N__89749),
            .I(N__89700));
    InMux I__21597 (
            .O(N__89748),
            .I(N__89697));
    CascadeMux I__21596 (
            .O(N__89747),
            .I(N__89693));
    CascadeMux I__21595 (
            .O(N__89746),
            .I(N__89689));
    Span4Mux_v I__21594 (
            .O(N__89743),
            .I(N__89686));
    LocalMux I__21593 (
            .O(N__89740),
            .I(N__89683));
    LocalMux I__21592 (
            .O(N__89737),
            .I(N__89678));
    LocalMux I__21591 (
            .O(N__89734),
            .I(N__89678));
    Span4Mux_v I__21590 (
            .O(N__89731),
            .I(N__89675));
    InMux I__21589 (
            .O(N__89730),
            .I(N__89672));
    Span4Mux_v I__21588 (
            .O(N__89727),
            .I(N__89665));
    Span4Mux_v I__21587 (
            .O(N__89724),
            .I(N__89665));
    Span4Mux_v I__21586 (
            .O(N__89721),
            .I(N__89665));
    LocalMux I__21585 (
            .O(N__89718),
            .I(N__89658));
    Span4Mux_v I__21584 (
            .O(N__89711),
            .I(N__89658));
    Span4Mux_v I__21583 (
            .O(N__89708),
            .I(N__89658));
    LocalMux I__21582 (
            .O(N__89705),
            .I(N__89655));
    Span4Mux_h I__21581 (
            .O(N__89700),
            .I(N__89652));
    LocalMux I__21580 (
            .O(N__89697),
            .I(N__89649));
    InMux I__21579 (
            .O(N__89696),
            .I(N__89640));
    InMux I__21578 (
            .O(N__89693),
            .I(N__89640));
    InMux I__21577 (
            .O(N__89692),
            .I(N__89640));
    InMux I__21576 (
            .O(N__89689),
            .I(N__89640));
    Span4Mux_h I__21575 (
            .O(N__89686),
            .I(N__89635));
    Span4Mux_v I__21574 (
            .O(N__89683),
            .I(N__89635));
    Span4Mux_h I__21573 (
            .O(N__89678),
            .I(N__89628));
    Span4Mux_h I__21572 (
            .O(N__89675),
            .I(N__89628));
    LocalMux I__21571 (
            .O(N__89672),
            .I(N__89628));
    Span4Mux_s3_h I__21570 (
            .O(N__89665),
            .I(N__89623));
    Span4Mux_h I__21569 (
            .O(N__89658),
            .I(N__89623));
    Span12Mux_h I__21568 (
            .O(N__89655),
            .I(N__89618));
    Sp12to4 I__21567 (
            .O(N__89652),
            .I(N__89618));
    Odrv12 I__21566 (
            .O(N__89649),
            .I(xy_ki_0));
    LocalMux I__21565 (
            .O(N__89640),
            .I(xy_ki_0));
    Odrv4 I__21564 (
            .O(N__89635),
            .I(xy_ki_0));
    Odrv4 I__21563 (
            .O(N__89628),
            .I(xy_ki_0));
    Odrv4 I__21562 (
            .O(N__89623),
            .I(xy_ki_0));
    Odrv12 I__21561 (
            .O(N__89618),
            .I(xy_ki_0));
    CascadeMux I__21560 (
            .O(N__89605),
            .I(N__89598));
    InMux I__21559 (
            .O(N__89604),
            .I(N__89593));
    InMux I__21558 (
            .O(N__89603),
            .I(N__89593));
    CascadeMux I__21557 (
            .O(N__89602),
            .I(N__89587));
    CascadeMux I__21556 (
            .O(N__89601),
            .I(N__89583));
    InMux I__21555 (
            .O(N__89598),
            .I(N__89580));
    LocalMux I__21554 (
            .O(N__89593),
            .I(N__89577));
    CascadeMux I__21553 (
            .O(N__89592),
            .I(N__89573));
    InMux I__21552 (
            .O(N__89591),
            .I(N__89569));
    InMux I__21551 (
            .O(N__89590),
            .I(N__89564));
    InMux I__21550 (
            .O(N__89587),
            .I(N__89564));
    CascadeMux I__21549 (
            .O(N__89586),
            .I(N__89559));
    InMux I__21548 (
            .O(N__89583),
            .I(N__89556));
    LocalMux I__21547 (
            .O(N__89580),
            .I(N__89553));
    Span4Mux_v I__21546 (
            .O(N__89577),
            .I(N__89550));
    InMux I__21545 (
            .O(N__89576),
            .I(N__89547));
    InMux I__21544 (
            .O(N__89573),
            .I(N__89544));
    InMux I__21543 (
            .O(N__89572),
            .I(N__89541));
    LocalMux I__21542 (
            .O(N__89569),
            .I(N__89536));
    LocalMux I__21541 (
            .O(N__89564),
            .I(N__89536));
    InMux I__21540 (
            .O(N__89563),
            .I(N__89532));
    InMux I__21539 (
            .O(N__89562),
            .I(N__89527));
    InMux I__21538 (
            .O(N__89559),
            .I(N__89522));
    LocalMux I__21537 (
            .O(N__89556),
            .I(N__89518));
    Span4Mux_h I__21536 (
            .O(N__89553),
            .I(N__89509));
    Span4Mux_h I__21535 (
            .O(N__89550),
            .I(N__89509));
    LocalMux I__21534 (
            .O(N__89547),
            .I(N__89509));
    LocalMux I__21533 (
            .O(N__89544),
            .I(N__89509));
    LocalMux I__21532 (
            .O(N__89541),
            .I(N__89503));
    Span4Mux_v I__21531 (
            .O(N__89536),
            .I(N__89503));
    InMux I__21530 (
            .O(N__89535),
            .I(N__89499));
    LocalMux I__21529 (
            .O(N__89532),
            .I(N__89496));
    CascadeMux I__21528 (
            .O(N__89531),
            .I(N__89491));
    CascadeMux I__21527 (
            .O(N__89530),
            .I(N__89488));
    LocalMux I__21526 (
            .O(N__89527),
            .I(N__89485));
    InMux I__21525 (
            .O(N__89526),
            .I(N__89480));
    InMux I__21524 (
            .O(N__89525),
            .I(N__89480));
    LocalMux I__21523 (
            .O(N__89522),
            .I(N__89477));
    CascadeMux I__21522 (
            .O(N__89521),
            .I(N__89474));
    Span4Mux_h I__21521 (
            .O(N__89518),
            .I(N__89469));
    Span4Mux_v I__21520 (
            .O(N__89509),
            .I(N__89469));
    CascadeMux I__21519 (
            .O(N__89508),
            .I(N__89465));
    Span4Mux_h I__21518 (
            .O(N__89503),
            .I(N__89462));
    InMux I__21517 (
            .O(N__89502),
            .I(N__89459));
    LocalMux I__21516 (
            .O(N__89499),
            .I(N__89454));
    Span4Mux_v I__21515 (
            .O(N__89496),
            .I(N__89454));
    InMux I__21514 (
            .O(N__89495),
            .I(N__89451));
    InMux I__21513 (
            .O(N__89494),
            .I(N__89444));
    InMux I__21512 (
            .O(N__89491),
            .I(N__89444));
    InMux I__21511 (
            .O(N__89488),
            .I(N__89444));
    Span4Mux_v I__21510 (
            .O(N__89485),
            .I(N__89439));
    LocalMux I__21509 (
            .O(N__89480),
            .I(N__89439));
    Span4Mux_h I__21508 (
            .O(N__89477),
            .I(N__89433));
    InMux I__21507 (
            .O(N__89474),
            .I(N__89430));
    Span4Mux_h I__21506 (
            .O(N__89469),
            .I(N__89427));
    InMux I__21505 (
            .O(N__89468),
            .I(N__89422));
    InMux I__21504 (
            .O(N__89465),
            .I(N__89422));
    Span4Mux_h I__21503 (
            .O(N__89462),
            .I(N__89411));
    LocalMux I__21502 (
            .O(N__89459),
            .I(N__89411));
    Span4Mux_h I__21501 (
            .O(N__89454),
            .I(N__89411));
    LocalMux I__21500 (
            .O(N__89451),
            .I(N__89411));
    LocalMux I__21499 (
            .O(N__89444),
            .I(N__89411));
    Span4Mux_h I__21498 (
            .O(N__89439),
            .I(N__89408));
    InMux I__21497 (
            .O(N__89438),
            .I(N__89405));
    InMux I__21496 (
            .O(N__89437),
            .I(N__89400));
    InMux I__21495 (
            .O(N__89436),
            .I(N__89400));
    Span4Mux_v I__21494 (
            .O(N__89433),
            .I(N__89391));
    LocalMux I__21493 (
            .O(N__89430),
            .I(N__89391));
    Span4Mux_s3_h I__21492 (
            .O(N__89427),
            .I(N__89391));
    LocalMux I__21491 (
            .O(N__89422),
            .I(N__89391));
    Span4Mux_v I__21490 (
            .O(N__89411),
            .I(N__89386));
    Span4Mux_s3_h I__21489 (
            .O(N__89408),
            .I(N__89386));
    LocalMux I__21488 (
            .O(N__89405),
            .I(xy_ki_2_rep2));
    LocalMux I__21487 (
            .O(N__89400),
            .I(xy_ki_2_rep2));
    Odrv4 I__21486 (
            .O(N__89391),
            .I(xy_ki_2_rep2));
    Odrv4 I__21485 (
            .O(N__89386),
            .I(xy_ki_2_rep2));
    InMux I__21484 (
            .O(N__89377),
            .I(N__89369));
    CascadeMux I__21483 (
            .O(N__89376),
            .I(N__89366));
    CascadeMux I__21482 (
            .O(N__89375),
            .I(N__89363));
    CascadeMux I__21481 (
            .O(N__89374),
            .I(N__89360));
    InMux I__21480 (
            .O(N__89373),
            .I(N__89355));
    InMux I__21479 (
            .O(N__89372),
            .I(N__89355));
    LocalMux I__21478 (
            .O(N__89369),
            .I(N__89348));
    InMux I__21477 (
            .O(N__89366),
            .I(N__89342));
    InMux I__21476 (
            .O(N__89363),
            .I(N__89339));
    InMux I__21475 (
            .O(N__89360),
            .I(N__89335));
    LocalMux I__21474 (
            .O(N__89355),
            .I(N__89331));
    InMux I__21473 (
            .O(N__89354),
            .I(N__89324));
    InMux I__21472 (
            .O(N__89353),
            .I(N__89324));
    InMux I__21471 (
            .O(N__89352),
            .I(N__89324));
    InMux I__21470 (
            .O(N__89351),
            .I(N__89321));
    Span4Mux_h I__21469 (
            .O(N__89348),
            .I(N__89317));
    InMux I__21468 (
            .O(N__89347),
            .I(N__89312));
    InMux I__21467 (
            .O(N__89346),
            .I(N__89312));
    InMux I__21466 (
            .O(N__89345),
            .I(N__89308));
    LocalMux I__21465 (
            .O(N__89342),
            .I(N__89301));
    LocalMux I__21464 (
            .O(N__89339),
            .I(N__89301));
    InMux I__21463 (
            .O(N__89338),
            .I(N__89297));
    LocalMux I__21462 (
            .O(N__89335),
            .I(N__89294));
    CascadeMux I__21461 (
            .O(N__89334),
            .I(N__89288));
    Span4Mux_v I__21460 (
            .O(N__89331),
            .I(N__89281));
    LocalMux I__21459 (
            .O(N__89324),
            .I(N__89281));
    LocalMux I__21458 (
            .O(N__89321),
            .I(N__89278));
    InMux I__21457 (
            .O(N__89320),
            .I(N__89275));
    Span4Mux_v I__21456 (
            .O(N__89317),
            .I(N__89270));
    LocalMux I__21455 (
            .O(N__89312),
            .I(N__89270));
    CascadeMux I__21454 (
            .O(N__89311),
            .I(N__89267));
    LocalMux I__21453 (
            .O(N__89308),
            .I(N__89264));
    InMux I__21452 (
            .O(N__89307),
            .I(N__89259));
    InMux I__21451 (
            .O(N__89306),
            .I(N__89259));
    Span4Mux_v I__21450 (
            .O(N__89301),
            .I(N__89256));
    InMux I__21449 (
            .O(N__89300),
            .I(N__89253));
    LocalMux I__21448 (
            .O(N__89297),
            .I(N__89247));
    Span4Mux_v I__21447 (
            .O(N__89294),
            .I(N__89247));
    InMux I__21446 (
            .O(N__89293),
            .I(N__89242));
    InMux I__21445 (
            .O(N__89292),
            .I(N__89239));
    InMux I__21444 (
            .O(N__89291),
            .I(N__89234));
    InMux I__21443 (
            .O(N__89288),
            .I(N__89234));
    InMux I__21442 (
            .O(N__89287),
            .I(N__89229));
    InMux I__21441 (
            .O(N__89286),
            .I(N__89226));
    Span4Mux_v I__21440 (
            .O(N__89281),
            .I(N__89223));
    Span4Mux_h I__21439 (
            .O(N__89278),
            .I(N__89216));
    LocalMux I__21438 (
            .O(N__89275),
            .I(N__89216));
    Span4Mux_v I__21437 (
            .O(N__89270),
            .I(N__89216));
    InMux I__21436 (
            .O(N__89267),
            .I(N__89213));
    Span4Mux_h I__21435 (
            .O(N__89264),
            .I(N__89204));
    LocalMux I__21434 (
            .O(N__89259),
            .I(N__89204));
    Span4Mux_h I__21433 (
            .O(N__89256),
            .I(N__89204));
    LocalMux I__21432 (
            .O(N__89253),
            .I(N__89204));
    InMux I__21431 (
            .O(N__89252),
            .I(N__89201));
    Span4Mux_h I__21430 (
            .O(N__89247),
            .I(N__89198));
    InMux I__21429 (
            .O(N__89246),
            .I(N__89193));
    InMux I__21428 (
            .O(N__89245),
            .I(N__89193));
    LocalMux I__21427 (
            .O(N__89242),
            .I(N__89188));
    LocalMux I__21426 (
            .O(N__89239),
            .I(N__89188));
    LocalMux I__21425 (
            .O(N__89234),
            .I(N__89185));
    InMux I__21424 (
            .O(N__89233),
            .I(N__89182));
    InMux I__21423 (
            .O(N__89232),
            .I(N__89179));
    LocalMux I__21422 (
            .O(N__89229),
            .I(N__89172));
    LocalMux I__21421 (
            .O(N__89226),
            .I(N__89172));
    Span4Mux_h I__21420 (
            .O(N__89223),
            .I(N__89172));
    Span4Mux_h I__21419 (
            .O(N__89216),
            .I(N__89169));
    LocalMux I__21418 (
            .O(N__89213),
            .I(N__89164));
    Span4Mux_h I__21417 (
            .O(N__89204),
            .I(N__89164));
    LocalMux I__21416 (
            .O(N__89201),
            .I(N__89156));
    Span4Mux_v I__21415 (
            .O(N__89198),
            .I(N__89156));
    LocalMux I__21414 (
            .O(N__89193),
            .I(N__89156));
    Span4Mux_v I__21413 (
            .O(N__89188),
            .I(N__89149));
    Span4Mux_h I__21412 (
            .O(N__89185),
            .I(N__89149));
    LocalMux I__21411 (
            .O(N__89182),
            .I(N__89149));
    LocalMux I__21410 (
            .O(N__89179),
            .I(N__89144));
    Sp12to4 I__21409 (
            .O(N__89172),
            .I(N__89144));
    Span4Mux_s2_h I__21408 (
            .O(N__89169),
            .I(N__89139));
    Span4Mux_h I__21407 (
            .O(N__89164),
            .I(N__89139));
    InMux I__21406 (
            .O(N__89163),
            .I(N__89136));
    Span4Mux_h I__21405 (
            .O(N__89156),
            .I(N__89133));
    Span4Mux_h I__21404 (
            .O(N__89149),
            .I(N__89130));
    Span12Mux_v I__21403 (
            .O(N__89144),
            .I(N__89127));
    Span4Mux_v I__21402 (
            .O(N__89139),
            .I(N__89124));
    LocalMux I__21401 (
            .O(N__89136),
            .I(xy_ki_3));
    Odrv4 I__21400 (
            .O(N__89133),
            .I(xy_ki_3));
    Odrv4 I__21399 (
            .O(N__89130),
            .I(xy_ki_3));
    Odrv12 I__21398 (
            .O(N__89127),
            .I(xy_ki_3));
    Odrv4 I__21397 (
            .O(N__89124),
            .I(xy_ki_3));
    CascadeMux I__21396 (
            .O(N__89113),
            .I(N__89106));
    InMux I__21395 (
            .O(N__89112),
            .I(N__89103));
    InMux I__21394 (
            .O(N__89111),
            .I(N__89100));
    InMux I__21393 (
            .O(N__89110),
            .I(N__89094));
    InMux I__21392 (
            .O(N__89109),
            .I(N__89091));
    InMux I__21391 (
            .O(N__89106),
            .I(N__89088));
    LocalMux I__21390 (
            .O(N__89103),
            .I(N__89083));
    LocalMux I__21389 (
            .O(N__89100),
            .I(N__89083));
    CascadeMux I__21388 (
            .O(N__89099),
            .I(N__89074));
    InMux I__21387 (
            .O(N__89098),
            .I(N__89069));
    InMux I__21386 (
            .O(N__89097),
            .I(N__89062));
    LocalMux I__21385 (
            .O(N__89094),
            .I(N__89059));
    LocalMux I__21384 (
            .O(N__89091),
            .I(N__89054));
    LocalMux I__21383 (
            .O(N__89088),
            .I(N__89054));
    Span4Mux_h I__21382 (
            .O(N__89083),
            .I(N__89051));
    InMux I__21381 (
            .O(N__89082),
            .I(N__89044));
    InMux I__21380 (
            .O(N__89081),
            .I(N__89044));
    InMux I__21379 (
            .O(N__89080),
            .I(N__89044));
    InMux I__21378 (
            .O(N__89079),
            .I(N__89038));
    InMux I__21377 (
            .O(N__89078),
            .I(N__89038));
    InMux I__21376 (
            .O(N__89077),
            .I(N__89034));
    InMux I__21375 (
            .O(N__89074),
            .I(N__89029));
    InMux I__21374 (
            .O(N__89073),
            .I(N__89029));
    CascadeMux I__21373 (
            .O(N__89072),
            .I(N__89024));
    LocalMux I__21372 (
            .O(N__89069),
            .I(N__89021));
    InMux I__21371 (
            .O(N__89068),
            .I(N__89016));
    InMux I__21370 (
            .O(N__89067),
            .I(N__89016));
    InMux I__21369 (
            .O(N__89066),
            .I(N__89011));
    InMux I__21368 (
            .O(N__89065),
            .I(N__89011));
    LocalMux I__21367 (
            .O(N__89062),
            .I(N__89004));
    Span4Mux_h I__21366 (
            .O(N__89059),
            .I(N__89004));
    Span4Mux_v I__21365 (
            .O(N__89054),
            .I(N__89004));
    Span4Mux_h I__21364 (
            .O(N__89051),
            .I(N__88999));
    LocalMux I__21363 (
            .O(N__89044),
            .I(N__88999));
    InMux I__21362 (
            .O(N__89043),
            .I(N__88996));
    LocalMux I__21361 (
            .O(N__89038),
            .I(N__88993));
    InMux I__21360 (
            .O(N__89037),
            .I(N__88990));
    LocalMux I__21359 (
            .O(N__89034),
            .I(N__88985));
    LocalMux I__21358 (
            .O(N__89029),
            .I(N__88985));
    InMux I__21357 (
            .O(N__89028),
            .I(N__88981));
    InMux I__21356 (
            .O(N__89027),
            .I(N__88976));
    InMux I__21355 (
            .O(N__89024),
            .I(N__88976));
    Span4Mux_v I__21354 (
            .O(N__89021),
            .I(N__88973));
    LocalMux I__21353 (
            .O(N__89016),
            .I(N__88966));
    LocalMux I__21352 (
            .O(N__89011),
            .I(N__88966));
    Span4Mux_h I__21351 (
            .O(N__89004),
            .I(N__88961));
    Span4Mux_v I__21350 (
            .O(N__88999),
            .I(N__88961));
    LocalMux I__21349 (
            .O(N__88996),
            .I(N__88958));
    Span4Mux_v I__21348 (
            .O(N__88993),
            .I(N__88951));
    LocalMux I__21347 (
            .O(N__88990),
            .I(N__88951));
    Span4Mux_v I__21346 (
            .O(N__88985),
            .I(N__88951));
    InMux I__21345 (
            .O(N__88984),
            .I(N__88948));
    LocalMux I__21344 (
            .O(N__88981),
            .I(N__88943));
    LocalMux I__21343 (
            .O(N__88976),
            .I(N__88943));
    Span4Mux_h I__21342 (
            .O(N__88973),
            .I(N__88940));
    InMux I__21341 (
            .O(N__88972),
            .I(N__88937));
    InMux I__21340 (
            .O(N__88971),
            .I(N__88934));
    Span4Mux_h I__21339 (
            .O(N__88966),
            .I(N__88931));
    Span4Mux_h I__21338 (
            .O(N__88961),
            .I(N__88928));
    Span4Mux_v I__21337 (
            .O(N__88958),
            .I(N__88923));
    Span4Mux_h I__21336 (
            .O(N__88951),
            .I(N__88923));
    LocalMux I__21335 (
            .O(N__88948),
            .I(N__88920));
    Span4Mux_v I__21334 (
            .O(N__88943),
            .I(N__88917));
    Span4Mux_h I__21333 (
            .O(N__88940),
            .I(N__88912));
    LocalMux I__21332 (
            .O(N__88937),
            .I(N__88912));
    LocalMux I__21331 (
            .O(N__88934),
            .I(N__88905));
    Span4Mux_h I__21330 (
            .O(N__88931),
            .I(N__88905));
    Span4Mux_s0_h I__21329 (
            .O(N__88928),
            .I(N__88905));
    Span4Mux_h I__21328 (
            .O(N__88923),
            .I(N__88902));
    Span4Mux_h I__21327 (
            .O(N__88920),
            .I(N__88895));
    Span4Mux_h I__21326 (
            .O(N__88917),
            .I(N__88895));
    Span4Mux_v I__21325 (
            .O(N__88912),
            .I(N__88895));
    Odrv4 I__21324 (
            .O(N__88905),
            .I(xy_ki_1_rep2));
    Odrv4 I__21323 (
            .O(N__88902),
            .I(xy_ki_1_rep2));
    Odrv4 I__21322 (
            .O(N__88895),
            .I(xy_ki_1_rep2));
    InMux I__21321 (
            .O(N__88888),
            .I(N__88885));
    LocalMux I__21320 (
            .O(N__88885),
            .I(N__88882));
    Span4Mux_v I__21319 (
            .O(N__88882),
            .I(N__88878));
    InMux I__21318 (
            .O(N__88881),
            .I(N__88875));
    Span4Mux_h I__21317 (
            .O(N__88878),
            .I(N__88872));
    LocalMux I__21316 (
            .O(N__88875),
            .I(N__88869));
    Span4Mux_h I__21315 (
            .O(N__88872),
            .I(N__88864));
    Span4Mux_v I__21314 (
            .O(N__88869),
            .I(N__88864));
    Odrv4 I__21313 (
            .O(N__88864),
            .I(pid_front_N_463_1));
    InMux I__21312 (
            .O(N__88861),
            .I(N__88855));
    InMux I__21311 (
            .O(N__88860),
            .I(N__88851));
    InMux I__21310 (
            .O(N__88859),
            .I(N__88848));
    InMux I__21309 (
            .O(N__88858),
            .I(N__88843));
    LocalMux I__21308 (
            .O(N__88855),
            .I(N__88840));
    InMux I__21307 (
            .O(N__88854),
            .I(N__88837));
    LocalMux I__21306 (
            .O(N__88851),
            .I(N__88834));
    LocalMux I__21305 (
            .O(N__88848),
            .I(N__88831));
    InMux I__21304 (
            .O(N__88847),
            .I(N__88825));
    InMux I__21303 (
            .O(N__88846),
            .I(N__88822));
    LocalMux I__21302 (
            .O(N__88843),
            .I(N__88817));
    Span4Mux_h I__21301 (
            .O(N__88840),
            .I(N__88817));
    LocalMux I__21300 (
            .O(N__88837),
            .I(N__88814));
    Span4Mux_v I__21299 (
            .O(N__88834),
            .I(N__88810));
    Span12Mux_s5_h I__21298 (
            .O(N__88831),
            .I(N__88807));
    InMux I__21297 (
            .O(N__88830),
            .I(N__88802));
    InMux I__21296 (
            .O(N__88829),
            .I(N__88802));
    InMux I__21295 (
            .O(N__88828),
            .I(N__88799));
    LocalMux I__21294 (
            .O(N__88825),
            .I(N__88795));
    LocalMux I__21293 (
            .O(N__88822),
            .I(N__88792));
    Span4Mux_v I__21292 (
            .O(N__88817),
            .I(N__88789));
    Span12Mux_s5_h I__21291 (
            .O(N__88814),
            .I(N__88786));
    InMux I__21290 (
            .O(N__88813),
            .I(N__88783));
    Sp12to4 I__21289 (
            .O(N__88810),
            .I(N__88778));
    Span12Mux_v I__21288 (
            .O(N__88807),
            .I(N__88778));
    LocalMux I__21287 (
            .O(N__88802),
            .I(N__88775));
    LocalMux I__21286 (
            .O(N__88799),
            .I(N__88772));
    InMux I__21285 (
            .O(N__88798),
            .I(N__88769));
    Span4Mux_v I__21284 (
            .O(N__88795),
            .I(N__88762));
    Span4Mux_h I__21283 (
            .O(N__88792),
            .I(N__88762));
    Span4Mux_h I__21282 (
            .O(N__88789),
            .I(N__88759));
    Span12Mux_h I__21281 (
            .O(N__88786),
            .I(N__88756));
    LocalMux I__21280 (
            .O(N__88783),
            .I(N__88751));
    Span12Mux_h I__21279 (
            .O(N__88778),
            .I(N__88751));
    Span4Mux_h I__21278 (
            .O(N__88775),
            .I(N__88744));
    Span4Mux_v I__21277 (
            .O(N__88772),
            .I(N__88744));
    LocalMux I__21276 (
            .O(N__88769),
            .I(N__88744));
    InMux I__21275 (
            .O(N__88768),
            .I(N__88739));
    InMux I__21274 (
            .O(N__88767),
            .I(N__88739));
    Odrv4 I__21273 (
            .O(N__88762),
            .I(uart_pc_data_4));
    Odrv4 I__21272 (
            .O(N__88759),
            .I(uart_pc_data_4));
    Odrv12 I__21271 (
            .O(N__88756),
            .I(uart_pc_data_4));
    Odrv12 I__21270 (
            .O(N__88751),
            .I(uart_pc_data_4));
    Odrv4 I__21269 (
            .O(N__88744),
            .I(uart_pc_data_4));
    LocalMux I__21268 (
            .O(N__88739),
            .I(uart_pc_data_4));
    InMux I__21267 (
            .O(N__88726),
            .I(N__88723));
    LocalMux I__21266 (
            .O(N__88723),
            .I(N__88719));
    InMux I__21265 (
            .O(N__88722),
            .I(N__88716));
    Span4Mux_s2_h I__21264 (
            .O(N__88719),
            .I(N__88713));
    LocalMux I__21263 (
            .O(N__88716),
            .I(N__88710));
    Span4Mux_v I__21262 (
            .O(N__88713),
            .I(N__88705));
    Span4Mux_s2_h I__21261 (
            .O(N__88710),
            .I(N__88705));
    Odrv4 I__21260 (
            .O(N__88705),
            .I(xy_kd_4));
    InMux I__21259 (
            .O(N__88702),
            .I(N__88696));
    InMux I__21258 (
            .O(N__88701),
            .I(N__88692));
    InMux I__21257 (
            .O(N__88700),
            .I(N__88689));
    InMux I__21256 (
            .O(N__88699),
            .I(N__88686));
    LocalMux I__21255 (
            .O(N__88696),
            .I(N__88682));
    InMux I__21254 (
            .O(N__88695),
            .I(N__88679));
    LocalMux I__21253 (
            .O(N__88692),
            .I(N__88676));
    LocalMux I__21252 (
            .O(N__88689),
            .I(N__88673));
    LocalMux I__21251 (
            .O(N__88686),
            .I(N__88670));
    InMux I__21250 (
            .O(N__88685),
            .I(N__88667));
    Span4Mux_v I__21249 (
            .O(N__88682),
            .I(N__88658));
    LocalMux I__21248 (
            .O(N__88679),
            .I(N__88658));
    Span4Mux_v I__21247 (
            .O(N__88676),
            .I(N__88655));
    Span4Mux_v I__21246 (
            .O(N__88673),
            .I(N__88650));
    Span4Mux_v I__21245 (
            .O(N__88670),
            .I(N__88650));
    LocalMux I__21244 (
            .O(N__88667),
            .I(N__88647));
    InMux I__21243 (
            .O(N__88666),
            .I(N__88643));
    InMux I__21242 (
            .O(N__88665),
            .I(N__88637));
    InMux I__21241 (
            .O(N__88664),
            .I(N__88633));
    InMux I__21240 (
            .O(N__88663),
            .I(N__88630));
    Span4Mux_h I__21239 (
            .O(N__88658),
            .I(N__88627));
    Span4Mux_h I__21238 (
            .O(N__88655),
            .I(N__88624));
    Span4Mux_h I__21237 (
            .O(N__88650),
            .I(N__88621));
    Span4Mux_v I__21236 (
            .O(N__88647),
            .I(N__88618));
    InMux I__21235 (
            .O(N__88646),
            .I(N__88615));
    LocalMux I__21234 (
            .O(N__88643),
            .I(N__88612));
    InMux I__21233 (
            .O(N__88642),
            .I(N__88607));
    InMux I__21232 (
            .O(N__88641),
            .I(N__88607));
    CascadeMux I__21231 (
            .O(N__88640),
            .I(N__88604));
    LocalMux I__21230 (
            .O(N__88637),
            .I(N__88601));
    InMux I__21229 (
            .O(N__88636),
            .I(N__88598));
    LocalMux I__21228 (
            .O(N__88633),
            .I(N__88595));
    LocalMux I__21227 (
            .O(N__88630),
            .I(N__88588));
    Span4Mux_v I__21226 (
            .O(N__88627),
            .I(N__88588));
    Span4Mux_h I__21225 (
            .O(N__88624),
            .I(N__88588));
    Span4Mux_h I__21224 (
            .O(N__88621),
            .I(N__88585));
    Span4Mux_h I__21223 (
            .O(N__88618),
            .I(N__88580));
    LocalMux I__21222 (
            .O(N__88615),
            .I(N__88580));
    Span4Mux_v I__21221 (
            .O(N__88612),
            .I(N__88575));
    LocalMux I__21220 (
            .O(N__88607),
            .I(N__88575));
    InMux I__21219 (
            .O(N__88604),
            .I(N__88571));
    Span4Mux_h I__21218 (
            .O(N__88601),
            .I(N__88568));
    LocalMux I__21217 (
            .O(N__88598),
            .I(N__88563));
    Span4Mux_v I__21216 (
            .O(N__88595),
            .I(N__88563));
    Span4Mux_h I__21215 (
            .O(N__88588),
            .I(N__88560));
    Span4Mux_h I__21214 (
            .O(N__88585),
            .I(N__88555));
    Span4Mux_v I__21213 (
            .O(N__88580),
            .I(N__88555));
    Span4Mux_h I__21212 (
            .O(N__88575),
            .I(N__88552));
    InMux I__21211 (
            .O(N__88574),
            .I(N__88549));
    LocalMux I__21210 (
            .O(N__88571),
            .I(uart_pc_data_5));
    Odrv4 I__21209 (
            .O(N__88568),
            .I(uart_pc_data_5));
    Odrv4 I__21208 (
            .O(N__88563),
            .I(uart_pc_data_5));
    Odrv4 I__21207 (
            .O(N__88560),
            .I(uart_pc_data_5));
    Odrv4 I__21206 (
            .O(N__88555),
            .I(uart_pc_data_5));
    Odrv4 I__21205 (
            .O(N__88552),
            .I(uart_pc_data_5));
    LocalMux I__21204 (
            .O(N__88549),
            .I(uart_pc_data_5));
    InMux I__21203 (
            .O(N__88534),
            .I(N__88531));
    LocalMux I__21202 (
            .O(N__88531),
            .I(N__88527));
    InMux I__21201 (
            .O(N__88530),
            .I(N__88524));
    Span4Mux_s0_h I__21200 (
            .O(N__88527),
            .I(N__88521));
    LocalMux I__21199 (
            .O(N__88524),
            .I(N__88518));
    Span4Mux_v I__21198 (
            .O(N__88521),
            .I(N__88513));
    Span4Mux_v I__21197 (
            .O(N__88518),
            .I(N__88513));
    Odrv4 I__21196 (
            .O(N__88513),
            .I(xy_kd_5));
    InMux I__21195 (
            .O(N__88510),
            .I(N__88502));
    InMux I__21194 (
            .O(N__88509),
            .I(N__88499));
    InMux I__21193 (
            .O(N__88508),
            .I(N__88496));
    InMux I__21192 (
            .O(N__88507),
            .I(N__88493));
    InMux I__21191 (
            .O(N__88506),
            .I(N__88490));
    InMux I__21190 (
            .O(N__88505),
            .I(N__88486));
    LocalMux I__21189 (
            .O(N__88502),
            .I(N__88483));
    LocalMux I__21188 (
            .O(N__88499),
            .I(N__88477));
    LocalMux I__21187 (
            .O(N__88496),
            .I(N__88474));
    LocalMux I__21186 (
            .O(N__88493),
            .I(N__88471));
    LocalMux I__21185 (
            .O(N__88490),
            .I(N__88467));
    InMux I__21184 (
            .O(N__88489),
            .I(N__88464));
    LocalMux I__21183 (
            .O(N__88486),
            .I(N__88461));
    Span4Mux_v I__21182 (
            .O(N__88483),
            .I(N__88458));
    InMux I__21181 (
            .O(N__88482),
            .I(N__88454));
    InMux I__21180 (
            .O(N__88481),
            .I(N__88451));
    InMux I__21179 (
            .O(N__88480),
            .I(N__88448));
    Span4Mux_h I__21178 (
            .O(N__88477),
            .I(N__88445));
    Span4Mux_v I__21177 (
            .O(N__88474),
            .I(N__88440));
    Span4Mux_v I__21176 (
            .O(N__88471),
            .I(N__88440));
    InMux I__21175 (
            .O(N__88470),
            .I(N__88437));
    Span4Mux_h I__21174 (
            .O(N__88467),
            .I(N__88434));
    LocalMux I__21173 (
            .O(N__88464),
            .I(N__88431));
    Span4Mux_h I__21172 (
            .O(N__88461),
            .I(N__88426));
    Span4Mux_h I__21171 (
            .O(N__88458),
            .I(N__88426));
    CascadeMux I__21170 (
            .O(N__88457),
            .I(N__88422));
    LocalMux I__21169 (
            .O(N__88454),
            .I(N__88419));
    LocalMux I__21168 (
            .O(N__88451),
            .I(N__88416));
    LocalMux I__21167 (
            .O(N__88448),
            .I(N__88413));
    Span4Mux_v I__21166 (
            .O(N__88445),
            .I(N__88410));
    Sp12to4 I__21165 (
            .O(N__88440),
            .I(N__88407));
    LocalMux I__21164 (
            .O(N__88437),
            .I(N__88404));
    Span4Mux_v I__21163 (
            .O(N__88434),
            .I(N__88401));
    Span4Mux_v I__21162 (
            .O(N__88431),
            .I(N__88396));
    Span4Mux_v I__21161 (
            .O(N__88426),
            .I(N__88396));
    InMux I__21160 (
            .O(N__88425),
            .I(N__88393));
    InMux I__21159 (
            .O(N__88422),
            .I(N__88389));
    Span4Mux_h I__21158 (
            .O(N__88419),
            .I(N__88386));
    Span12Mux_s9_v I__21157 (
            .O(N__88416),
            .I(N__88381));
    Span12Mux_s8_h I__21156 (
            .O(N__88413),
            .I(N__88381));
    Span4Mux_h I__21155 (
            .O(N__88410),
            .I(N__88378));
    Span12Mux_s6_h I__21154 (
            .O(N__88407),
            .I(N__88375));
    Span4Mux_v I__21153 (
            .O(N__88404),
            .I(N__88366));
    Span4Mux_v I__21152 (
            .O(N__88401),
            .I(N__88366));
    Span4Mux_h I__21151 (
            .O(N__88396),
            .I(N__88366));
    LocalMux I__21150 (
            .O(N__88393),
            .I(N__88366));
    InMux I__21149 (
            .O(N__88392),
            .I(N__88363));
    LocalMux I__21148 (
            .O(N__88389),
            .I(uart_pc_data_6));
    Odrv4 I__21147 (
            .O(N__88386),
            .I(uart_pc_data_6));
    Odrv12 I__21146 (
            .O(N__88381),
            .I(uart_pc_data_6));
    Odrv4 I__21145 (
            .O(N__88378),
            .I(uart_pc_data_6));
    Odrv12 I__21144 (
            .O(N__88375),
            .I(uart_pc_data_6));
    Odrv4 I__21143 (
            .O(N__88366),
            .I(uart_pc_data_6));
    LocalMux I__21142 (
            .O(N__88363),
            .I(uart_pc_data_6));
    InMux I__21141 (
            .O(N__88348),
            .I(N__88345));
    LocalMux I__21140 (
            .O(N__88345),
            .I(N__88341));
    InMux I__21139 (
            .O(N__88344),
            .I(N__88338));
    Span4Mux_s2_h I__21138 (
            .O(N__88341),
            .I(N__88335));
    LocalMux I__21137 (
            .O(N__88338),
            .I(N__88332));
    Span4Mux_v I__21136 (
            .O(N__88335),
            .I(N__88327));
    Span4Mux_s2_h I__21135 (
            .O(N__88332),
            .I(N__88327));
    Odrv4 I__21134 (
            .O(N__88327),
            .I(xy_kd_6));
    InMux I__21133 (
            .O(N__88324),
            .I(N__88317));
    InMux I__21132 (
            .O(N__88323),
            .I(N__88314));
    InMux I__21131 (
            .O(N__88322),
            .I(N__88311));
    InMux I__21130 (
            .O(N__88321),
            .I(N__88308));
    InMux I__21129 (
            .O(N__88320),
            .I(N__88302));
    LocalMux I__21128 (
            .O(N__88317),
            .I(N__88297));
    LocalMux I__21127 (
            .O(N__88314),
            .I(N__88297));
    LocalMux I__21126 (
            .O(N__88311),
            .I(N__88294));
    LocalMux I__21125 (
            .O(N__88308),
            .I(N__88291));
    InMux I__21124 (
            .O(N__88307),
            .I(N__88288));
    InMux I__21123 (
            .O(N__88306),
            .I(N__88285));
    InMux I__21122 (
            .O(N__88305),
            .I(N__88282));
    LocalMux I__21121 (
            .O(N__88302),
            .I(N__88275));
    Span4Mux_v I__21120 (
            .O(N__88297),
            .I(N__88275));
    Span4Mux_h I__21119 (
            .O(N__88294),
            .I(N__88270));
    Span4Mux_v I__21118 (
            .O(N__88291),
            .I(N__88270));
    LocalMux I__21117 (
            .O(N__88288),
            .I(N__88267));
    LocalMux I__21116 (
            .O(N__88285),
            .I(N__88264));
    LocalMux I__21115 (
            .O(N__88282),
            .I(N__88257));
    InMux I__21114 (
            .O(N__88281),
            .I(N__88251));
    InMux I__21113 (
            .O(N__88280),
            .I(N__88248));
    Span4Mux_v I__21112 (
            .O(N__88275),
            .I(N__88245));
    Span4Mux_v I__21111 (
            .O(N__88270),
            .I(N__88242));
    Span4Mux_v I__21110 (
            .O(N__88267),
            .I(N__88239));
    Span4Mux_v I__21109 (
            .O(N__88264),
            .I(N__88236));
    InMux I__21108 (
            .O(N__88263),
            .I(N__88231));
    InMux I__21107 (
            .O(N__88262),
            .I(N__88231));
    InMux I__21106 (
            .O(N__88261),
            .I(N__88228));
    InMux I__21105 (
            .O(N__88260),
            .I(N__88225));
    Span4Mux_h I__21104 (
            .O(N__88257),
            .I(N__88222));
    InMux I__21103 (
            .O(N__88256),
            .I(N__88219));
    CascadeMux I__21102 (
            .O(N__88255),
            .I(N__88216));
    InMux I__21101 (
            .O(N__88254),
            .I(N__88213));
    LocalMux I__21100 (
            .O(N__88251),
            .I(N__88210));
    LocalMux I__21099 (
            .O(N__88248),
            .I(N__88207));
    Sp12to4 I__21098 (
            .O(N__88245),
            .I(N__88202));
    Sp12to4 I__21097 (
            .O(N__88242),
            .I(N__88202));
    Span4Mux_v I__21096 (
            .O(N__88239),
            .I(N__88195));
    Span4Mux_v I__21095 (
            .O(N__88236),
            .I(N__88195));
    LocalMux I__21094 (
            .O(N__88231),
            .I(N__88195));
    LocalMux I__21093 (
            .O(N__88228),
            .I(N__88191));
    LocalMux I__21092 (
            .O(N__88225),
            .I(N__88186));
    Span4Mux_h I__21091 (
            .O(N__88222),
            .I(N__88186));
    LocalMux I__21090 (
            .O(N__88219),
            .I(N__88183));
    InMux I__21089 (
            .O(N__88216),
            .I(N__88180));
    LocalMux I__21088 (
            .O(N__88213),
            .I(N__88175));
    Span4Mux_v I__21087 (
            .O(N__88210),
            .I(N__88175));
    Span12Mux_s9_h I__21086 (
            .O(N__88207),
            .I(N__88170));
    Span12Mux_h I__21085 (
            .O(N__88202),
            .I(N__88170));
    Span4Mux_h I__21084 (
            .O(N__88195),
            .I(N__88167));
    InMux I__21083 (
            .O(N__88194),
            .I(N__88164));
    Span4Mux_h I__21082 (
            .O(N__88191),
            .I(N__88157));
    Span4Mux_v I__21081 (
            .O(N__88186),
            .I(N__88157));
    Span4Mux_v I__21080 (
            .O(N__88183),
            .I(N__88157));
    LocalMux I__21079 (
            .O(N__88180),
            .I(uart_pc_data_0));
    Odrv4 I__21078 (
            .O(N__88175),
            .I(uart_pc_data_0));
    Odrv12 I__21077 (
            .O(N__88170),
            .I(uart_pc_data_0));
    Odrv4 I__21076 (
            .O(N__88167),
            .I(uart_pc_data_0));
    LocalMux I__21075 (
            .O(N__88164),
            .I(uart_pc_data_0));
    Odrv4 I__21074 (
            .O(N__88157),
            .I(uart_pc_data_0));
    InMux I__21073 (
            .O(N__88144),
            .I(N__88141));
    LocalMux I__21072 (
            .O(N__88141),
            .I(N__88137));
    InMux I__21071 (
            .O(N__88140),
            .I(N__88134));
    Span4Mux_s2_h I__21070 (
            .O(N__88137),
            .I(N__88131));
    LocalMux I__21069 (
            .O(N__88134),
            .I(N__88128));
    Span4Mux_v I__21068 (
            .O(N__88131),
            .I(N__88123));
    Span4Mux_s2_h I__21067 (
            .O(N__88128),
            .I(N__88123));
    Odrv4 I__21066 (
            .O(N__88123),
            .I(xy_kd_0));
    CEMux I__21065 (
            .O(N__88120),
            .I(N__88116));
    CEMux I__21064 (
            .O(N__88119),
            .I(N__88113));
    LocalMux I__21063 (
            .O(N__88116),
            .I(N__88108));
    LocalMux I__21062 (
            .O(N__88113),
            .I(N__88108));
    Span4Mux_v I__21061 (
            .O(N__88108),
            .I(N__88103));
    CEMux I__21060 (
            .O(N__88107),
            .I(N__88100));
    CEMux I__21059 (
            .O(N__88106),
            .I(N__88097));
    Span4Mux_h I__21058 (
            .O(N__88103),
            .I(N__88092));
    LocalMux I__21057 (
            .O(N__88100),
            .I(N__88092));
    LocalMux I__21056 (
            .O(N__88097),
            .I(N__88084));
    Span4Mux_v I__21055 (
            .O(N__88092),
            .I(N__88081));
    CEMux I__21054 (
            .O(N__88091),
            .I(N__88075));
    CEMux I__21053 (
            .O(N__88090),
            .I(N__88072));
    CEMux I__21052 (
            .O(N__88089),
            .I(N__88069));
    CEMux I__21051 (
            .O(N__88088),
            .I(N__88066));
    CEMux I__21050 (
            .O(N__88087),
            .I(N__88063));
    Span4Mux_v I__21049 (
            .O(N__88084),
            .I(N__88058));
    Span4Mux_h I__21048 (
            .O(N__88081),
            .I(N__88058));
    CEMux I__21047 (
            .O(N__88080),
            .I(N__88055));
    CEMux I__21046 (
            .O(N__88079),
            .I(N__88050));
    CEMux I__21045 (
            .O(N__88078),
            .I(N__88047));
    LocalMux I__21044 (
            .O(N__88075),
            .I(N__88044));
    LocalMux I__21043 (
            .O(N__88072),
            .I(N__88041));
    LocalMux I__21042 (
            .O(N__88069),
            .I(N__88038));
    LocalMux I__21041 (
            .O(N__88066),
            .I(N__88035));
    LocalMux I__21040 (
            .O(N__88063),
            .I(N__88032));
    Span4Mux_h I__21039 (
            .O(N__88058),
            .I(N__88027));
    LocalMux I__21038 (
            .O(N__88055),
            .I(N__88027));
    CEMux I__21037 (
            .O(N__88054),
            .I(N__88024));
    CEMux I__21036 (
            .O(N__88053),
            .I(N__88021));
    LocalMux I__21035 (
            .O(N__88050),
            .I(N__88017));
    LocalMux I__21034 (
            .O(N__88047),
            .I(N__88014));
    Span4Mux_s3_h I__21033 (
            .O(N__88044),
            .I(N__88009));
    Span4Mux_h I__21032 (
            .O(N__88041),
            .I(N__88009));
    Span4Mux_v I__21031 (
            .O(N__88038),
            .I(N__87998));
    Span4Mux_v I__21030 (
            .O(N__88035),
            .I(N__87998));
    Span4Mux_v I__21029 (
            .O(N__88032),
            .I(N__87998));
    Span4Mux_h I__21028 (
            .O(N__88027),
            .I(N__87998));
    LocalMux I__21027 (
            .O(N__88024),
            .I(N__87998));
    LocalMux I__21026 (
            .O(N__88021),
            .I(N__87995));
    CEMux I__21025 (
            .O(N__88020),
            .I(N__87992));
    Span4Mux_v I__21024 (
            .O(N__88017),
            .I(N__87988));
    Span4Mux_v I__21023 (
            .O(N__88014),
            .I(N__87983));
    Span4Mux_h I__21022 (
            .O(N__88009),
            .I(N__87983));
    Sp12to4 I__21021 (
            .O(N__87998),
            .I(N__87980));
    Span4Mux_v I__21020 (
            .O(N__87995),
            .I(N__87975));
    LocalMux I__21019 (
            .O(N__87992),
            .I(N__87975));
    CEMux I__21018 (
            .O(N__87991),
            .I(N__87972));
    Odrv4 I__21017 (
            .O(N__87988),
            .I(\pid_side.N_834_0 ));
    Odrv4 I__21016 (
            .O(N__87983),
            .I(\pid_side.N_834_0 ));
    Odrv12 I__21015 (
            .O(N__87980),
            .I(\pid_side.N_834_0 ));
    Odrv4 I__21014 (
            .O(N__87975),
            .I(\pid_side.N_834_0 ));
    LocalMux I__21013 (
            .O(N__87972),
            .I(\pid_side.N_834_0 ));
    SRMux I__21012 (
            .O(N__87961),
            .I(N__87955));
    InMux I__21011 (
            .O(N__87960),
            .I(N__87955));
    LocalMux I__21010 (
            .O(N__87955),
            .I(N__87937));
    SRMux I__21009 (
            .O(N__87954),
            .I(N__87904));
    SRMux I__21008 (
            .O(N__87953),
            .I(N__87904));
    SRMux I__21007 (
            .O(N__87952),
            .I(N__87904));
    SRMux I__21006 (
            .O(N__87951),
            .I(N__87904));
    SRMux I__21005 (
            .O(N__87950),
            .I(N__87904));
    SRMux I__21004 (
            .O(N__87949),
            .I(N__87904));
    SRMux I__21003 (
            .O(N__87948),
            .I(N__87904));
    SRMux I__21002 (
            .O(N__87947),
            .I(N__87904));
    SRMux I__21001 (
            .O(N__87946),
            .I(N__87904));
    SRMux I__21000 (
            .O(N__87945),
            .I(N__87904));
    SRMux I__20999 (
            .O(N__87944),
            .I(N__87904));
    SRMux I__20998 (
            .O(N__87943),
            .I(N__87904));
    SRMux I__20997 (
            .O(N__87942),
            .I(N__87904));
    SRMux I__20996 (
            .O(N__87941),
            .I(N__87904));
    SRMux I__20995 (
            .O(N__87940),
            .I(N__87904));
    Glb2LocalMux I__20994 (
            .O(N__87937),
            .I(N__87904));
    GlobalMux I__20993 (
            .O(N__87904),
            .I(N__87901));
    gio2CtrlBuf I__20992 (
            .O(N__87901),
            .I(\pid_side.N_2054_g ));
    InMux I__20991 (
            .O(N__87898),
            .I(N__87895));
    LocalMux I__20990 (
            .O(N__87895),
            .I(N__87892));
    Span4Mux_h I__20989 (
            .O(N__87892),
            .I(N__87889));
    Span4Mux_v I__20988 (
            .O(N__87889),
            .I(N__87886));
    Odrv4 I__20987 (
            .O(N__87886),
            .I(\pid_side.O_1_7 ));
    InMux I__20986 (
            .O(N__87883),
            .I(N__87874));
    InMux I__20985 (
            .O(N__87882),
            .I(N__87874));
    InMux I__20984 (
            .O(N__87881),
            .I(N__87874));
    LocalMux I__20983 (
            .O(N__87874),
            .I(N__87871));
    Odrv4 I__20982 (
            .O(N__87871),
            .I(\pid_side.error_d_regZ0Z_4 ));
    InMux I__20981 (
            .O(N__87868),
            .I(N__87864));
    InMux I__20980 (
            .O(N__87867),
            .I(N__87861));
    LocalMux I__20979 (
            .O(N__87864),
            .I(N__87856));
    LocalMux I__20978 (
            .O(N__87861),
            .I(N__87856));
    Odrv4 I__20977 (
            .O(N__87856),
            .I(\pid_side.error_d_reg_prevZ0Z_18 ));
    InMux I__20976 (
            .O(N__87853),
            .I(N__87850));
    LocalMux I__20975 (
            .O(N__87850),
            .I(N__87846));
    InMux I__20974 (
            .O(N__87849),
            .I(N__87843));
    Span12Mux_s8_v I__20973 (
            .O(N__87846),
            .I(N__87838));
    LocalMux I__20972 (
            .O(N__87843),
            .I(N__87838));
    Odrv12 I__20971 (
            .O(N__87838),
            .I(\pid_side.error_d_reg_prev_esr_RNIH7JO_0Z0Z_18 ));
    InMux I__20970 (
            .O(N__87835),
            .I(N__87832));
    LocalMux I__20969 (
            .O(N__87832),
            .I(N__87829));
    Span4Mux_h I__20968 (
            .O(N__87829),
            .I(N__87826));
    Odrv4 I__20967 (
            .O(N__87826),
            .I(\pid_side.O_2_12 ));
    InMux I__20966 (
            .O(N__87823),
            .I(N__87817));
    InMux I__20965 (
            .O(N__87822),
            .I(N__87817));
    LocalMux I__20964 (
            .O(N__87817),
            .I(N__87814));
    Span4Mux_h I__20963 (
            .O(N__87814),
            .I(N__87811));
    Span4Mux_h I__20962 (
            .O(N__87811),
            .I(N__87808));
    Odrv4 I__20961 (
            .O(N__87808),
            .I(\pid_side.error_p_regZ0Z_8 ));
    CascadeMux I__20960 (
            .O(N__87805),
            .I(N__87797));
    InMux I__20959 (
            .O(N__87804),
            .I(N__87794));
    CascadeMux I__20958 (
            .O(N__87803),
            .I(N__87791));
    CascadeMux I__20957 (
            .O(N__87802),
            .I(N__87787));
    InMux I__20956 (
            .O(N__87801),
            .I(N__87784));
    InMux I__20955 (
            .O(N__87800),
            .I(N__87781));
    InMux I__20954 (
            .O(N__87797),
            .I(N__87770));
    LocalMux I__20953 (
            .O(N__87794),
            .I(N__87767));
    InMux I__20952 (
            .O(N__87791),
            .I(N__87764));
    InMux I__20951 (
            .O(N__87790),
            .I(N__87761));
    InMux I__20950 (
            .O(N__87787),
            .I(N__87757));
    LocalMux I__20949 (
            .O(N__87784),
            .I(N__87752));
    LocalMux I__20948 (
            .O(N__87781),
            .I(N__87752));
    InMux I__20947 (
            .O(N__87780),
            .I(N__87746));
    InMux I__20946 (
            .O(N__87779),
            .I(N__87741));
    InMux I__20945 (
            .O(N__87778),
            .I(N__87741));
    InMux I__20944 (
            .O(N__87777),
            .I(N__87738));
    InMux I__20943 (
            .O(N__87776),
            .I(N__87733));
    InMux I__20942 (
            .O(N__87775),
            .I(N__87733));
    CascadeMux I__20941 (
            .O(N__87774),
            .I(N__87730));
    InMux I__20940 (
            .O(N__87773),
            .I(N__87727));
    LocalMux I__20939 (
            .O(N__87770),
            .I(N__87724));
    Span4Mux_v I__20938 (
            .O(N__87767),
            .I(N__87719));
    LocalMux I__20937 (
            .O(N__87764),
            .I(N__87719));
    LocalMux I__20936 (
            .O(N__87761),
            .I(N__87716));
    InMux I__20935 (
            .O(N__87760),
            .I(N__87713));
    LocalMux I__20934 (
            .O(N__87757),
            .I(N__87710));
    Span4Mux_v I__20933 (
            .O(N__87752),
            .I(N__87707));
    InMux I__20932 (
            .O(N__87751),
            .I(N__87704));
    InMux I__20931 (
            .O(N__87750),
            .I(N__87701));
    InMux I__20930 (
            .O(N__87749),
            .I(N__87698));
    LocalMux I__20929 (
            .O(N__87746),
            .I(N__87695));
    LocalMux I__20928 (
            .O(N__87741),
            .I(N__87692));
    LocalMux I__20927 (
            .O(N__87738),
            .I(N__87687));
    LocalMux I__20926 (
            .O(N__87733),
            .I(N__87687));
    InMux I__20925 (
            .O(N__87730),
            .I(N__87684));
    LocalMux I__20924 (
            .O(N__87727),
            .I(N__87681));
    Span4Mux_v I__20923 (
            .O(N__87724),
            .I(N__87676));
    Span4Mux_v I__20922 (
            .O(N__87719),
            .I(N__87676));
    Span4Mux_h I__20921 (
            .O(N__87716),
            .I(N__87671));
    LocalMux I__20920 (
            .O(N__87713),
            .I(N__87668));
    Span4Mux_h I__20919 (
            .O(N__87710),
            .I(N__87660));
    Span4Mux_v I__20918 (
            .O(N__87707),
            .I(N__87660));
    LocalMux I__20917 (
            .O(N__87704),
            .I(N__87660));
    LocalMux I__20916 (
            .O(N__87701),
            .I(N__87653));
    LocalMux I__20915 (
            .O(N__87698),
            .I(N__87653));
    Span4Mux_h I__20914 (
            .O(N__87695),
            .I(N__87653));
    Span4Mux_h I__20913 (
            .O(N__87692),
            .I(N__87648));
    Span4Mux_v I__20912 (
            .O(N__87687),
            .I(N__87648));
    LocalMux I__20911 (
            .O(N__87684),
            .I(N__87641));
    Span4Mux_v I__20910 (
            .O(N__87681),
            .I(N__87641));
    Span4Mux_h I__20909 (
            .O(N__87676),
            .I(N__87641));
    InMux I__20908 (
            .O(N__87675),
            .I(N__87638));
    InMux I__20907 (
            .O(N__87674),
            .I(N__87635));
    Span4Mux_h I__20906 (
            .O(N__87671),
            .I(N__87630));
    Span4Mux_h I__20905 (
            .O(N__87668),
            .I(N__87630));
    InMux I__20904 (
            .O(N__87667),
            .I(N__87627));
    Span4Mux_h I__20903 (
            .O(N__87660),
            .I(N__87624));
    Span4Mux_v I__20902 (
            .O(N__87653),
            .I(N__87619));
    Span4Mux_h I__20901 (
            .O(N__87648),
            .I(N__87619));
    Span4Mux_h I__20900 (
            .O(N__87641),
            .I(N__87616));
    LocalMux I__20899 (
            .O(N__87638),
            .I(pid_side_N_164));
    LocalMux I__20898 (
            .O(N__87635),
            .I(pid_side_N_164));
    Odrv4 I__20897 (
            .O(N__87630),
            .I(pid_side_N_164));
    LocalMux I__20896 (
            .O(N__87627),
            .I(pid_side_N_164));
    Odrv4 I__20895 (
            .O(N__87624),
            .I(pid_side_N_164));
    Odrv4 I__20894 (
            .O(N__87619),
            .I(pid_side_N_164));
    Odrv4 I__20893 (
            .O(N__87616),
            .I(pid_side_N_164));
    InMux I__20892 (
            .O(N__87601),
            .I(N__87597));
    InMux I__20891 (
            .O(N__87600),
            .I(N__87594));
    LocalMux I__20890 (
            .O(N__87597),
            .I(N__87590));
    LocalMux I__20889 (
            .O(N__87594),
            .I(N__87587));
    InMux I__20888 (
            .O(N__87593),
            .I(N__87583));
    Span4Mux_s3_h I__20887 (
            .O(N__87590),
            .I(N__87580));
    Span4Mux_v I__20886 (
            .O(N__87587),
            .I(N__87577));
    InMux I__20885 (
            .O(N__87586),
            .I(N__87574));
    LocalMux I__20884 (
            .O(N__87583),
            .I(\pid_side.N_589 ));
    Odrv4 I__20883 (
            .O(N__87580),
            .I(\pid_side.N_589 ));
    Odrv4 I__20882 (
            .O(N__87577),
            .I(\pid_side.N_589 ));
    LocalMux I__20881 (
            .O(N__87574),
            .I(\pid_side.N_589 ));
    CascadeMux I__20880 (
            .O(N__87565),
            .I(\pid_side.N_459_cascade_ ));
    InMux I__20879 (
            .O(N__87562),
            .I(N__87555));
    InMux I__20878 (
            .O(N__87561),
            .I(N__87551));
    InMux I__20877 (
            .O(N__87560),
            .I(N__87547));
    InMux I__20876 (
            .O(N__87559),
            .I(N__87544));
    InMux I__20875 (
            .O(N__87558),
            .I(N__87541));
    LocalMux I__20874 (
            .O(N__87555),
            .I(N__87537));
    InMux I__20873 (
            .O(N__87554),
            .I(N__87534));
    LocalMux I__20872 (
            .O(N__87551),
            .I(N__87530));
    InMux I__20871 (
            .O(N__87550),
            .I(N__87526));
    LocalMux I__20870 (
            .O(N__87547),
            .I(N__87523));
    LocalMux I__20869 (
            .O(N__87544),
            .I(N__87518));
    LocalMux I__20868 (
            .O(N__87541),
            .I(N__87518));
    InMux I__20867 (
            .O(N__87540),
            .I(N__87515));
    Span4Mux_s1_h I__20866 (
            .O(N__87537),
            .I(N__87512));
    LocalMux I__20865 (
            .O(N__87534),
            .I(N__87509));
    InMux I__20864 (
            .O(N__87533),
            .I(N__87506));
    Span4Mux_s1_h I__20863 (
            .O(N__87530),
            .I(N__87503));
    InMux I__20862 (
            .O(N__87529),
            .I(N__87500));
    LocalMux I__20861 (
            .O(N__87526),
            .I(N__87495));
    Span4Mux_v I__20860 (
            .O(N__87523),
            .I(N__87495));
    Span4Mux_v I__20859 (
            .O(N__87518),
            .I(N__87490));
    LocalMux I__20858 (
            .O(N__87515),
            .I(N__87490));
    Span4Mux_v I__20857 (
            .O(N__87512),
            .I(N__87487));
    Span4Mux_h I__20856 (
            .O(N__87509),
            .I(N__87480));
    LocalMux I__20855 (
            .O(N__87506),
            .I(N__87480));
    Span4Mux_h I__20854 (
            .O(N__87503),
            .I(N__87480));
    LocalMux I__20853 (
            .O(N__87500),
            .I(\pid_side.error_11 ));
    Odrv4 I__20852 (
            .O(N__87495),
            .I(\pid_side.error_11 ));
    Odrv4 I__20851 (
            .O(N__87490),
            .I(\pid_side.error_11 ));
    Odrv4 I__20850 (
            .O(N__87487),
            .I(\pid_side.error_11 ));
    Odrv4 I__20849 (
            .O(N__87480),
            .I(\pid_side.error_11 ));
    InMux I__20848 (
            .O(N__87469),
            .I(N__87465));
    InMux I__20847 (
            .O(N__87468),
            .I(N__87462));
    LocalMux I__20846 (
            .O(N__87465),
            .I(N__87456));
    LocalMux I__20845 (
            .O(N__87462),
            .I(N__87456));
    InMux I__20844 (
            .O(N__87461),
            .I(N__87453));
    Odrv12 I__20843 (
            .O(N__87456),
            .I(\pid_side.N_225 ));
    LocalMux I__20842 (
            .O(N__87453),
            .I(\pid_side.N_225 ));
    CascadeMux I__20841 (
            .O(N__87448),
            .I(N__87444));
    InMux I__20840 (
            .O(N__87447),
            .I(N__87440));
    InMux I__20839 (
            .O(N__87444),
            .I(N__87437));
    CascadeMux I__20838 (
            .O(N__87443),
            .I(N__87431));
    LocalMux I__20837 (
            .O(N__87440),
            .I(N__87423));
    LocalMux I__20836 (
            .O(N__87437),
            .I(N__87423));
    CascadeMux I__20835 (
            .O(N__87436),
            .I(N__87419));
    InMux I__20834 (
            .O(N__87435),
            .I(N__87411));
    InMux I__20833 (
            .O(N__87434),
            .I(N__87411));
    InMux I__20832 (
            .O(N__87431),
            .I(N__87405));
    CascadeMux I__20831 (
            .O(N__87430),
            .I(N__87400));
    InMux I__20830 (
            .O(N__87429),
            .I(N__87396));
    InMux I__20829 (
            .O(N__87428),
            .I(N__87393));
    Span4Mux_v I__20828 (
            .O(N__87423),
            .I(N__87390));
    InMux I__20827 (
            .O(N__87422),
            .I(N__87383));
    InMux I__20826 (
            .O(N__87419),
            .I(N__87383));
    InMux I__20825 (
            .O(N__87418),
            .I(N__87380));
    CascadeMux I__20824 (
            .O(N__87417),
            .I(N__87377));
    CascadeMux I__20823 (
            .O(N__87416),
            .I(N__87371));
    LocalMux I__20822 (
            .O(N__87411),
            .I(N__87368));
    InMux I__20821 (
            .O(N__87410),
            .I(N__87365));
    InMux I__20820 (
            .O(N__87409),
            .I(N__87362));
    InMux I__20819 (
            .O(N__87408),
            .I(N__87359));
    LocalMux I__20818 (
            .O(N__87405),
            .I(N__87355));
    CascadeMux I__20817 (
            .O(N__87404),
            .I(N__87352));
    InMux I__20816 (
            .O(N__87403),
            .I(N__87349));
    InMux I__20815 (
            .O(N__87400),
            .I(N__87343));
    InMux I__20814 (
            .O(N__87399),
            .I(N__87343));
    LocalMux I__20813 (
            .O(N__87396),
            .I(N__87340));
    LocalMux I__20812 (
            .O(N__87393),
            .I(N__87337));
    Span4Mux_h I__20811 (
            .O(N__87390),
            .I(N__87334));
    InMux I__20810 (
            .O(N__87389),
            .I(N__87331));
    InMux I__20809 (
            .O(N__87388),
            .I(N__87326));
    LocalMux I__20808 (
            .O(N__87383),
            .I(N__87321));
    LocalMux I__20807 (
            .O(N__87380),
            .I(N__87321));
    InMux I__20806 (
            .O(N__87377),
            .I(N__87318));
    InMux I__20805 (
            .O(N__87376),
            .I(N__87313));
    InMux I__20804 (
            .O(N__87375),
            .I(N__87313));
    InMux I__20803 (
            .O(N__87374),
            .I(N__87308));
    InMux I__20802 (
            .O(N__87371),
            .I(N__87308));
    Span4Mux_h I__20801 (
            .O(N__87368),
            .I(N__87301));
    LocalMux I__20800 (
            .O(N__87365),
            .I(N__87301));
    LocalMux I__20799 (
            .O(N__87362),
            .I(N__87301));
    LocalMux I__20798 (
            .O(N__87359),
            .I(N__87298));
    CascadeMux I__20797 (
            .O(N__87358),
            .I(N__87295));
    Span4Mux_v I__20796 (
            .O(N__87355),
            .I(N__87292));
    InMux I__20795 (
            .O(N__87352),
            .I(N__87289));
    LocalMux I__20794 (
            .O(N__87349),
            .I(N__87286));
    InMux I__20793 (
            .O(N__87348),
            .I(N__87283));
    LocalMux I__20792 (
            .O(N__87343),
            .I(N__87280));
    Span4Mux_v I__20791 (
            .O(N__87340),
            .I(N__87273));
    Span4Mux_v I__20790 (
            .O(N__87337),
            .I(N__87273));
    Sp12to4 I__20789 (
            .O(N__87334),
            .I(N__87265));
    LocalMux I__20788 (
            .O(N__87331),
            .I(N__87265));
    CascadeMux I__20787 (
            .O(N__87330),
            .I(N__87262));
    CascadeMux I__20786 (
            .O(N__87329),
            .I(N__87259));
    LocalMux I__20785 (
            .O(N__87326),
            .I(N__87253));
    Span4Mux_v I__20784 (
            .O(N__87321),
            .I(N__87253));
    LocalMux I__20783 (
            .O(N__87318),
            .I(N__87242));
    LocalMux I__20782 (
            .O(N__87313),
            .I(N__87242));
    LocalMux I__20781 (
            .O(N__87308),
            .I(N__87242));
    Span4Mux_v I__20780 (
            .O(N__87301),
            .I(N__87242));
    Span4Mux_v I__20779 (
            .O(N__87298),
            .I(N__87242));
    InMux I__20778 (
            .O(N__87295),
            .I(N__87239));
    Span4Mux_h I__20777 (
            .O(N__87292),
            .I(N__87230));
    LocalMux I__20776 (
            .O(N__87289),
            .I(N__87230));
    Span4Mux_h I__20775 (
            .O(N__87286),
            .I(N__87230));
    LocalMux I__20774 (
            .O(N__87283),
            .I(N__87230));
    Span4Mux_h I__20773 (
            .O(N__87280),
            .I(N__87227));
    InMux I__20772 (
            .O(N__87279),
            .I(N__87224));
    InMux I__20771 (
            .O(N__87278),
            .I(N__87221));
    Span4Mux_h I__20770 (
            .O(N__87273),
            .I(N__87218));
    InMux I__20769 (
            .O(N__87272),
            .I(N__87213));
    InMux I__20768 (
            .O(N__87271),
            .I(N__87213));
    InMux I__20767 (
            .O(N__87270),
            .I(N__87210));
    Span12Mux_h I__20766 (
            .O(N__87265),
            .I(N__87207));
    InMux I__20765 (
            .O(N__87262),
            .I(N__87200));
    InMux I__20764 (
            .O(N__87259),
            .I(N__87200));
    InMux I__20763 (
            .O(N__87258),
            .I(N__87200));
    Sp12to4 I__20762 (
            .O(N__87253),
            .I(N__87195));
    Sp12to4 I__20761 (
            .O(N__87242),
            .I(N__87195));
    LocalMux I__20760 (
            .O(N__87239),
            .I(N__87188));
    Span4Mux_v I__20759 (
            .O(N__87230),
            .I(N__87188));
    Span4Mux_v I__20758 (
            .O(N__87227),
            .I(N__87188));
    LocalMux I__20757 (
            .O(N__87224),
            .I(xy_ki_1));
    LocalMux I__20756 (
            .O(N__87221),
            .I(xy_ki_1));
    Odrv4 I__20755 (
            .O(N__87218),
            .I(xy_ki_1));
    LocalMux I__20754 (
            .O(N__87213),
            .I(xy_ki_1));
    LocalMux I__20753 (
            .O(N__87210),
            .I(xy_ki_1));
    Odrv12 I__20752 (
            .O(N__87207),
            .I(xy_ki_1));
    LocalMux I__20751 (
            .O(N__87200),
            .I(xy_ki_1));
    Odrv12 I__20750 (
            .O(N__87195),
            .I(xy_ki_1));
    Odrv4 I__20749 (
            .O(N__87188),
            .I(xy_ki_1));
    CascadeMux I__20748 (
            .O(N__87169),
            .I(\pid_side.m23_2_03_0_2_cascade_ ));
    InMux I__20747 (
            .O(N__87166),
            .I(N__87160));
    InMux I__20746 (
            .O(N__87165),
            .I(N__87160));
    LocalMux I__20745 (
            .O(N__87160),
            .I(\pid_side.un4_error_i_reg_29_ns_sn ));
    CascadeMux I__20744 (
            .O(N__87157),
            .I(N__87154));
    InMux I__20743 (
            .O(N__87154),
            .I(N__87148));
    InMux I__20742 (
            .O(N__87153),
            .I(N__87148));
    LocalMux I__20741 (
            .O(N__87148),
            .I(\pid_side.un4_error_i_reg_29_ns_rn_0 ));
    CascadeMux I__20740 (
            .O(N__87145),
            .I(N__87135));
    CascadeMux I__20739 (
            .O(N__87144),
            .I(N__87132));
    InMux I__20738 (
            .O(N__87143),
            .I(N__87129));
    CascadeMux I__20737 (
            .O(N__87142),
            .I(N__87125));
    InMux I__20736 (
            .O(N__87141),
            .I(N__87118));
    InMux I__20735 (
            .O(N__87140),
            .I(N__87118));
    InMux I__20734 (
            .O(N__87139),
            .I(N__87118));
    InMux I__20733 (
            .O(N__87138),
            .I(N__87115));
    InMux I__20732 (
            .O(N__87135),
            .I(N__87110));
    InMux I__20731 (
            .O(N__87132),
            .I(N__87107));
    LocalMux I__20730 (
            .O(N__87129),
            .I(N__87099));
    CascadeMux I__20729 (
            .O(N__87128),
            .I(N__87095));
    InMux I__20728 (
            .O(N__87125),
            .I(N__87090));
    LocalMux I__20727 (
            .O(N__87118),
            .I(N__87083));
    LocalMux I__20726 (
            .O(N__87115),
            .I(N__87083));
    InMux I__20725 (
            .O(N__87114),
            .I(N__87080));
    InMux I__20724 (
            .O(N__87113),
            .I(N__87077));
    LocalMux I__20723 (
            .O(N__87110),
            .I(N__87074));
    LocalMux I__20722 (
            .O(N__87107),
            .I(N__87069));
    InMux I__20721 (
            .O(N__87106),
            .I(N__87064));
    InMux I__20720 (
            .O(N__87105),
            .I(N__87064));
    InMux I__20719 (
            .O(N__87104),
            .I(N__87061));
    InMux I__20718 (
            .O(N__87103),
            .I(N__87056));
    InMux I__20717 (
            .O(N__87102),
            .I(N__87056));
    Span4Mux_v I__20716 (
            .O(N__87099),
            .I(N__87052));
    InMux I__20715 (
            .O(N__87098),
            .I(N__87049));
    InMux I__20714 (
            .O(N__87095),
            .I(N__87044));
    InMux I__20713 (
            .O(N__87094),
            .I(N__87039));
    InMux I__20712 (
            .O(N__87093),
            .I(N__87039));
    LocalMux I__20711 (
            .O(N__87090),
            .I(N__87036));
    CascadeMux I__20710 (
            .O(N__87089),
            .I(N__87027));
    InMux I__20709 (
            .O(N__87088),
            .I(N__87022));
    Span4Mux_v I__20708 (
            .O(N__87083),
            .I(N__87019));
    LocalMux I__20707 (
            .O(N__87080),
            .I(N__87014));
    LocalMux I__20706 (
            .O(N__87077),
            .I(N__87014));
    Span4Mux_h I__20705 (
            .O(N__87074),
            .I(N__87011));
    InMux I__20704 (
            .O(N__87073),
            .I(N__87006));
    InMux I__20703 (
            .O(N__87072),
            .I(N__87006));
    Span4Mux_v I__20702 (
            .O(N__87069),
            .I(N__87001));
    LocalMux I__20701 (
            .O(N__87064),
            .I(N__87001));
    LocalMux I__20700 (
            .O(N__87061),
            .I(N__86996));
    LocalMux I__20699 (
            .O(N__87056),
            .I(N__86996));
    CascadeMux I__20698 (
            .O(N__87055),
            .I(N__86993));
    Span4Mux_h I__20697 (
            .O(N__87052),
            .I(N__86985));
    LocalMux I__20696 (
            .O(N__87049),
            .I(N__86985));
    InMux I__20695 (
            .O(N__87048),
            .I(N__86982));
    InMux I__20694 (
            .O(N__87047),
            .I(N__86979));
    LocalMux I__20693 (
            .O(N__87044),
            .I(N__86972));
    LocalMux I__20692 (
            .O(N__87039),
            .I(N__86972));
    Span4Mux_h I__20691 (
            .O(N__87036),
            .I(N__86972));
    InMux I__20690 (
            .O(N__87035),
            .I(N__86967));
    InMux I__20689 (
            .O(N__87034),
            .I(N__86958));
    InMux I__20688 (
            .O(N__87033),
            .I(N__86958));
    InMux I__20687 (
            .O(N__87032),
            .I(N__86958));
    InMux I__20686 (
            .O(N__87031),
            .I(N__86958));
    InMux I__20685 (
            .O(N__87030),
            .I(N__86953));
    InMux I__20684 (
            .O(N__87027),
            .I(N__86953));
    InMux I__20683 (
            .O(N__87026),
            .I(N__86948));
    InMux I__20682 (
            .O(N__87025),
            .I(N__86948));
    LocalMux I__20681 (
            .O(N__87022),
            .I(N__86941));
    Span4Mux_h I__20680 (
            .O(N__87019),
            .I(N__86941));
    Span4Mux_v I__20679 (
            .O(N__87014),
            .I(N__86941));
    Span4Mux_v I__20678 (
            .O(N__87011),
            .I(N__86927));
    LocalMux I__20677 (
            .O(N__87006),
            .I(N__86927));
    Span4Mux_h I__20676 (
            .O(N__87001),
            .I(N__86927));
    Span4Mux_v I__20675 (
            .O(N__86996),
            .I(N__86924));
    InMux I__20674 (
            .O(N__86993),
            .I(N__86915));
    InMux I__20673 (
            .O(N__86992),
            .I(N__86915));
    InMux I__20672 (
            .O(N__86991),
            .I(N__86915));
    InMux I__20671 (
            .O(N__86990),
            .I(N__86915));
    Span4Mux_v I__20670 (
            .O(N__86985),
            .I(N__86912));
    LocalMux I__20669 (
            .O(N__86982),
            .I(N__86909));
    LocalMux I__20668 (
            .O(N__86979),
            .I(N__86904));
    Span4Mux_h I__20667 (
            .O(N__86972),
            .I(N__86904));
    InMux I__20666 (
            .O(N__86971),
            .I(N__86899));
    InMux I__20665 (
            .O(N__86970),
            .I(N__86896));
    LocalMux I__20664 (
            .O(N__86967),
            .I(N__86891));
    LocalMux I__20663 (
            .O(N__86958),
            .I(N__86891));
    LocalMux I__20662 (
            .O(N__86953),
            .I(N__86888));
    LocalMux I__20661 (
            .O(N__86948),
            .I(N__86883));
    Span4Mux_v I__20660 (
            .O(N__86941),
            .I(N__86883));
    InMux I__20659 (
            .O(N__86940),
            .I(N__86876));
    InMux I__20658 (
            .O(N__86939),
            .I(N__86876));
    InMux I__20657 (
            .O(N__86938),
            .I(N__86876));
    InMux I__20656 (
            .O(N__86937),
            .I(N__86871));
    InMux I__20655 (
            .O(N__86936),
            .I(N__86871));
    InMux I__20654 (
            .O(N__86935),
            .I(N__86868));
    InMux I__20653 (
            .O(N__86934),
            .I(N__86865));
    Span4Mux_h I__20652 (
            .O(N__86927),
            .I(N__86862));
    Span4Mux_h I__20651 (
            .O(N__86924),
            .I(N__86855));
    LocalMux I__20650 (
            .O(N__86915),
            .I(N__86855));
    Span4Mux_h I__20649 (
            .O(N__86912),
            .I(N__86855));
    Span4Mux_h I__20648 (
            .O(N__86909),
            .I(N__86850));
    Span4Mux_v I__20647 (
            .O(N__86904),
            .I(N__86850));
    InMux I__20646 (
            .O(N__86903),
            .I(N__86845));
    InMux I__20645 (
            .O(N__86902),
            .I(N__86845));
    LocalMux I__20644 (
            .O(N__86899),
            .I(N__86838));
    LocalMux I__20643 (
            .O(N__86896),
            .I(N__86838));
    Sp12to4 I__20642 (
            .O(N__86891),
            .I(N__86838));
    Span4Mux_h I__20641 (
            .O(N__86888),
            .I(N__86831));
    Span4Mux_h I__20640 (
            .O(N__86883),
            .I(N__86831));
    LocalMux I__20639 (
            .O(N__86876),
            .I(N__86831));
    LocalMux I__20638 (
            .O(N__86871),
            .I(pid_front_N_335));
    LocalMux I__20637 (
            .O(N__86868),
            .I(pid_front_N_335));
    LocalMux I__20636 (
            .O(N__86865),
            .I(pid_front_N_335));
    Odrv4 I__20635 (
            .O(N__86862),
            .I(pid_front_N_335));
    Odrv4 I__20634 (
            .O(N__86855),
            .I(pid_front_N_335));
    Odrv4 I__20633 (
            .O(N__86850),
            .I(pid_front_N_335));
    LocalMux I__20632 (
            .O(N__86845),
            .I(pid_front_N_335));
    Odrv12 I__20631 (
            .O(N__86838),
            .I(pid_front_N_335));
    Odrv4 I__20630 (
            .O(N__86831),
            .I(pid_front_N_335));
    InMux I__20629 (
            .O(N__86812),
            .I(N__86809));
    LocalMux I__20628 (
            .O(N__86809),
            .I(\pid_side.m23_2_03_0_1 ));
    CascadeMux I__20627 (
            .O(N__86806),
            .I(\pid_side.error_i_reg_esr_RNO_2Z0Z_19_cascade_ ));
    InMux I__20626 (
            .O(N__86803),
            .I(N__86800));
    LocalMux I__20625 (
            .O(N__86800),
            .I(\pid_side.error_i_reg_esr_RNO_1Z0Z_19 ));
    InMux I__20624 (
            .O(N__86797),
            .I(N__86794));
    LocalMux I__20623 (
            .O(N__86794),
            .I(N__86791));
    Span12Mux_h I__20622 (
            .O(N__86791),
            .I(N__86788));
    Odrv12 I__20621 (
            .O(N__86788),
            .I(\pid_side.error_i_regZ0Z_19 ));
    CEMux I__20620 (
            .O(N__86785),
            .I(N__86779));
    CEMux I__20619 (
            .O(N__86784),
            .I(N__86771));
    CEMux I__20618 (
            .O(N__86783),
            .I(N__86768));
    CEMux I__20617 (
            .O(N__86782),
            .I(N__86765));
    LocalMux I__20616 (
            .O(N__86779),
            .I(N__86762));
    CEMux I__20615 (
            .O(N__86778),
            .I(N__86756));
    CEMux I__20614 (
            .O(N__86777),
            .I(N__86752));
    CEMux I__20613 (
            .O(N__86776),
            .I(N__86748));
    CEMux I__20612 (
            .O(N__86775),
            .I(N__86745));
    CEMux I__20611 (
            .O(N__86774),
            .I(N__86741));
    LocalMux I__20610 (
            .O(N__86771),
            .I(N__86738));
    LocalMux I__20609 (
            .O(N__86768),
            .I(N__86735));
    LocalMux I__20608 (
            .O(N__86765),
            .I(N__86732));
    Span4Mux_h I__20607 (
            .O(N__86762),
            .I(N__86729));
    CEMux I__20606 (
            .O(N__86761),
            .I(N__86726));
    CEMux I__20605 (
            .O(N__86760),
            .I(N__86723));
    CEMux I__20604 (
            .O(N__86759),
            .I(N__86720));
    LocalMux I__20603 (
            .O(N__86756),
            .I(N__86717));
    CEMux I__20602 (
            .O(N__86755),
            .I(N__86714));
    LocalMux I__20601 (
            .O(N__86752),
            .I(N__86711));
    CEMux I__20600 (
            .O(N__86751),
            .I(N__86708));
    LocalMux I__20599 (
            .O(N__86748),
            .I(N__86705));
    LocalMux I__20598 (
            .O(N__86745),
            .I(N__86702));
    CEMux I__20597 (
            .O(N__86744),
            .I(N__86699));
    LocalMux I__20596 (
            .O(N__86741),
            .I(N__86694));
    Span4Mux_h I__20595 (
            .O(N__86738),
            .I(N__86694));
    Span4Mux_v I__20594 (
            .O(N__86735),
            .I(N__86689));
    Span4Mux_h I__20593 (
            .O(N__86732),
            .I(N__86689));
    Span4Mux_h I__20592 (
            .O(N__86729),
            .I(N__86686));
    LocalMux I__20591 (
            .O(N__86726),
            .I(N__86683));
    LocalMux I__20590 (
            .O(N__86723),
            .I(N__86680));
    LocalMux I__20589 (
            .O(N__86720),
            .I(N__86673));
    Span4Mux_h I__20588 (
            .O(N__86717),
            .I(N__86673));
    LocalMux I__20587 (
            .O(N__86714),
            .I(N__86673));
    Span4Mux_v I__20586 (
            .O(N__86711),
            .I(N__86668));
    LocalMux I__20585 (
            .O(N__86708),
            .I(N__86668));
    Span4Mux_h I__20584 (
            .O(N__86705),
            .I(N__86663));
    Span4Mux_h I__20583 (
            .O(N__86702),
            .I(N__86663));
    LocalMux I__20582 (
            .O(N__86699),
            .I(N__86658));
    Span4Mux_h I__20581 (
            .O(N__86694),
            .I(N__86658));
    Span4Mux_v I__20580 (
            .O(N__86689),
            .I(N__86655));
    Span4Mux_h I__20579 (
            .O(N__86686),
            .I(N__86652));
    Span4Mux_v I__20578 (
            .O(N__86683),
            .I(N__86649));
    Span4Mux_h I__20577 (
            .O(N__86680),
            .I(N__86644));
    Span4Mux_v I__20576 (
            .O(N__86673),
            .I(N__86644));
    Span4Mux_v I__20575 (
            .O(N__86668),
            .I(N__86641));
    Span4Mux_h I__20574 (
            .O(N__86663),
            .I(N__86638));
    Span4Mux_v I__20573 (
            .O(N__86658),
            .I(N__86635));
    Span4Mux_h I__20572 (
            .O(N__86655),
            .I(N__86630));
    Span4Mux_v I__20571 (
            .O(N__86652),
            .I(N__86630));
    Span4Mux_h I__20570 (
            .O(N__86649),
            .I(N__86625));
    Span4Mux_v I__20569 (
            .O(N__86644),
            .I(N__86625));
    Span4Mux_h I__20568 (
            .O(N__86641),
            .I(N__86620));
    Span4Mux_v I__20567 (
            .O(N__86638),
            .I(N__86620));
    Span4Mux_h I__20566 (
            .O(N__86635),
            .I(N__86617));
    Span4Mux_v I__20565 (
            .O(N__86630),
            .I(N__86614));
    Span4Mux_h I__20564 (
            .O(N__86625),
            .I(N__86611));
    Odrv4 I__20563 (
            .O(N__86620),
            .I(\pid_side.state_ns_0_0 ));
    Odrv4 I__20562 (
            .O(N__86617),
            .I(\pid_side.state_ns_0_0 ));
    Odrv4 I__20561 (
            .O(N__86614),
            .I(\pid_side.state_ns_0_0 ));
    Odrv4 I__20560 (
            .O(N__86611),
            .I(\pid_side.state_ns_0_0 ));
    InMux I__20559 (
            .O(N__86602),
            .I(N__86577));
    InMux I__20558 (
            .O(N__86601),
            .I(N__86572));
    InMux I__20557 (
            .O(N__86600),
            .I(N__86572));
    SRMux I__20556 (
            .O(N__86599),
            .I(N__86567));
    InMux I__20555 (
            .O(N__86598),
            .I(N__86567));
    SRMux I__20554 (
            .O(N__86597),
            .I(N__86562));
    InMux I__20553 (
            .O(N__86596),
            .I(N__86562));
    InMux I__20552 (
            .O(N__86595),
            .I(N__86559));
    InMux I__20551 (
            .O(N__86594),
            .I(N__86546));
    InMux I__20550 (
            .O(N__86593),
            .I(N__86546));
    InMux I__20549 (
            .O(N__86592),
            .I(N__86546));
    InMux I__20548 (
            .O(N__86591),
            .I(N__86546));
    InMux I__20547 (
            .O(N__86590),
            .I(N__86546));
    InMux I__20546 (
            .O(N__86589),
            .I(N__86546));
    InMux I__20545 (
            .O(N__86588),
            .I(N__86543));
    InMux I__20544 (
            .O(N__86587),
            .I(N__86540));
    InMux I__20543 (
            .O(N__86586),
            .I(N__86535));
    InMux I__20542 (
            .O(N__86585),
            .I(N__86535));
    InMux I__20541 (
            .O(N__86584),
            .I(N__86532));
    InMux I__20540 (
            .O(N__86583),
            .I(N__86529));
    InMux I__20539 (
            .O(N__86582),
            .I(N__86526));
    InMux I__20538 (
            .O(N__86581),
            .I(N__86523));
    InMux I__20537 (
            .O(N__86580),
            .I(N__86520));
    LocalMux I__20536 (
            .O(N__86577),
            .I(N__86349));
    LocalMux I__20535 (
            .O(N__86572),
            .I(N__86346));
    LocalMux I__20534 (
            .O(N__86567),
            .I(N__86343));
    LocalMux I__20533 (
            .O(N__86562),
            .I(N__86340));
    LocalMux I__20532 (
            .O(N__86559),
            .I(N__86337));
    LocalMux I__20531 (
            .O(N__86546),
            .I(N__86334));
    LocalMux I__20530 (
            .O(N__86543),
            .I(N__86331));
    LocalMux I__20529 (
            .O(N__86540),
            .I(N__86328));
    LocalMux I__20528 (
            .O(N__86535),
            .I(N__86325));
    LocalMux I__20527 (
            .O(N__86532),
            .I(N__86322));
    LocalMux I__20526 (
            .O(N__86529),
            .I(N__86319));
    LocalMux I__20525 (
            .O(N__86526),
            .I(N__86316));
    LocalMux I__20524 (
            .O(N__86523),
            .I(N__86313));
    LocalMux I__20523 (
            .O(N__86520),
            .I(N__86310));
    SRMux I__20522 (
            .O(N__86519),
            .I(N__85945));
    SRMux I__20521 (
            .O(N__86518),
            .I(N__85945));
    SRMux I__20520 (
            .O(N__86517),
            .I(N__85945));
    SRMux I__20519 (
            .O(N__86516),
            .I(N__85945));
    SRMux I__20518 (
            .O(N__86515),
            .I(N__85945));
    SRMux I__20517 (
            .O(N__86514),
            .I(N__85945));
    SRMux I__20516 (
            .O(N__86513),
            .I(N__85945));
    SRMux I__20515 (
            .O(N__86512),
            .I(N__85945));
    SRMux I__20514 (
            .O(N__86511),
            .I(N__85945));
    SRMux I__20513 (
            .O(N__86510),
            .I(N__85945));
    SRMux I__20512 (
            .O(N__86509),
            .I(N__85945));
    SRMux I__20511 (
            .O(N__86508),
            .I(N__85945));
    SRMux I__20510 (
            .O(N__86507),
            .I(N__85945));
    SRMux I__20509 (
            .O(N__86506),
            .I(N__85945));
    SRMux I__20508 (
            .O(N__86505),
            .I(N__85945));
    SRMux I__20507 (
            .O(N__86504),
            .I(N__85945));
    SRMux I__20506 (
            .O(N__86503),
            .I(N__85945));
    SRMux I__20505 (
            .O(N__86502),
            .I(N__85945));
    SRMux I__20504 (
            .O(N__86501),
            .I(N__85945));
    SRMux I__20503 (
            .O(N__86500),
            .I(N__85945));
    SRMux I__20502 (
            .O(N__86499),
            .I(N__85945));
    SRMux I__20501 (
            .O(N__86498),
            .I(N__85945));
    SRMux I__20500 (
            .O(N__86497),
            .I(N__85945));
    SRMux I__20499 (
            .O(N__86496),
            .I(N__85945));
    SRMux I__20498 (
            .O(N__86495),
            .I(N__85945));
    SRMux I__20497 (
            .O(N__86494),
            .I(N__85945));
    SRMux I__20496 (
            .O(N__86493),
            .I(N__85945));
    SRMux I__20495 (
            .O(N__86492),
            .I(N__85945));
    SRMux I__20494 (
            .O(N__86491),
            .I(N__85945));
    SRMux I__20493 (
            .O(N__86490),
            .I(N__85945));
    SRMux I__20492 (
            .O(N__86489),
            .I(N__85945));
    SRMux I__20491 (
            .O(N__86488),
            .I(N__85945));
    SRMux I__20490 (
            .O(N__86487),
            .I(N__85945));
    SRMux I__20489 (
            .O(N__86486),
            .I(N__85945));
    SRMux I__20488 (
            .O(N__86485),
            .I(N__85945));
    SRMux I__20487 (
            .O(N__86484),
            .I(N__85945));
    SRMux I__20486 (
            .O(N__86483),
            .I(N__85945));
    SRMux I__20485 (
            .O(N__86482),
            .I(N__85945));
    SRMux I__20484 (
            .O(N__86481),
            .I(N__85945));
    SRMux I__20483 (
            .O(N__86480),
            .I(N__85945));
    SRMux I__20482 (
            .O(N__86479),
            .I(N__85945));
    SRMux I__20481 (
            .O(N__86478),
            .I(N__85945));
    SRMux I__20480 (
            .O(N__86477),
            .I(N__85945));
    SRMux I__20479 (
            .O(N__86476),
            .I(N__85945));
    SRMux I__20478 (
            .O(N__86475),
            .I(N__85945));
    SRMux I__20477 (
            .O(N__86474),
            .I(N__85945));
    SRMux I__20476 (
            .O(N__86473),
            .I(N__85945));
    SRMux I__20475 (
            .O(N__86472),
            .I(N__85945));
    SRMux I__20474 (
            .O(N__86471),
            .I(N__85945));
    SRMux I__20473 (
            .O(N__86470),
            .I(N__85945));
    SRMux I__20472 (
            .O(N__86469),
            .I(N__85945));
    SRMux I__20471 (
            .O(N__86468),
            .I(N__85945));
    SRMux I__20470 (
            .O(N__86467),
            .I(N__85945));
    SRMux I__20469 (
            .O(N__86466),
            .I(N__85945));
    SRMux I__20468 (
            .O(N__86465),
            .I(N__85945));
    SRMux I__20467 (
            .O(N__86464),
            .I(N__85945));
    SRMux I__20466 (
            .O(N__86463),
            .I(N__85945));
    SRMux I__20465 (
            .O(N__86462),
            .I(N__85945));
    SRMux I__20464 (
            .O(N__86461),
            .I(N__85945));
    SRMux I__20463 (
            .O(N__86460),
            .I(N__85945));
    SRMux I__20462 (
            .O(N__86459),
            .I(N__85945));
    SRMux I__20461 (
            .O(N__86458),
            .I(N__85945));
    SRMux I__20460 (
            .O(N__86457),
            .I(N__85945));
    SRMux I__20459 (
            .O(N__86456),
            .I(N__85945));
    SRMux I__20458 (
            .O(N__86455),
            .I(N__85945));
    SRMux I__20457 (
            .O(N__86454),
            .I(N__85945));
    SRMux I__20456 (
            .O(N__86453),
            .I(N__85945));
    SRMux I__20455 (
            .O(N__86452),
            .I(N__85945));
    SRMux I__20454 (
            .O(N__86451),
            .I(N__85945));
    SRMux I__20453 (
            .O(N__86450),
            .I(N__85945));
    SRMux I__20452 (
            .O(N__86449),
            .I(N__85945));
    SRMux I__20451 (
            .O(N__86448),
            .I(N__85945));
    SRMux I__20450 (
            .O(N__86447),
            .I(N__85945));
    SRMux I__20449 (
            .O(N__86446),
            .I(N__85945));
    SRMux I__20448 (
            .O(N__86445),
            .I(N__85945));
    SRMux I__20447 (
            .O(N__86444),
            .I(N__85945));
    SRMux I__20446 (
            .O(N__86443),
            .I(N__85945));
    SRMux I__20445 (
            .O(N__86442),
            .I(N__85945));
    SRMux I__20444 (
            .O(N__86441),
            .I(N__85945));
    SRMux I__20443 (
            .O(N__86440),
            .I(N__85945));
    SRMux I__20442 (
            .O(N__86439),
            .I(N__85945));
    SRMux I__20441 (
            .O(N__86438),
            .I(N__85945));
    SRMux I__20440 (
            .O(N__86437),
            .I(N__85945));
    SRMux I__20439 (
            .O(N__86436),
            .I(N__85945));
    SRMux I__20438 (
            .O(N__86435),
            .I(N__85945));
    SRMux I__20437 (
            .O(N__86434),
            .I(N__85945));
    SRMux I__20436 (
            .O(N__86433),
            .I(N__85945));
    SRMux I__20435 (
            .O(N__86432),
            .I(N__85945));
    SRMux I__20434 (
            .O(N__86431),
            .I(N__85945));
    SRMux I__20433 (
            .O(N__86430),
            .I(N__85945));
    SRMux I__20432 (
            .O(N__86429),
            .I(N__85945));
    SRMux I__20431 (
            .O(N__86428),
            .I(N__85945));
    SRMux I__20430 (
            .O(N__86427),
            .I(N__85945));
    SRMux I__20429 (
            .O(N__86426),
            .I(N__85945));
    SRMux I__20428 (
            .O(N__86425),
            .I(N__85945));
    SRMux I__20427 (
            .O(N__86424),
            .I(N__85945));
    SRMux I__20426 (
            .O(N__86423),
            .I(N__85945));
    SRMux I__20425 (
            .O(N__86422),
            .I(N__85945));
    SRMux I__20424 (
            .O(N__86421),
            .I(N__85945));
    SRMux I__20423 (
            .O(N__86420),
            .I(N__85945));
    SRMux I__20422 (
            .O(N__86419),
            .I(N__85945));
    SRMux I__20421 (
            .O(N__86418),
            .I(N__85945));
    SRMux I__20420 (
            .O(N__86417),
            .I(N__85945));
    SRMux I__20419 (
            .O(N__86416),
            .I(N__85945));
    SRMux I__20418 (
            .O(N__86415),
            .I(N__85945));
    SRMux I__20417 (
            .O(N__86414),
            .I(N__85945));
    SRMux I__20416 (
            .O(N__86413),
            .I(N__85945));
    SRMux I__20415 (
            .O(N__86412),
            .I(N__85945));
    SRMux I__20414 (
            .O(N__86411),
            .I(N__85945));
    SRMux I__20413 (
            .O(N__86410),
            .I(N__85945));
    SRMux I__20412 (
            .O(N__86409),
            .I(N__85945));
    SRMux I__20411 (
            .O(N__86408),
            .I(N__85945));
    SRMux I__20410 (
            .O(N__86407),
            .I(N__85945));
    SRMux I__20409 (
            .O(N__86406),
            .I(N__85945));
    SRMux I__20408 (
            .O(N__86405),
            .I(N__85945));
    SRMux I__20407 (
            .O(N__86404),
            .I(N__85945));
    SRMux I__20406 (
            .O(N__86403),
            .I(N__85945));
    SRMux I__20405 (
            .O(N__86402),
            .I(N__85945));
    SRMux I__20404 (
            .O(N__86401),
            .I(N__85945));
    SRMux I__20403 (
            .O(N__86400),
            .I(N__85945));
    SRMux I__20402 (
            .O(N__86399),
            .I(N__85945));
    SRMux I__20401 (
            .O(N__86398),
            .I(N__85945));
    SRMux I__20400 (
            .O(N__86397),
            .I(N__85945));
    SRMux I__20399 (
            .O(N__86396),
            .I(N__85945));
    SRMux I__20398 (
            .O(N__86395),
            .I(N__85945));
    SRMux I__20397 (
            .O(N__86394),
            .I(N__85945));
    SRMux I__20396 (
            .O(N__86393),
            .I(N__85945));
    SRMux I__20395 (
            .O(N__86392),
            .I(N__85945));
    SRMux I__20394 (
            .O(N__86391),
            .I(N__85945));
    SRMux I__20393 (
            .O(N__86390),
            .I(N__85945));
    SRMux I__20392 (
            .O(N__86389),
            .I(N__85945));
    SRMux I__20391 (
            .O(N__86388),
            .I(N__85945));
    SRMux I__20390 (
            .O(N__86387),
            .I(N__85945));
    SRMux I__20389 (
            .O(N__86386),
            .I(N__85945));
    SRMux I__20388 (
            .O(N__86385),
            .I(N__85945));
    SRMux I__20387 (
            .O(N__86384),
            .I(N__85945));
    SRMux I__20386 (
            .O(N__86383),
            .I(N__85945));
    SRMux I__20385 (
            .O(N__86382),
            .I(N__85945));
    SRMux I__20384 (
            .O(N__86381),
            .I(N__85945));
    SRMux I__20383 (
            .O(N__86380),
            .I(N__85945));
    SRMux I__20382 (
            .O(N__86379),
            .I(N__85945));
    SRMux I__20381 (
            .O(N__86378),
            .I(N__85945));
    SRMux I__20380 (
            .O(N__86377),
            .I(N__85945));
    SRMux I__20379 (
            .O(N__86376),
            .I(N__85945));
    SRMux I__20378 (
            .O(N__86375),
            .I(N__85945));
    SRMux I__20377 (
            .O(N__86374),
            .I(N__85945));
    SRMux I__20376 (
            .O(N__86373),
            .I(N__85945));
    SRMux I__20375 (
            .O(N__86372),
            .I(N__85945));
    SRMux I__20374 (
            .O(N__86371),
            .I(N__85945));
    SRMux I__20373 (
            .O(N__86370),
            .I(N__85945));
    SRMux I__20372 (
            .O(N__86369),
            .I(N__85945));
    SRMux I__20371 (
            .O(N__86368),
            .I(N__85945));
    SRMux I__20370 (
            .O(N__86367),
            .I(N__85945));
    SRMux I__20369 (
            .O(N__86366),
            .I(N__85945));
    SRMux I__20368 (
            .O(N__86365),
            .I(N__85945));
    SRMux I__20367 (
            .O(N__86364),
            .I(N__85945));
    SRMux I__20366 (
            .O(N__86363),
            .I(N__85945));
    SRMux I__20365 (
            .O(N__86362),
            .I(N__85945));
    SRMux I__20364 (
            .O(N__86361),
            .I(N__85945));
    SRMux I__20363 (
            .O(N__86360),
            .I(N__85945));
    SRMux I__20362 (
            .O(N__86359),
            .I(N__85945));
    SRMux I__20361 (
            .O(N__86358),
            .I(N__85945));
    SRMux I__20360 (
            .O(N__86357),
            .I(N__85945));
    SRMux I__20359 (
            .O(N__86356),
            .I(N__85945));
    SRMux I__20358 (
            .O(N__86355),
            .I(N__85945));
    SRMux I__20357 (
            .O(N__86354),
            .I(N__85945));
    SRMux I__20356 (
            .O(N__86353),
            .I(N__85945));
    SRMux I__20355 (
            .O(N__86352),
            .I(N__85945));
    Glb2LocalMux I__20354 (
            .O(N__86349),
            .I(N__85945));
    Glb2LocalMux I__20353 (
            .O(N__86346),
            .I(N__85945));
    Glb2LocalMux I__20352 (
            .O(N__86343),
            .I(N__85945));
    Glb2LocalMux I__20351 (
            .O(N__86340),
            .I(N__85945));
    Glb2LocalMux I__20350 (
            .O(N__86337),
            .I(N__85945));
    Glb2LocalMux I__20349 (
            .O(N__86334),
            .I(N__85945));
    Glb2LocalMux I__20348 (
            .O(N__86331),
            .I(N__85945));
    Glb2LocalMux I__20347 (
            .O(N__86328),
            .I(N__85945));
    Glb2LocalMux I__20346 (
            .O(N__86325),
            .I(N__85945));
    Glb2LocalMux I__20345 (
            .O(N__86322),
            .I(N__85945));
    Glb2LocalMux I__20344 (
            .O(N__86319),
            .I(N__85945));
    Glb2LocalMux I__20343 (
            .O(N__86316),
            .I(N__85945));
    Glb2LocalMux I__20342 (
            .O(N__86313),
            .I(N__85945));
    Glb2LocalMux I__20341 (
            .O(N__86310),
            .I(N__85945));
    GlobalMux I__20340 (
            .O(N__85945),
            .I(N__85942));
    gio2CtrlBuf I__20339 (
            .O(N__85942),
            .I(reset_module_System_reset_iso_g));
    InMux I__20338 (
            .O(N__85939),
            .I(N__85931));
    InMux I__20337 (
            .O(N__85938),
            .I(N__85920));
    InMux I__20336 (
            .O(N__85937),
            .I(N__85916));
    InMux I__20335 (
            .O(N__85936),
            .I(N__85913));
    InMux I__20334 (
            .O(N__85935),
            .I(N__85904));
    InMux I__20333 (
            .O(N__85934),
            .I(N__85904));
    LocalMux I__20332 (
            .O(N__85931),
            .I(N__85901));
    InMux I__20331 (
            .O(N__85930),
            .I(N__85892));
    InMux I__20330 (
            .O(N__85929),
            .I(N__85892));
    InMux I__20329 (
            .O(N__85928),
            .I(N__85892));
    InMux I__20328 (
            .O(N__85927),
            .I(N__85892));
    InMux I__20327 (
            .O(N__85926),
            .I(N__85889));
    InMux I__20326 (
            .O(N__85925),
            .I(N__85886));
    InMux I__20325 (
            .O(N__85924),
            .I(N__85883));
    InMux I__20324 (
            .O(N__85923),
            .I(N__85880));
    LocalMux I__20323 (
            .O(N__85920),
            .I(N__85877));
    InMux I__20322 (
            .O(N__85919),
            .I(N__85874));
    LocalMux I__20321 (
            .O(N__85916),
            .I(N__85871));
    LocalMux I__20320 (
            .O(N__85913),
            .I(N__85868));
    InMux I__20319 (
            .O(N__85912),
            .I(N__85861));
    InMux I__20318 (
            .O(N__85911),
            .I(N__85861));
    InMux I__20317 (
            .O(N__85910),
            .I(N__85861));
    InMux I__20316 (
            .O(N__85909),
            .I(N__85857));
    LocalMux I__20315 (
            .O(N__85904),
            .I(N__85850));
    Span4Mux_h I__20314 (
            .O(N__85901),
            .I(N__85850));
    LocalMux I__20313 (
            .O(N__85892),
            .I(N__85850));
    LocalMux I__20312 (
            .O(N__85889),
            .I(N__85846));
    LocalMux I__20311 (
            .O(N__85886),
            .I(N__85843));
    LocalMux I__20310 (
            .O(N__85883),
            .I(N__85832));
    LocalMux I__20309 (
            .O(N__85880),
            .I(N__85832));
    Span4Mux_v I__20308 (
            .O(N__85877),
            .I(N__85832));
    LocalMux I__20307 (
            .O(N__85874),
            .I(N__85832));
    Span4Mux_v I__20306 (
            .O(N__85871),
            .I(N__85825));
    Span4Mux_v I__20305 (
            .O(N__85868),
            .I(N__85825));
    LocalMux I__20304 (
            .O(N__85861),
            .I(N__85825));
    InMux I__20303 (
            .O(N__85860),
            .I(N__85822));
    LocalMux I__20302 (
            .O(N__85857),
            .I(N__85817));
    Span4Mux_h I__20301 (
            .O(N__85850),
            .I(N__85817));
    InMux I__20300 (
            .O(N__85849),
            .I(N__85814));
    Span4Mux_v I__20299 (
            .O(N__85846),
            .I(N__85809));
    Span4Mux_h I__20298 (
            .O(N__85843),
            .I(N__85809));
    InMux I__20297 (
            .O(N__85842),
            .I(N__85804));
    InMux I__20296 (
            .O(N__85841),
            .I(N__85804));
    Span4Mux_h I__20295 (
            .O(N__85832),
            .I(N__85799));
    Span4Mux_h I__20294 (
            .O(N__85825),
            .I(N__85799));
    LocalMux I__20293 (
            .O(N__85822),
            .I(N__85794));
    Span4Mux_v I__20292 (
            .O(N__85817),
            .I(N__85794));
    LocalMux I__20291 (
            .O(N__85814),
            .I(\pid_side.error_15 ));
    Odrv4 I__20290 (
            .O(N__85809),
            .I(\pid_side.error_15 ));
    LocalMux I__20289 (
            .O(N__85804),
            .I(\pid_side.error_15 ));
    Odrv4 I__20288 (
            .O(N__85799),
            .I(\pid_side.error_15 ));
    Odrv4 I__20287 (
            .O(N__85794),
            .I(\pid_side.error_15 ));
    InMux I__20286 (
            .O(N__85783),
            .I(N__85780));
    LocalMux I__20285 (
            .O(N__85780),
            .I(\pid_side.N_622 ));
    InMux I__20284 (
            .O(N__85777),
            .I(N__85772));
    InMux I__20283 (
            .O(N__85776),
            .I(N__85765));
    CascadeMux I__20282 (
            .O(N__85775),
            .I(N__85760));
    LocalMux I__20281 (
            .O(N__85772),
            .I(N__85757));
    InMux I__20280 (
            .O(N__85771),
            .I(N__85754));
    CascadeMux I__20279 (
            .O(N__85770),
            .I(N__85751));
    CascadeMux I__20278 (
            .O(N__85769),
            .I(N__85743));
    CascadeMux I__20277 (
            .O(N__85768),
            .I(N__85740));
    LocalMux I__20276 (
            .O(N__85765),
            .I(N__85734));
    InMux I__20275 (
            .O(N__85764),
            .I(N__85728));
    InMux I__20274 (
            .O(N__85763),
            .I(N__85728));
    InMux I__20273 (
            .O(N__85760),
            .I(N__85725));
    Span4Mux_v I__20272 (
            .O(N__85757),
            .I(N__85720));
    LocalMux I__20271 (
            .O(N__85754),
            .I(N__85720));
    InMux I__20270 (
            .O(N__85751),
            .I(N__85717));
    InMux I__20269 (
            .O(N__85750),
            .I(N__85713));
    InMux I__20268 (
            .O(N__85749),
            .I(N__85710));
    InMux I__20267 (
            .O(N__85748),
            .I(N__85707));
    InMux I__20266 (
            .O(N__85747),
            .I(N__85704));
    InMux I__20265 (
            .O(N__85746),
            .I(N__85701));
    InMux I__20264 (
            .O(N__85743),
            .I(N__85698));
    InMux I__20263 (
            .O(N__85740),
            .I(N__85695));
    InMux I__20262 (
            .O(N__85739),
            .I(N__85692));
    InMux I__20261 (
            .O(N__85738),
            .I(N__85687));
    InMux I__20260 (
            .O(N__85737),
            .I(N__85687));
    Span4Mux_v I__20259 (
            .O(N__85734),
            .I(N__85684));
    InMux I__20258 (
            .O(N__85733),
            .I(N__85681));
    LocalMux I__20257 (
            .O(N__85728),
            .I(N__85678));
    LocalMux I__20256 (
            .O(N__85725),
            .I(N__85675));
    Span4Mux_h I__20255 (
            .O(N__85720),
            .I(N__85670));
    LocalMux I__20254 (
            .O(N__85717),
            .I(N__85670));
    InMux I__20253 (
            .O(N__85716),
            .I(N__85667));
    LocalMux I__20252 (
            .O(N__85713),
            .I(N__85662));
    LocalMux I__20251 (
            .O(N__85710),
            .I(N__85662));
    LocalMux I__20250 (
            .O(N__85707),
            .I(N__85655));
    LocalMux I__20249 (
            .O(N__85704),
            .I(N__85655));
    LocalMux I__20248 (
            .O(N__85701),
            .I(N__85655));
    LocalMux I__20247 (
            .O(N__85698),
            .I(N__85648));
    LocalMux I__20246 (
            .O(N__85695),
            .I(N__85648));
    LocalMux I__20245 (
            .O(N__85692),
            .I(N__85648));
    LocalMux I__20244 (
            .O(N__85687),
            .I(N__85645));
    Sp12to4 I__20243 (
            .O(N__85684),
            .I(N__85640));
    LocalMux I__20242 (
            .O(N__85681),
            .I(N__85640));
    Span4Mux_h I__20241 (
            .O(N__85678),
            .I(N__85633));
    Span4Mux_v I__20240 (
            .O(N__85675),
            .I(N__85633));
    Span4Mux_h I__20239 (
            .O(N__85670),
            .I(N__85633));
    LocalMux I__20238 (
            .O(N__85667),
            .I(N__85628));
    Span4Mux_v I__20237 (
            .O(N__85662),
            .I(N__85628));
    Span4Mux_h I__20236 (
            .O(N__85655),
            .I(N__85625));
    Span4Mux_v I__20235 (
            .O(N__85648),
            .I(N__85620));
    Span4Mux_v I__20234 (
            .O(N__85645),
            .I(N__85620));
    Span12Mux_h I__20233 (
            .O(N__85640),
            .I(N__85617));
    Span4Mux_v I__20232 (
            .O(N__85633),
            .I(N__85614));
    Span4Mux_h I__20231 (
            .O(N__85628),
            .I(N__85609));
    Span4Mux_h I__20230 (
            .O(N__85625),
            .I(N__85609));
    Odrv4 I__20229 (
            .O(N__85620),
            .I(pid_side_N_493));
    Odrv12 I__20228 (
            .O(N__85617),
            .I(pid_side_N_493));
    Odrv4 I__20227 (
            .O(N__85614),
            .I(pid_side_N_493));
    Odrv4 I__20226 (
            .O(N__85609),
            .I(pid_side_N_493));
    InMux I__20225 (
            .O(N__85600),
            .I(N__85596));
    InMux I__20224 (
            .O(N__85599),
            .I(N__85593));
    LocalMux I__20223 (
            .O(N__85596),
            .I(N__85589));
    LocalMux I__20222 (
            .O(N__85593),
            .I(N__85586));
    InMux I__20221 (
            .O(N__85592),
            .I(N__85583));
    Span4Mux_h I__20220 (
            .O(N__85589),
            .I(N__85580));
    Odrv4 I__20219 (
            .O(N__85586),
            .I(\pid_side.N_226 ));
    LocalMux I__20218 (
            .O(N__85583),
            .I(\pid_side.N_226 ));
    Odrv4 I__20217 (
            .O(N__85580),
            .I(\pid_side.N_226 ));
    CascadeMux I__20216 (
            .O(N__85573),
            .I(N__85570));
    InMux I__20215 (
            .O(N__85570),
            .I(N__85567));
    LocalMux I__20214 (
            .O(N__85567),
            .I(N__85563));
    CascadeMux I__20213 (
            .O(N__85566),
            .I(N__85560));
    Span4Mux_h I__20212 (
            .O(N__85563),
            .I(N__85557));
    InMux I__20211 (
            .O(N__85560),
            .I(N__85554));
    Odrv4 I__20210 (
            .O(N__85557),
            .I(pid_side_m22_2_03_0_a2_0));
    LocalMux I__20209 (
            .O(N__85554),
            .I(pid_side_m22_2_03_0_a2_0));
    InMux I__20208 (
            .O(N__85549),
            .I(N__85546));
    LocalMux I__20207 (
            .O(N__85546),
            .I(\pid_side.N_254 ));
    InMux I__20206 (
            .O(N__85543),
            .I(N__85540));
    LocalMux I__20205 (
            .O(N__85540),
            .I(N__85537));
    Odrv12 I__20204 (
            .O(N__85537),
            .I(\pid_side.m22_2_03_0_0 ));
    InMux I__20203 (
            .O(N__85534),
            .I(N__85531));
    LocalMux I__20202 (
            .O(N__85531),
            .I(N__85523));
    InMux I__20201 (
            .O(N__85530),
            .I(N__85520));
    InMux I__20200 (
            .O(N__85529),
            .I(N__85517));
    InMux I__20199 (
            .O(N__85528),
            .I(N__85514));
    InMux I__20198 (
            .O(N__85527),
            .I(N__85510));
    InMux I__20197 (
            .O(N__85526),
            .I(N__85506));
    Span4Mux_h I__20196 (
            .O(N__85523),
            .I(N__85499));
    LocalMux I__20195 (
            .O(N__85520),
            .I(N__85499));
    LocalMux I__20194 (
            .O(N__85517),
            .I(N__85499));
    LocalMux I__20193 (
            .O(N__85514),
            .I(N__85496));
    InMux I__20192 (
            .O(N__85513),
            .I(N__85493));
    LocalMux I__20191 (
            .O(N__85510),
            .I(N__85490));
    InMux I__20190 (
            .O(N__85509),
            .I(N__85486));
    LocalMux I__20189 (
            .O(N__85506),
            .I(N__85482));
    Span4Mux_v I__20188 (
            .O(N__85499),
            .I(N__85477));
    Span4Mux_v I__20187 (
            .O(N__85496),
            .I(N__85472));
    LocalMux I__20186 (
            .O(N__85493),
            .I(N__85472));
    Span4Mux_h I__20185 (
            .O(N__85490),
            .I(N__85469));
    InMux I__20184 (
            .O(N__85489),
            .I(N__85465));
    LocalMux I__20183 (
            .O(N__85486),
            .I(N__85461));
    InMux I__20182 (
            .O(N__85485),
            .I(N__85458));
    Span4Mux_h I__20181 (
            .O(N__85482),
            .I(N__85454));
    InMux I__20180 (
            .O(N__85481),
            .I(N__85449));
    InMux I__20179 (
            .O(N__85480),
            .I(N__85449));
    Span4Mux_h I__20178 (
            .O(N__85477),
            .I(N__85446));
    Span4Mux_h I__20177 (
            .O(N__85472),
            .I(N__85442));
    Span4Mux_v I__20176 (
            .O(N__85469),
            .I(N__85439));
    InMux I__20175 (
            .O(N__85468),
            .I(N__85436));
    LocalMux I__20174 (
            .O(N__85465),
            .I(N__85433));
    InMux I__20173 (
            .O(N__85464),
            .I(N__85430));
    Span4Mux_v I__20172 (
            .O(N__85461),
            .I(N__85427));
    LocalMux I__20171 (
            .O(N__85458),
            .I(N__85424));
    InMux I__20170 (
            .O(N__85457),
            .I(N__85421));
    Span4Mux_v I__20169 (
            .O(N__85454),
            .I(N__85418));
    LocalMux I__20168 (
            .O(N__85449),
            .I(N__85415));
    Sp12to4 I__20167 (
            .O(N__85446),
            .I(N__85411));
    InMux I__20166 (
            .O(N__85445),
            .I(N__85408));
    Span4Mux_h I__20165 (
            .O(N__85442),
            .I(N__85403));
    Span4Mux_h I__20164 (
            .O(N__85439),
            .I(N__85403));
    LocalMux I__20163 (
            .O(N__85436),
            .I(N__85396));
    Span12Mux_s9_h I__20162 (
            .O(N__85433),
            .I(N__85396));
    LocalMux I__20161 (
            .O(N__85430),
            .I(N__85396));
    Span4Mux_v I__20160 (
            .O(N__85427),
            .I(N__85389));
    Span4Mux_h I__20159 (
            .O(N__85424),
            .I(N__85389));
    LocalMux I__20158 (
            .O(N__85421),
            .I(N__85389));
    Span4Mux_v I__20157 (
            .O(N__85418),
            .I(N__85384));
    Span4Mux_h I__20156 (
            .O(N__85415),
            .I(N__85384));
    InMux I__20155 (
            .O(N__85414),
            .I(N__85381));
    Odrv12 I__20154 (
            .O(N__85411),
            .I(uart_pc_data_1));
    LocalMux I__20153 (
            .O(N__85408),
            .I(uart_pc_data_1));
    Odrv4 I__20152 (
            .O(N__85403),
            .I(uart_pc_data_1));
    Odrv12 I__20151 (
            .O(N__85396),
            .I(uart_pc_data_1));
    Odrv4 I__20150 (
            .O(N__85389),
            .I(uart_pc_data_1));
    Odrv4 I__20149 (
            .O(N__85384),
            .I(uart_pc_data_1));
    LocalMux I__20148 (
            .O(N__85381),
            .I(uart_pc_data_1));
    CascadeMux I__20147 (
            .O(N__85366),
            .I(N__85363));
    InMux I__20146 (
            .O(N__85363),
            .I(N__85360));
    LocalMux I__20145 (
            .O(N__85360),
            .I(N__85357));
    Odrv12 I__20144 (
            .O(N__85357),
            .I(side_command_1));
    CascadeMux I__20143 (
            .O(N__85354),
            .I(N__85351));
    InMux I__20142 (
            .O(N__85351),
            .I(N__85348));
    LocalMux I__20141 (
            .O(N__85348),
            .I(N__85345));
    Span4Mux_h I__20140 (
            .O(N__85345),
            .I(N__85342));
    Odrv4 I__20139 (
            .O(N__85342),
            .I(side_command_2));
    CascadeMux I__20138 (
            .O(N__85339),
            .I(N__85336));
    InMux I__20137 (
            .O(N__85336),
            .I(N__85333));
    LocalMux I__20136 (
            .O(N__85333),
            .I(N__85330));
    Odrv12 I__20135 (
            .O(N__85330),
            .I(side_command_3));
    CascadeMux I__20134 (
            .O(N__85327),
            .I(N__85324));
    InMux I__20133 (
            .O(N__85324),
            .I(N__85321));
    LocalMux I__20132 (
            .O(N__85321),
            .I(N__85318));
    Span4Mux_v I__20131 (
            .O(N__85318),
            .I(N__85315));
    Odrv4 I__20130 (
            .O(N__85315),
            .I(side_command_4));
    CascadeMux I__20129 (
            .O(N__85312),
            .I(N__85309));
    InMux I__20128 (
            .O(N__85309),
            .I(N__85306));
    LocalMux I__20127 (
            .O(N__85306),
            .I(N__85303));
    Span4Mux_v I__20126 (
            .O(N__85303),
            .I(N__85300));
    Sp12to4 I__20125 (
            .O(N__85300),
            .I(N__85297));
    Odrv12 I__20124 (
            .O(N__85297),
            .I(side_command_5));
    CascadeMux I__20123 (
            .O(N__85294),
            .I(N__85291));
    InMux I__20122 (
            .O(N__85291),
            .I(N__85288));
    LocalMux I__20121 (
            .O(N__85288),
            .I(N__85285));
    Span4Mux_h I__20120 (
            .O(N__85285),
            .I(N__85282));
    Odrv4 I__20119 (
            .O(N__85282),
            .I(side_command_6));
    CascadeMux I__20118 (
            .O(N__85279),
            .I(N__85276));
    InMux I__20117 (
            .O(N__85276),
            .I(N__85270));
    InMux I__20116 (
            .O(N__85275),
            .I(N__85270));
    LocalMux I__20115 (
            .O(N__85270),
            .I(N__85267));
    Odrv12 I__20114 (
            .O(N__85267),
            .I(side_command_7));
    CEMux I__20113 (
            .O(N__85264),
            .I(N__85261));
    LocalMux I__20112 (
            .O(N__85261),
            .I(N__85258));
    Span12Mux_s4_h I__20111 (
            .O(N__85258),
            .I(N__85255));
    Odrv12 I__20110 (
            .O(N__85255),
            .I(\Commands_frame_decoder.source_CH2data_1_sqmuxa_0 ));
    CascadeMux I__20109 (
            .O(N__85252),
            .I(N__85247));
    InMux I__20108 (
            .O(N__85251),
            .I(N__85243));
    InMux I__20107 (
            .O(N__85250),
            .I(N__85240));
    InMux I__20106 (
            .O(N__85247),
            .I(N__85237));
    CascadeMux I__20105 (
            .O(N__85246),
            .I(N__85234));
    LocalMux I__20104 (
            .O(N__85243),
            .I(N__85229));
    LocalMux I__20103 (
            .O(N__85240),
            .I(N__85226));
    LocalMux I__20102 (
            .O(N__85237),
            .I(N__85222));
    InMux I__20101 (
            .O(N__85234),
            .I(N__85217));
    InMux I__20100 (
            .O(N__85233),
            .I(N__85217));
    InMux I__20099 (
            .O(N__85232),
            .I(N__85214));
    Span4Mux_s2_h I__20098 (
            .O(N__85229),
            .I(N__85211));
    Span4Mux_s0_h I__20097 (
            .O(N__85226),
            .I(N__85208));
    InMux I__20096 (
            .O(N__85225),
            .I(N__85205));
    Span4Mux_v I__20095 (
            .O(N__85222),
            .I(N__85200));
    LocalMux I__20094 (
            .O(N__85217),
            .I(N__85200));
    LocalMux I__20093 (
            .O(N__85214),
            .I(N__85195));
    Span4Mux_v I__20092 (
            .O(N__85211),
            .I(N__85195));
    Span4Mux_h I__20091 (
            .O(N__85208),
            .I(N__85190));
    LocalMux I__20090 (
            .O(N__85205),
            .I(N__85190));
    Span4Mux_h I__20089 (
            .O(N__85200),
            .I(N__85187));
    Odrv4 I__20088 (
            .O(N__85195),
            .I(\pid_side.error_8 ));
    Odrv4 I__20087 (
            .O(N__85190),
            .I(\pid_side.error_8 ));
    Odrv4 I__20086 (
            .O(N__85187),
            .I(\pid_side.error_8 ));
    CascadeMux I__20085 (
            .O(N__85180),
            .I(N__85175));
    CascadeMux I__20084 (
            .O(N__85179),
            .I(N__85172));
    CascadeMux I__20083 (
            .O(N__85178),
            .I(N__85169));
    InMux I__20082 (
            .O(N__85175),
            .I(N__85166));
    InMux I__20081 (
            .O(N__85172),
            .I(N__85162));
    InMux I__20080 (
            .O(N__85169),
            .I(N__85153));
    LocalMux I__20079 (
            .O(N__85166),
            .I(N__85150));
    InMux I__20078 (
            .O(N__85165),
            .I(N__85147));
    LocalMux I__20077 (
            .O(N__85162),
            .I(N__85144));
    InMux I__20076 (
            .O(N__85161),
            .I(N__85141));
    CascadeMux I__20075 (
            .O(N__85160),
            .I(N__85138));
    CascadeMux I__20074 (
            .O(N__85159),
            .I(N__85134));
    InMux I__20073 (
            .O(N__85158),
            .I(N__85129));
    InMux I__20072 (
            .O(N__85157),
            .I(N__85124));
    CascadeMux I__20071 (
            .O(N__85156),
            .I(N__85121));
    LocalMux I__20070 (
            .O(N__85153),
            .I(N__85118));
    Span4Mux_h I__20069 (
            .O(N__85150),
            .I(N__85111));
    LocalMux I__20068 (
            .O(N__85147),
            .I(N__85104));
    Span4Mux_v I__20067 (
            .O(N__85144),
            .I(N__85104));
    LocalMux I__20066 (
            .O(N__85141),
            .I(N__85104));
    InMux I__20065 (
            .O(N__85138),
            .I(N__85101));
    InMux I__20064 (
            .O(N__85137),
            .I(N__85096));
    InMux I__20063 (
            .O(N__85134),
            .I(N__85096));
    InMux I__20062 (
            .O(N__85133),
            .I(N__85091));
    InMux I__20061 (
            .O(N__85132),
            .I(N__85091));
    LocalMux I__20060 (
            .O(N__85129),
            .I(N__85088));
    InMux I__20059 (
            .O(N__85128),
            .I(N__85085));
    InMux I__20058 (
            .O(N__85127),
            .I(N__85081));
    LocalMux I__20057 (
            .O(N__85124),
            .I(N__85078));
    InMux I__20056 (
            .O(N__85121),
            .I(N__85073));
    Span4Mux_h I__20055 (
            .O(N__85118),
            .I(N__85070));
    InMux I__20054 (
            .O(N__85117),
            .I(N__85062));
    InMux I__20053 (
            .O(N__85116),
            .I(N__85055));
    InMux I__20052 (
            .O(N__85115),
            .I(N__85055));
    InMux I__20051 (
            .O(N__85114),
            .I(N__85055));
    Span4Mux_v I__20050 (
            .O(N__85111),
            .I(N__85045));
    Span4Mux_h I__20049 (
            .O(N__85104),
            .I(N__85045));
    LocalMux I__20048 (
            .O(N__85101),
            .I(N__85045));
    LocalMux I__20047 (
            .O(N__85096),
            .I(N__85045));
    LocalMux I__20046 (
            .O(N__85091),
            .I(N__85038));
    Span4Mux_v I__20045 (
            .O(N__85088),
            .I(N__85038));
    LocalMux I__20044 (
            .O(N__85085),
            .I(N__85038));
    InMux I__20043 (
            .O(N__85084),
            .I(N__85035));
    LocalMux I__20042 (
            .O(N__85081),
            .I(N__85029));
    Span4Mux_h I__20041 (
            .O(N__85078),
            .I(N__85029));
    CascadeMux I__20040 (
            .O(N__85077),
            .I(N__85026));
    CascadeMux I__20039 (
            .O(N__85076),
            .I(N__85022));
    LocalMux I__20038 (
            .O(N__85073),
            .I(N__85019));
    Span4Mux_h I__20037 (
            .O(N__85070),
            .I(N__85016));
    InMux I__20036 (
            .O(N__85069),
            .I(N__85013));
    InMux I__20035 (
            .O(N__85068),
            .I(N__85006));
    InMux I__20034 (
            .O(N__85067),
            .I(N__85006));
    InMux I__20033 (
            .O(N__85066),
            .I(N__85006));
    CascadeMux I__20032 (
            .O(N__85065),
            .I(N__85002));
    LocalMux I__20031 (
            .O(N__85062),
            .I(N__84997));
    LocalMux I__20030 (
            .O(N__85055),
            .I(N__84997));
    InMux I__20029 (
            .O(N__85054),
            .I(N__84994));
    Span4Mux_v I__20028 (
            .O(N__85045),
            .I(N__84989));
    Span4Mux_h I__20027 (
            .O(N__85038),
            .I(N__84989));
    LocalMux I__20026 (
            .O(N__85035),
            .I(N__84986));
    InMux I__20025 (
            .O(N__85034),
            .I(N__84983));
    Span4Mux_v I__20024 (
            .O(N__85029),
            .I(N__84980));
    InMux I__20023 (
            .O(N__85026),
            .I(N__84973));
    InMux I__20022 (
            .O(N__85025),
            .I(N__84973));
    InMux I__20021 (
            .O(N__85022),
            .I(N__84973));
    Span4Mux_v I__20020 (
            .O(N__85019),
            .I(N__84964));
    Span4Mux_s3_h I__20019 (
            .O(N__85016),
            .I(N__84964));
    LocalMux I__20018 (
            .O(N__85013),
            .I(N__84964));
    LocalMux I__20017 (
            .O(N__85006),
            .I(N__84964));
    InMux I__20016 (
            .O(N__85005),
            .I(N__84959));
    InMux I__20015 (
            .O(N__85002),
            .I(N__84959));
    Span4Mux_v I__20014 (
            .O(N__84997),
            .I(N__84954));
    LocalMux I__20013 (
            .O(N__84994),
            .I(N__84954));
    Span4Mux_h I__20012 (
            .O(N__84989),
            .I(N__84951));
    Odrv12 I__20011 (
            .O(N__84986),
            .I(xy_ki_3_rep2));
    LocalMux I__20010 (
            .O(N__84983),
            .I(xy_ki_3_rep2));
    Odrv4 I__20009 (
            .O(N__84980),
            .I(xy_ki_3_rep2));
    LocalMux I__20008 (
            .O(N__84973),
            .I(xy_ki_3_rep2));
    Odrv4 I__20007 (
            .O(N__84964),
            .I(xy_ki_3_rep2));
    LocalMux I__20006 (
            .O(N__84959),
            .I(xy_ki_3_rep2));
    Odrv4 I__20005 (
            .O(N__84954),
            .I(xy_ki_3_rep2));
    Odrv4 I__20004 (
            .O(N__84951),
            .I(xy_ki_3_rep2));
    InMux I__20003 (
            .O(N__84934),
            .I(N__84929));
    InMux I__20002 (
            .O(N__84933),
            .I(N__84926));
    InMux I__20001 (
            .O(N__84932),
            .I(N__84923));
    LocalMux I__20000 (
            .O(N__84929),
            .I(N__84919));
    LocalMux I__19999 (
            .O(N__84926),
            .I(N__84916));
    LocalMux I__19998 (
            .O(N__84923),
            .I(N__84912));
    InMux I__19997 (
            .O(N__84922),
            .I(N__84908));
    Span4Mux_h I__19996 (
            .O(N__84919),
            .I(N__84905));
    Span4Mux_v I__19995 (
            .O(N__84916),
            .I(N__84902));
    InMux I__19994 (
            .O(N__84915),
            .I(N__84899));
    Span4Mux_s1_h I__19993 (
            .O(N__84912),
            .I(N__84893));
    InMux I__19992 (
            .O(N__84911),
            .I(N__84890));
    LocalMux I__19991 (
            .O(N__84908),
            .I(N__84887));
    Span4Mux_v I__19990 (
            .O(N__84905),
            .I(N__84884));
    Span4Mux_h I__19989 (
            .O(N__84902),
            .I(N__84879));
    LocalMux I__19988 (
            .O(N__84899),
            .I(N__84879));
    InMux I__19987 (
            .O(N__84898),
            .I(N__84872));
    InMux I__19986 (
            .O(N__84897),
            .I(N__84872));
    InMux I__19985 (
            .O(N__84896),
            .I(N__84872));
    Span4Mux_v I__19984 (
            .O(N__84893),
            .I(N__84867));
    LocalMux I__19983 (
            .O(N__84890),
            .I(N__84867));
    Span4Mux_h I__19982 (
            .O(N__84887),
            .I(N__84864));
    Odrv4 I__19981 (
            .O(N__84884),
            .I(\pid_side.error_12 ));
    Odrv4 I__19980 (
            .O(N__84879),
            .I(\pid_side.error_12 ));
    LocalMux I__19979 (
            .O(N__84872),
            .I(\pid_side.error_12 ));
    Odrv4 I__19978 (
            .O(N__84867),
            .I(\pid_side.error_12 ));
    Odrv4 I__19977 (
            .O(N__84864),
            .I(\pid_side.error_12 ));
    CascadeMux I__19976 (
            .O(N__84853),
            .I(\pid_side.N_226_cascade_ ));
    CascadeMux I__19975 (
            .O(N__84850),
            .I(N__84847));
    InMux I__19974 (
            .O(N__84847),
            .I(N__84844));
    LocalMux I__19973 (
            .O(N__84844),
            .I(N__84841));
    Odrv4 I__19972 (
            .O(N__84841),
            .I(\pid_side.m58_0_a2_1_sxZ0 ));
    InMux I__19971 (
            .O(N__84838),
            .I(N__84828));
    CascadeMux I__19970 (
            .O(N__84837),
            .I(N__84823));
    InMux I__19969 (
            .O(N__84836),
            .I(N__84820));
    InMux I__19968 (
            .O(N__84835),
            .I(N__84817));
    InMux I__19967 (
            .O(N__84834),
            .I(N__84812));
    CascadeMux I__19966 (
            .O(N__84833),
            .I(N__84809));
    InMux I__19965 (
            .O(N__84832),
            .I(N__84806));
    InMux I__19964 (
            .O(N__84831),
            .I(N__84803));
    LocalMux I__19963 (
            .O(N__84828),
            .I(N__84800));
    InMux I__19962 (
            .O(N__84827),
            .I(N__84797));
    InMux I__19961 (
            .O(N__84826),
            .I(N__84794));
    InMux I__19960 (
            .O(N__84823),
            .I(N__84791));
    LocalMux I__19959 (
            .O(N__84820),
            .I(N__84788));
    LocalMux I__19958 (
            .O(N__84817),
            .I(N__84782));
    InMux I__19957 (
            .O(N__84816),
            .I(N__84777));
    InMux I__19956 (
            .O(N__84815),
            .I(N__84777));
    LocalMux I__19955 (
            .O(N__84812),
            .I(N__84774));
    InMux I__19954 (
            .O(N__84809),
            .I(N__84771));
    LocalMux I__19953 (
            .O(N__84806),
            .I(N__84765));
    LocalMux I__19952 (
            .O(N__84803),
            .I(N__84762));
    Span4Mux_v I__19951 (
            .O(N__84800),
            .I(N__84758));
    LocalMux I__19950 (
            .O(N__84797),
            .I(N__84753));
    LocalMux I__19949 (
            .O(N__84794),
            .I(N__84753));
    LocalMux I__19948 (
            .O(N__84791),
            .I(N__84748));
    Span4Mux_v I__19947 (
            .O(N__84788),
            .I(N__84748));
    InMux I__19946 (
            .O(N__84787),
            .I(N__84745));
    InMux I__19945 (
            .O(N__84786),
            .I(N__84740));
    InMux I__19944 (
            .O(N__84785),
            .I(N__84740));
    Span4Mux_h I__19943 (
            .O(N__84782),
            .I(N__84735));
    LocalMux I__19942 (
            .O(N__84777),
            .I(N__84735));
    Span4Mux_v I__19941 (
            .O(N__84774),
            .I(N__84732));
    LocalMux I__19940 (
            .O(N__84771),
            .I(N__84729));
    InMux I__19939 (
            .O(N__84770),
            .I(N__84722));
    InMux I__19938 (
            .O(N__84769),
            .I(N__84722));
    InMux I__19937 (
            .O(N__84768),
            .I(N__84722));
    Span12Mux_v I__19936 (
            .O(N__84765),
            .I(N__84719));
    Span4Mux_h I__19935 (
            .O(N__84762),
            .I(N__84716));
    InMux I__19934 (
            .O(N__84761),
            .I(N__84713));
    Span4Mux_v I__19933 (
            .O(N__84758),
            .I(N__84706));
    Span4Mux_h I__19932 (
            .O(N__84753),
            .I(N__84706));
    Span4Mux_h I__19931 (
            .O(N__84748),
            .I(N__84706));
    LocalMux I__19930 (
            .O(N__84745),
            .I(N__84699));
    LocalMux I__19929 (
            .O(N__84740),
            .I(N__84699));
    Sp12to4 I__19928 (
            .O(N__84735),
            .I(N__84699));
    Odrv4 I__19927 (
            .O(N__84732),
            .I(pid_side_N_216));
    Odrv4 I__19926 (
            .O(N__84729),
            .I(pid_side_N_216));
    LocalMux I__19925 (
            .O(N__84722),
            .I(pid_side_N_216));
    Odrv12 I__19924 (
            .O(N__84719),
            .I(pid_side_N_216));
    Odrv4 I__19923 (
            .O(N__84716),
            .I(pid_side_N_216));
    LocalMux I__19922 (
            .O(N__84713),
            .I(pid_side_N_216));
    Odrv4 I__19921 (
            .O(N__84706),
            .I(pid_side_N_216));
    Odrv12 I__19920 (
            .O(N__84699),
            .I(pid_side_N_216));
    CascadeMux I__19919 (
            .O(N__84682),
            .I(N__84679));
    InMux I__19918 (
            .O(N__84679),
            .I(N__84675));
    CascadeMux I__19917 (
            .O(N__84678),
            .I(N__84672));
    LocalMux I__19916 (
            .O(N__84675),
            .I(N__84668));
    InMux I__19915 (
            .O(N__84672),
            .I(N__84663));
    InMux I__19914 (
            .O(N__84671),
            .I(N__84663));
    Span4Mux_v I__19913 (
            .O(N__84668),
            .I(N__84656));
    LocalMux I__19912 (
            .O(N__84663),
            .I(N__84653));
    InMux I__19911 (
            .O(N__84662),
            .I(N__84650));
    InMux I__19910 (
            .O(N__84661),
            .I(N__84647));
    CascadeMux I__19909 (
            .O(N__84660),
            .I(N__84644));
    CascadeMux I__19908 (
            .O(N__84659),
            .I(N__84641));
    Span4Mux_v I__19907 (
            .O(N__84656),
            .I(N__84638));
    Span4Mux_v I__19906 (
            .O(N__84653),
            .I(N__84635));
    LocalMux I__19905 (
            .O(N__84650),
            .I(N__84632));
    LocalMux I__19904 (
            .O(N__84647),
            .I(N__84629));
    InMux I__19903 (
            .O(N__84644),
            .I(N__84623));
    InMux I__19902 (
            .O(N__84641),
            .I(N__84623));
    Sp12to4 I__19901 (
            .O(N__84638),
            .I(N__84616));
    Sp12to4 I__19900 (
            .O(N__84635),
            .I(N__84616));
    Span12Mux_v I__19899 (
            .O(N__84632),
            .I(N__84616));
    Span12Mux_s1_h I__19898 (
            .O(N__84629),
            .I(N__84613));
    InMux I__19897 (
            .O(N__84628),
            .I(N__84610));
    LocalMux I__19896 (
            .O(N__84623),
            .I(N__84607));
    Span12Mux_h I__19895 (
            .O(N__84616),
            .I(N__84602));
    Span12Mux_h I__19894 (
            .O(N__84613),
            .I(N__84602));
    LocalMux I__19893 (
            .O(N__84610),
            .I(drone_H_disp_front_0));
    Odrv4 I__19892 (
            .O(N__84607),
            .I(drone_H_disp_front_0));
    Odrv12 I__19891 (
            .O(N__84602),
            .I(drone_H_disp_front_0));
    InMux I__19890 (
            .O(N__84595),
            .I(N__84592));
    LocalMux I__19889 (
            .O(N__84592),
            .I(N__84589));
    Span4Mux_v I__19888 (
            .O(N__84589),
            .I(N__84586));
    Span4Mux_h I__19887 (
            .O(N__84586),
            .I(N__84583));
    Span4Mux_s3_h I__19886 (
            .O(N__84583),
            .I(N__84580));
    Odrv4 I__19885 (
            .O(N__84580),
            .I(\pid_front.m0_2_03 ));
    CascadeMux I__19884 (
            .O(N__84577),
            .I(N__84572));
    InMux I__19883 (
            .O(N__84576),
            .I(N__84565));
    InMux I__19882 (
            .O(N__84575),
            .I(N__84565));
    InMux I__19881 (
            .O(N__84572),
            .I(N__84565));
    LocalMux I__19880 (
            .O(N__84565),
            .I(N__84557));
    InMux I__19879 (
            .O(N__84564),
            .I(N__84554));
    InMux I__19878 (
            .O(N__84563),
            .I(N__84551));
    InMux I__19877 (
            .O(N__84562),
            .I(N__84530));
    InMux I__19876 (
            .O(N__84561),
            .I(N__84530));
    InMux I__19875 (
            .O(N__84560),
            .I(N__84530));
    Span4Mux_v I__19874 (
            .O(N__84557),
            .I(N__84523));
    LocalMux I__19873 (
            .O(N__84554),
            .I(N__84523));
    LocalMux I__19872 (
            .O(N__84551),
            .I(N__84523));
    InMux I__19871 (
            .O(N__84550),
            .I(N__84518));
    InMux I__19870 (
            .O(N__84549),
            .I(N__84510));
    InMux I__19869 (
            .O(N__84548),
            .I(N__84510));
    InMux I__19868 (
            .O(N__84547),
            .I(N__84505));
    InMux I__19867 (
            .O(N__84546),
            .I(N__84501));
    InMux I__19866 (
            .O(N__84545),
            .I(N__84493));
    InMux I__19865 (
            .O(N__84544),
            .I(N__84493));
    InMux I__19864 (
            .O(N__84543),
            .I(N__84493));
    InMux I__19863 (
            .O(N__84542),
            .I(N__84488));
    InMux I__19862 (
            .O(N__84541),
            .I(N__84483));
    InMux I__19861 (
            .O(N__84540),
            .I(N__84478));
    InMux I__19860 (
            .O(N__84539),
            .I(N__84478));
    InMux I__19859 (
            .O(N__84538),
            .I(N__84470));
    InMux I__19858 (
            .O(N__84537),
            .I(N__84465));
    LocalMux I__19857 (
            .O(N__84530),
            .I(N__84460));
    Span4Mux_v I__19856 (
            .O(N__84523),
            .I(N__84460));
    InMux I__19855 (
            .O(N__84522),
            .I(N__84457));
    InMux I__19854 (
            .O(N__84521),
            .I(N__84454));
    LocalMux I__19853 (
            .O(N__84518),
            .I(N__84451));
    InMux I__19852 (
            .O(N__84517),
            .I(N__84444));
    InMux I__19851 (
            .O(N__84516),
            .I(N__84444));
    InMux I__19850 (
            .O(N__84515),
            .I(N__84444));
    LocalMux I__19849 (
            .O(N__84510),
            .I(N__84441));
    InMux I__19848 (
            .O(N__84509),
            .I(N__84436));
    InMux I__19847 (
            .O(N__84508),
            .I(N__84436));
    LocalMux I__19846 (
            .O(N__84505),
            .I(N__84429));
    InMux I__19845 (
            .O(N__84504),
            .I(N__84426));
    LocalMux I__19844 (
            .O(N__84501),
            .I(N__84423));
    InMux I__19843 (
            .O(N__84500),
            .I(N__84420));
    LocalMux I__19842 (
            .O(N__84493),
            .I(N__84416));
    InMux I__19841 (
            .O(N__84492),
            .I(N__84408));
    InMux I__19840 (
            .O(N__84491),
            .I(N__84408));
    LocalMux I__19839 (
            .O(N__84488),
            .I(N__84405));
    InMux I__19838 (
            .O(N__84487),
            .I(N__84398));
    InMux I__19837 (
            .O(N__84486),
            .I(N__84395));
    LocalMux I__19836 (
            .O(N__84483),
            .I(N__84390));
    LocalMux I__19835 (
            .O(N__84478),
            .I(N__84390));
    InMux I__19834 (
            .O(N__84477),
            .I(N__84385));
    InMux I__19833 (
            .O(N__84476),
            .I(N__84385));
    InMux I__19832 (
            .O(N__84475),
            .I(N__84378));
    InMux I__19831 (
            .O(N__84474),
            .I(N__84378));
    InMux I__19830 (
            .O(N__84473),
            .I(N__84378));
    LocalMux I__19829 (
            .O(N__84470),
            .I(N__84375));
    InMux I__19828 (
            .O(N__84469),
            .I(N__84370));
    InMux I__19827 (
            .O(N__84468),
            .I(N__84370));
    LocalMux I__19826 (
            .O(N__84465),
            .I(N__84367));
    Span4Mux_h I__19825 (
            .O(N__84460),
            .I(N__84362));
    LocalMux I__19824 (
            .O(N__84457),
            .I(N__84362));
    LocalMux I__19823 (
            .O(N__84454),
            .I(N__84355));
    Span4Mux_v I__19822 (
            .O(N__84451),
            .I(N__84355));
    LocalMux I__19821 (
            .O(N__84444),
            .I(N__84355));
    Span4Mux_v I__19820 (
            .O(N__84441),
            .I(N__84350));
    LocalMux I__19819 (
            .O(N__84436),
            .I(N__84350));
    InMux I__19818 (
            .O(N__84435),
            .I(N__84345));
    InMux I__19817 (
            .O(N__84434),
            .I(N__84345));
    InMux I__19816 (
            .O(N__84433),
            .I(N__84342));
    InMux I__19815 (
            .O(N__84432),
            .I(N__84339));
    Span4Mux_v I__19814 (
            .O(N__84429),
            .I(N__84330));
    LocalMux I__19813 (
            .O(N__84426),
            .I(N__84330));
    Span4Mux_v I__19812 (
            .O(N__84423),
            .I(N__84330));
    LocalMux I__19811 (
            .O(N__84420),
            .I(N__84330));
    InMux I__19810 (
            .O(N__84419),
            .I(N__84327));
    Span4Mux_v I__19809 (
            .O(N__84416),
            .I(N__84324));
    InMux I__19808 (
            .O(N__84415),
            .I(N__84316));
    InMux I__19807 (
            .O(N__84414),
            .I(N__84316));
    InMux I__19806 (
            .O(N__84413),
            .I(N__84313));
    LocalMux I__19805 (
            .O(N__84408),
            .I(N__84308));
    Span4Mux_v I__19804 (
            .O(N__84405),
            .I(N__84308));
    InMux I__19803 (
            .O(N__84404),
            .I(N__84303));
    InMux I__19802 (
            .O(N__84403),
            .I(N__84303));
    InMux I__19801 (
            .O(N__84402),
            .I(N__84298));
    InMux I__19800 (
            .O(N__84401),
            .I(N__84298));
    LocalMux I__19799 (
            .O(N__84398),
            .I(N__84287));
    LocalMux I__19798 (
            .O(N__84395),
            .I(N__84287));
    Span4Mux_h I__19797 (
            .O(N__84390),
            .I(N__84287));
    LocalMux I__19796 (
            .O(N__84385),
            .I(N__84287));
    LocalMux I__19795 (
            .O(N__84378),
            .I(N__84287));
    Span4Mux_v I__19794 (
            .O(N__84375),
            .I(N__84284));
    LocalMux I__19793 (
            .O(N__84370),
            .I(N__84281));
    Span4Mux_v I__19792 (
            .O(N__84367),
            .I(N__84278));
    Span4Mux_v I__19791 (
            .O(N__84362),
            .I(N__84267));
    Span4Mux_v I__19790 (
            .O(N__84355),
            .I(N__84267));
    Span4Mux_h I__19789 (
            .O(N__84350),
            .I(N__84267));
    LocalMux I__19788 (
            .O(N__84345),
            .I(N__84267));
    LocalMux I__19787 (
            .O(N__84342),
            .I(N__84267));
    LocalMux I__19786 (
            .O(N__84339),
            .I(N__84260));
    Span4Mux_v I__19785 (
            .O(N__84330),
            .I(N__84260));
    LocalMux I__19784 (
            .O(N__84327),
            .I(N__84260));
    Span4Mux_v I__19783 (
            .O(N__84324),
            .I(N__84257));
    InMux I__19782 (
            .O(N__84323),
            .I(N__84252));
    InMux I__19781 (
            .O(N__84322),
            .I(N__84249));
    InMux I__19780 (
            .O(N__84321),
            .I(N__84246));
    LocalMux I__19779 (
            .O(N__84316),
            .I(N__84233));
    LocalMux I__19778 (
            .O(N__84313),
            .I(N__84233));
    Sp12to4 I__19777 (
            .O(N__84308),
            .I(N__84233));
    LocalMux I__19776 (
            .O(N__84303),
            .I(N__84233));
    LocalMux I__19775 (
            .O(N__84298),
            .I(N__84233));
    Sp12to4 I__19774 (
            .O(N__84287),
            .I(N__84233));
    Span4Mux_h I__19773 (
            .O(N__84284),
            .I(N__84224));
    Span4Mux_v I__19772 (
            .O(N__84281),
            .I(N__84224));
    Span4Mux_h I__19771 (
            .O(N__84278),
            .I(N__84224));
    Span4Mux_v I__19770 (
            .O(N__84267),
            .I(N__84224));
    Span4Mux_v I__19769 (
            .O(N__84260),
            .I(N__84219));
    Span4Mux_h I__19768 (
            .O(N__84257),
            .I(N__84219));
    InMux I__19767 (
            .O(N__84256),
            .I(N__84214));
    InMux I__19766 (
            .O(N__84255),
            .I(N__84214));
    LocalMux I__19765 (
            .O(N__84252),
            .I(xy_ki_4));
    LocalMux I__19764 (
            .O(N__84249),
            .I(xy_ki_4));
    LocalMux I__19763 (
            .O(N__84246),
            .I(xy_ki_4));
    Odrv12 I__19762 (
            .O(N__84233),
            .I(xy_ki_4));
    Odrv4 I__19761 (
            .O(N__84224),
            .I(xy_ki_4));
    Odrv4 I__19760 (
            .O(N__84219),
            .I(xy_ki_4));
    LocalMux I__19759 (
            .O(N__84214),
            .I(xy_ki_4));
    InMux I__19758 (
            .O(N__84199),
            .I(N__84196));
    LocalMux I__19757 (
            .O(N__84196),
            .I(\pid_side.error_i_reg_9_sx_18 ));
    CascadeMux I__19756 (
            .O(N__84193),
            .I(N__84189));
    InMux I__19755 (
            .O(N__84192),
            .I(N__84183));
    InMux I__19754 (
            .O(N__84189),
            .I(N__84175));
    InMux I__19753 (
            .O(N__84188),
            .I(N__84172));
    CascadeMux I__19752 (
            .O(N__84187),
            .I(N__84169));
    CascadeMux I__19751 (
            .O(N__84186),
            .I(N__84165));
    LocalMux I__19750 (
            .O(N__84183),
            .I(N__84162));
    CascadeMux I__19749 (
            .O(N__84182),
            .I(N__84159));
    InMux I__19748 (
            .O(N__84181),
            .I(N__84155));
    InMux I__19747 (
            .O(N__84180),
            .I(N__84150));
    InMux I__19746 (
            .O(N__84179),
            .I(N__84150));
    InMux I__19745 (
            .O(N__84178),
            .I(N__84147));
    LocalMux I__19744 (
            .O(N__84175),
            .I(N__84144));
    LocalMux I__19743 (
            .O(N__84172),
            .I(N__84141));
    InMux I__19742 (
            .O(N__84169),
            .I(N__84138));
    CascadeMux I__19741 (
            .O(N__84168),
            .I(N__84135));
    InMux I__19740 (
            .O(N__84165),
            .I(N__84129));
    Span4Mux_v I__19739 (
            .O(N__84162),
            .I(N__84126));
    InMux I__19738 (
            .O(N__84159),
            .I(N__84123));
    CascadeMux I__19737 (
            .O(N__84158),
            .I(N__84120));
    LocalMux I__19736 (
            .O(N__84155),
            .I(N__84113));
    LocalMux I__19735 (
            .O(N__84150),
            .I(N__84108));
    LocalMux I__19734 (
            .O(N__84147),
            .I(N__84108));
    Span4Mux_v I__19733 (
            .O(N__84144),
            .I(N__84101));
    Span4Mux_h I__19732 (
            .O(N__84141),
            .I(N__84101));
    LocalMux I__19731 (
            .O(N__84138),
            .I(N__84101));
    InMux I__19730 (
            .O(N__84135),
            .I(N__84097));
    CascadeMux I__19729 (
            .O(N__84134),
            .I(N__84094));
    InMux I__19728 (
            .O(N__84133),
            .I(N__84088));
    CascadeMux I__19727 (
            .O(N__84132),
            .I(N__84084));
    LocalMux I__19726 (
            .O(N__84129),
            .I(N__84078));
    Span4Mux_h I__19725 (
            .O(N__84126),
            .I(N__84073));
    LocalMux I__19724 (
            .O(N__84123),
            .I(N__84073));
    InMux I__19723 (
            .O(N__84120),
            .I(N__84070));
    InMux I__19722 (
            .O(N__84119),
            .I(N__84067));
    CascadeMux I__19721 (
            .O(N__84118),
            .I(N__84064));
    CascadeMux I__19720 (
            .O(N__84117),
            .I(N__84060));
    CascadeMux I__19719 (
            .O(N__84116),
            .I(N__84057));
    Span4Mux_h I__19718 (
            .O(N__84113),
            .I(N__84053));
    Span4Mux_h I__19717 (
            .O(N__84108),
            .I(N__84048));
    Span4Mux_v I__19716 (
            .O(N__84101),
            .I(N__84048));
    InMux I__19715 (
            .O(N__84100),
            .I(N__84045));
    LocalMux I__19714 (
            .O(N__84097),
            .I(N__84042));
    InMux I__19713 (
            .O(N__84094),
            .I(N__84039));
    InMux I__19712 (
            .O(N__84093),
            .I(N__84036));
    InMux I__19711 (
            .O(N__84092),
            .I(N__84031));
    InMux I__19710 (
            .O(N__84091),
            .I(N__84031));
    LocalMux I__19709 (
            .O(N__84088),
            .I(N__84028));
    InMux I__19708 (
            .O(N__84087),
            .I(N__84024));
    InMux I__19707 (
            .O(N__84084),
            .I(N__84019));
    InMux I__19706 (
            .O(N__84083),
            .I(N__84019));
    InMux I__19705 (
            .O(N__84082),
            .I(N__84014));
    InMux I__19704 (
            .O(N__84081),
            .I(N__84014));
    Span4Mux_h I__19703 (
            .O(N__84078),
            .I(N__84011));
    Span4Mux_v I__19702 (
            .O(N__84073),
            .I(N__84008));
    LocalMux I__19701 (
            .O(N__84070),
            .I(N__84003));
    LocalMux I__19700 (
            .O(N__84067),
            .I(N__84003));
    InMux I__19699 (
            .O(N__84064),
            .I(N__83996));
    InMux I__19698 (
            .O(N__84063),
            .I(N__83996));
    InMux I__19697 (
            .O(N__84060),
            .I(N__83996));
    InMux I__19696 (
            .O(N__84057),
            .I(N__83993));
    InMux I__19695 (
            .O(N__84056),
            .I(N__83990));
    Span4Mux_h I__19694 (
            .O(N__84053),
            .I(N__83983));
    Span4Mux_h I__19693 (
            .O(N__84048),
            .I(N__83983));
    LocalMux I__19692 (
            .O(N__84045),
            .I(N__83983));
    Span4Mux_v I__19691 (
            .O(N__84042),
            .I(N__83978));
    LocalMux I__19690 (
            .O(N__84039),
            .I(N__83978));
    LocalMux I__19689 (
            .O(N__84036),
            .I(N__83973));
    LocalMux I__19688 (
            .O(N__84031),
            .I(N__83973));
    Span4Mux_h I__19687 (
            .O(N__84028),
            .I(N__83970));
    CascadeMux I__19686 (
            .O(N__84027),
            .I(N__83967));
    LocalMux I__19685 (
            .O(N__84024),
            .I(N__83964));
    LocalMux I__19684 (
            .O(N__84019),
            .I(N__83959));
    LocalMux I__19683 (
            .O(N__84014),
            .I(N__83959));
    Span4Mux_v I__19682 (
            .O(N__84011),
            .I(N__83952));
    Span4Mux_h I__19681 (
            .O(N__84008),
            .I(N__83952));
    Span4Mux_h I__19680 (
            .O(N__84003),
            .I(N__83952));
    LocalMux I__19679 (
            .O(N__83996),
            .I(N__83949));
    LocalMux I__19678 (
            .O(N__83993),
            .I(N__83938));
    LocalMux I__19677 (
            .O(N__83990),
            .I(N__83938));
    Span4Mux_v I__19676 (
            .O(N__83983),
            .I(N__83938));
    Span4Mux_h I__19675 (
            .O(N__83978),
            .I(N__83938));
    Span4Mux_v I__19674 (
            .O(N__83973),
            .I(N__83938));
    Span4Mux_v I__19673 (
            .O(N__83970),
            .I(N__83935));
    InMux I__19672 (
            .O(N__83967),
            .I(N__83932));
    Span4Mux_v I__19671 (
            .O(N__83964),
            .I(N__83927));
    Span4Mux_v I__19670 (
            .O(N__83959),
            .I(N__83927));
    Span4Mux_h I__19669 (
            .O(N__83952),
            .I(N__83924));
    Span12Mux_h I__19668 (
            .O(N__83949),
            .I(N__83921));
    Span4Mux_h I__19667 (
            .O(N__83938),
            .I(N__83918));
    Odrv4 I__19666 (
            .O(N__83935),
            .I(xy_ki_2));
    LocalMux I__19665 (
            .O(N__83932),
            .I(xy_ki_2));
    Odrv4 I__19664 (
            .O(N__83927),
            .I(xy_ki_2));
    Odrv4 I__19663 (
            .O(N__83924),
            .I(xy_ki_2));
    Odrv12 I__19662 (
            .O(N__83921),
            .I(xy_ki_2));
    Odrv4 I__19661 (
            .O(N__83918),
            .I(xy_ki_2));
    CEMux I__19660 (
            .O(N__83905),
            .I(N__83902));
    LocalMux I__19659 (
            .O(N__83902),
            .I(N__83895));
    CEMux I__19658 (
            .O(N__83901),
            .I(N__83891));
    CEMux I__19657 (
            .O(N__83900),
            .I(N__83885));
    CEMux I__19656 (
            .O(N__83899),
            .I(N__83882));
    CEMux I__19655 (
            .O(N__83898),
            .I(N__83879));
    Span4Mux_v I__19654 (
            .O(N__83895),
            .I(N__83874));
    CEMux I__19653 (
            .O(N__83894),
            .I(N__83871));
    LocalMux I__19652 (
            .O(N__83891),
            .I(N__83868));
    CEMux I__19651 (
            .O(N__83890),
            .I(N__83865));
    CEMux I__19650 (
            .O(N__83889),
            .I(N__83862));
    CEMux I__19649 (
            .O(N__83888),
            .I(N__83859));
    LocalMux I__19648 (
            .O(N__83885),
            .I(N__83856));
    LocalMux I__19647 (
            .O(N__83882),
            .I(N__83851));
    LocalMux I__19646 (
            .O(N__83879),
            .I(N__83851));
    CEMux I__19645 (
            .O(N__83878),
            .I(N__83848));
    CEMux I__19644 (
            .O(N__83877),
            .I(N__83845));
    Span4Mux_v I__19643 (
            .O(N__83874),
            .I(N__83840));
    LocalMux I__19642 (
            .O(N__83871),
            .I(N__83840));
    Span4Mux_v I__19641 (
            .O(N__83868),
            .I(N__83837));
    LocalMux I__19640 (
            .O(N__83865),
            .I(N__83834));
    LocalMux I__19639 (
            .O(N__83862),
            .I(N__83831));
    LocalMux I__19638 (
            .O(N__83859),
            .I(N__83824));
    Span4Mux_v I__19637 (
            .O(N__83856),
            .I(N__83824));
    Span4Mux_h I__19636 (
            .O(N__83851),
            .I(N__83824));
    LocalMux I__19635 (
            .O(N__83848),
            .I(N__83821));
    LocalMux I__19634 (
            .O(N__83845),
            .I(N__83818));
    Span4Mux_h I__19633 (
            .O(N__83840),
            .I(N__83815));
    Span4Mux_v I__19632 (
            .O(N__83837),
            .I(N__83812));
    Span4Mux_h I__19631 (
            .O(N__83834),
            .I(N__83809));
    Span4Mux_h I__19630 (
            .O(N__83831),
            .I(N__83806));
    Span4Mux_h I__19629 (
            .O(N__83824),
            .I(N__83803));
    Span4Mux_h I__19628 (
            .O(N__83821),
            .I(N__83798));
    Span4Mux_v I__19627 (
            .O(N__83818),
            .I(N__83798));
    Span4Mux_h I__19626 (
            .O(N__83815),
            .I(N__83795));
    Span4Mux_h I__19625 (
            .O(N__83812),
            .I(N__83792));
    Span4Mux_h I__19624 (
            .O(N__83809),
            .I(N__83787));
    Span4Mux_v I__19623 (
            .O(N__83806),
            .I(N__83787));
    Span4Mux_h I__19622 (
            .O(N__83803),
            .I(N__83784));
    Span4Mux_v I__19621 (
            .O(N__83798),
            .I(N__83781));
    Span4Mux_v I__19620 (
            .O(N__83795),
            .I(N__83778));
    Span4Mux_h I__19619 (
            .O(N__83792),
            .I(N__83775));
    Span4Mux_h I__19618 (
            .O(N__83787),
            .I(N__83772));
    Span4Mux_v I__19617 (
            .O(N__83784),
            .I(N__83769));
    Sp12to4 I__19616 (
            .O(N__83781),
            .I(N__83766));
    Sp12to4 I__19615 (
            .O(N__83778),
            .I(N__83763));
    Odrv4 I__19614 (
            .O(N__83775),
            .I(\Commands_frame_decoder.source_xy_ki_1_sqmuxa_0 ));
    Odrv4 I__19613 (
            .O(N__83772),
            .I(\Commands_frame_decoder.source_xy_ki_1_sqmuxa_0 ));
    Odrv4 I__19612 (
            .O(N__83769),
            .I(\Commands_frame_decoder.source_xy_ki_1_sqmuxa_0 ));
    Odrv12 I__19611 (
            .O(N__83766),
            .I(\Commands_frame_decoder.source_xy_ki_1_sqmuxa_0 ));
    Odrv12 I__19610 (
            .O(N__83763),
            .I(\Commands_frame_decoder.source_xy_ki_1_sqmuxa_0 ));
    CascadeMux I__19609 (
            .O(N__83752),
            .I(N__83749));
    InMux I__19608 (
            .O(N__83749),
            .I(N__83746));
    LocalMux I__19607 (
            .O(N__83746),
            .I(N__83743));
    Odrv12 I__19606 (
            .O(N__83743),
            .I(side_command_0));
    InMux I__19605 (
            .O(N__83740),
            .I(N__83737));
    LocalMux I__19604 (
            .O(N__83737),
            .I(N__83734));
    Span4Mux_h I__19603 (
            .O(N__83734),
            .I(N__83731));
    Span4Mux_v I__19602 (
            .O(N__83731),
            .I(N__83728));
    Odrv4 I__19601 (
            .O(N__83728),
            .I(\pid_side.O_1_14 ));
    InMux I__19600 (
            .O(N__83725),
            .I(N__83716));
    InMux I__19599 (
            .O(N__83724),
            .I(N__83716));
    InMux I__19598 (
            .O(N__83723),
            .I(N__83709));
    InMux I__19597 (
            .O(N__83722),
            .I(N__83709));
    InMux I__19596 (
            .O(N__83721),
            .I(N__83709));
    LocalMux I__19595 (
            .O(N__83716),
            .I(\pid_side.error_d_regZ0Z_11 ));
    LocalMux I__19594 (
            .O(N__83709),
            .I(\pid_side.error_d_regZ0Z_11 ));
    InMux I__19593 (
            .O(N__83704),
            .I(N__83701));
    LocalMux I__19592 (
            .O(N__83701),
            .I(\pid_side.m24_2_03_0 ));
    CascadeMux I__19591 (
            .O(N__83698),
            .I(N__83695));
    InMux I__19590 (
            .O(N__83695),
            .I(N__83692));
    LocalMux I__19589 (
            .O(N__83692),
            .I(N__83689));
    Span4Mux_h I__19588 (
            .O(N__83689),
            .I(N__83686));
    Span4Mux_h I__19587 (
            .O(N__83686),
            .I(N__83683));
    Odrv4 I__19586 (
            .O(N__83683),
            .I(\pid_side.error_i_regZ0Z_20 ));
    InMux I__19585 (
            .O(N__83680),
            .I(N__83677));
    LocalMux I__19584 (
            .O(N__83677),
            .I(N__83672));
    InMux I__19583 (
            .O(N__83676),
            .I(N__83669));
    InMux I__19582 (
            .O(N__83675),
            .I(N__83666));
    Span4Mux_h I__19581 (
            .O(N__83672),
            .I(N__83663));
    LocalMux I__19580 (
            .O(N__83669),
            .I(N__83660));
    LocalMux I__19579 (
            .O(N__83666),
            .I(N__83656));
    Span4Mux_h I__19578 (
            .O(N__83663),
            .I(N__83651));
    Span4Mux_h I__19577 (
            .O(N__83660),
            .I(N__83651));
    InMux I__19576 (
            .O(N__83659),
            .I(N__83648));
    Odrv4 I__19575 (
            .O(N__83656),
            .I(\pid_side.N_156 ));
    Odrv4 I__19574 (
            .O(N__83651),
            .I(\pid_side.N_156 ));
    LocalMux I__19573 (
            .O(N__83648),
            .I(\pid_side.N_156 ));
    InMux I__19572 (
            .O(N__83641),
            .I(N__83632));
    InMux I__19571 (
            .O(N__83640),
            .I(N__83629));
    InMux I__19570 (
            .O(N__83639),
            .I(N__83625));
    InMux I__19569 (
            .O(N__83638),
            .I(N__83620));
    InMux I__19568 (
            .O(N__83637),
            .I(N__83620));
    InMux I__19567 (
            .O(N__83636),
            .I(N__83617));
    InMux I__19566 (
            .O(N__83635),
            .I(N__83614));
    LocalMux I__19565 (
            .O(N__83632),
            .I(N__83611));
    LocalMux I__19564 (
            .O(N__83629),
            .I(N__83608));
    InMux I__19563 (
            .O(N__83628),
            .I(N__83605));
    LocalMux I__19562 (
            .O(N__83625),
            .I(N__83600));
    LocalMux I__19561 (
            .O(N__83620),
            .I(N__83600));
    LocalMux I__19560 (
            .O(N__83617),
            .I(N__83597));
    LocalMux I__19559 (
            .O(N__83614),
            .I(N__83592));
    Span4Mux_s1_h I__19558 (
            .O(N__83611),
            .I(N__83592));
    Span4Mux_s1_h I__19557 (
            .O(N__83608),
            .I(N__83589));
    LocalMux I__19556 (
            .O(N__83605),
            .I(N__83585));
    Span4Mux_h I__19555 (
            .O(N__83600),
            .I(N__83582));
    Span4Mux_h I__19554 (
            .O(N__83597),
            .I(N__83577));
    Span4Mux_h I__19553 (
            .O(N__83592),
            .I(N__83577));
    Span4Mux_h I__19552 (
            .O(N__83589),
            .I(N__83574));
    InMux I__19551 (
            .O(N__83588),
            .I(N__83571));
    Odrv4 I__19550 (
            .O(N__83585),
            .I(\pid_side.error_7 ));
    Odrv4 I__19549 (
            .O(N__83582),
            .I(\pid_side.error_7 ));
    Odrv4 I__19548 (
            .O(N__83577),
            .I(\pid_side.error_7 ));
    Odrv4 I__19547 (
            .O(N__83574),
            .I(\pid_side.error_7 ));
    LocalMux I__19546 (
            .O(N__83571),
            .I(\pid_side.error_7 ));
    CascadeMux I__19545 (
            .O(N__83560),
            .I(\pid_side.N_551_cascade_ ));
    InMux I__19544 (
            .O(N__83557),
            .I(N__83554));
    LocalMux I__19543 (
            .O(N__83554),
            .I(\pid_side.m8_2_03_3_i_0 ));
    InMux I__19542 (
            .O(N__83551),
            .I(N__83545));
    InMux I__19541 (
            .O(N__83550),
            .I(N__83545));
    LocalMux I__19540 (
            .O(N__83545),
            .I(N__83542));
    Span4Mux_h I__19539 (
            .O(N__83542),
            .I(N__83539));
    Span4Mux_h I__19538 (
            .O(N__83539),
            .I(N__83535));
    InMux I__19537 (
            .O(N__83538),
            .I(N__83532));
    Odrv4 I__19536 (
            .O(N__83535),
            .I(\pid_side.N_230 ));
    LocalMux I__19535 (
            .O(N__83532),
            .I(\pid_side.N_230 ));
    CascadeMux I__19534 (
            .O(N__83527),
            .I(N__83524));
    InMux I__19533 (
            .O(N__83524),
            .I(N__83519));
    CascadeMux I__19532 (
            .O(N__83523),
            .I(N__83516));
    CascadeMux I__19531 (
            .O(N__83522),
            .I(N__83511));
    LocalMux I__19530 (
            .O(N__83519),
            .I(N__83507));
    InMux I__19529 (
            .O(N__83516),
            .I(N__83497));
    InMux I__19528 (
            .O(N__83515),
            .I(N__83497));
    InMux I__19527 (
            .O(N__83514),
            .I(N__83497));
    InMux I__19526 (
            .O(N__83511),
            .I(N__83497));
    CascadeMux I__19525 (
            .O(N__83510),
            .I(N__83493));
    Span4Mux_v I__19524 (
            .O(N__83507),
            .I(N__83488));
    InMux I__19523 (
            .O(N__83506),
            .I(N__83485));
    LocalMux I__19522 (
            .O(N__83497),
            .I(N__83482));
    InMux I__19521 (
            .O(N__83496),
            .I(N__83478));
    InMux I__19520 (
            .O(N__83493),
            .I(N__83470));
    InMux I__19519 (
            .O(N__83492),
            .I(N__83470));
    InMux I__19518 (
            .O(N__83491),
            .I(N__83467));
    Span4Mux_v I__19517 (
            .O(N__83488),
            .I(N__83462));
    LocalMux I__19516 (
            .O(N__83485),
            .I(N__83462));
    Span4Mux_v I__19515 (
            .O(N__83482),
            .I(N__83459));
    InMux I__19514 (
            .O(N__83481),
            .I(N__83456));
    LocalMux I__19513 (
            .O(N__83478),
            .I(N__83453));
    InMux I__19512 (
            .O(N__83477),
            .I(N__83450));
    InMux I__19511 (
            .O(N__83476),
            .I(N__83447));
    InMux I__19510 (
            .O(N__83475),
            .I(N__83444));
    LocalMux I__19509 (
            .O(N__83470),
            .I(N__83441));
    LocalMux I__19508 (
            .O(N__83467),
            .I(N__83438));
    Span4Mux_v I__19507 (
            .O(N__83462),
            .I(N__83435));
    Span4Mux_h I__19506 (
            .O(N__83459),
            .I(N__83430));
    LocalMux I__19505 (
            .O(N__83456),
            .I(N__83430));
    Span4Mux_h I__19504 (
            .O(N__83453),
            .I(N__83427));
    LocalMux I__19503 (
            .O(N__83450),
            .I(N__83422));
    LocalMux I__19502 (
            .O(N__83447),
            .I(N__83422));
    LocalMux I__19501 (
            .O(N__83444),
            .I(N__83419));
    Span4Mux_v I__19500 (
            .O(N__83441),
            .I(N__83412));
    Span4Mux_v I__19499 (
            .O(N__83438),
            .I(N__83412));
    Span4Mux_h I__19498 (
            .O(N__83435),
            .I(N__83412));
    Span4Mux_v I__19497 (
            .O(N__83430),
            .I(N__83409));
    Span4Mux_h I__19496 (
            .O(N__83427),
            .I(N__83406));
    Span4Mux_v I__19495 (
            .O(N__83422),
            .I(N__83403));
    Span12Mux_v I__19494 (
            .O(N__83419),
            .I(N__83400));
    Odrv4 I__19493 (
            .O(N__83412),
            .I(pid_side_N_496));
    Odrv4 I__19492 (
            .O(N__83409),
            .I(pid_side_N_496));
    Odrv4 I__19491 (
            .O(N__83406),
            .I(pid_side_N_496));
    Odrv4 I__19490 (
            .O(N__83403),
            .I(pid_side_N_496));
    Odrv12 I__19489 (
            .O(N__83400),
            .I(pid_side_N_496));
    InMux I__19488 (
            .O(N__83389),
            .I(N__83386));
    LocalMux I__19487 (
            .O(N__83386),
            .I(\pid_side.N_551 ));
    CascadeMux I__19486 (
            .O(N__83383),
            .I(\pid_side.error_i_reg_esr_RNO_0Z0Z_4_cascade_ ));
    InMux I__19485 (
            .O(N__83380),
            .I(N__83371));
    InMux I__19484 (
            .O(N__83379),
            .I(N__83362));
    InMux I__19483 (
            .O(N__83378),
            .I(N__83359));
    InMux I__19482 (
            .O(N__83377),
            .I(N__83356));
    InMux I__19481 (
            .O(N__83376),
            .I(N__83351));
    CascadeMux I__19480 (
            .O(N__83375),
            .I(N__83347));
    CascadeMux I__19479 (
            .O(N__83374),
            .I(N__83344));
    LocalMux I__19478 (
            .O(N__83371),
            .I(N__83341));
    InMux I__19477 (
            .O(N__83370),
            .I(N__83334));
    InMux I__19476 (
            .O(N__83369),
            .I(N__83334));
    InMux I__19475 (
            .O(N__83368),
            .I(N__83334));
    InMux I__19474 (
            .O(N__83367),
            .I(N__83331));
    InMux I__19473 (
            .O(N__83366),
            .I(N__83328));
    InMux I__19472 (
            .O(N__83365),
            .I(N__83325));
    LocalMux I__19471 (
            .O(N__83362),
            .I(N__83320));
    LocalMux I__19470 (
            .O(N__83359),
            .I(N__83320));
    LocalMux I__19469 (
            .O(N__83356),
            .I(N__83315));
    InMux I__19468 (
            .O(N__83355),
            .I(N__83312));
    InMux I__19467 (
            .O(N__83354),
            .I(N__83308));
    LocalMux I__19466 (
            .O(N__83351),
            .I(N__83305));
    InMux I__19465 (
            .O(N__83350),
            .I(N__83302));
    InMux I__19464 (
            .O(N__83347),
            .I(N__83297));
    InMux I__19463 (
            .O(N__83344),
            .I(N__83297));
    Span4Mux_v I__19462 (
            .O(N__83341),
            .I(N__83292));
    LocalMux I__19461 (
            .O(N__83334),
            .I(N__83292));
    LocalMux I__19460 (
            .O(N__83331),
            .I(N__83289));
    LocalMux I__19459 (
            .O(N__83328),
            .I(N__83286));
    LocalMux I__19458 (
            .O(N__83325),
            .I(N__83283));
    Span4Mux_v I__19457 (
            .O(N__83320),
            .I(N__83280));
    InMux I__19456 (
            .O(N__83319),
            .I(N__83275));
    InMux I__19455 (
            .O(N__83318),
            .I(N__83275));
    Span4Mux_h I__19454 (
            .O(N__83315),
            .I(N__83272));
    LocalMux I__19453 (
            .O(N__83312),
            .I(N__83269));
    CascadeMux I__19452 (
            .O(N__83311),
            .I(N__83264));
    LocalMux I__19451 (
            .O(N__83308),
            .I(N__83261));
    Span4Mux_h I__19450 (
            .O(N__83305),
            .I(N__83252));
    LocalMux I__19449 (
            .O(N__83302),
            .I(N__83252));
    LocalMux I__19448 (
            .O(N__83297),
            .I(N__83252));
    Span4Mux_h I__19447 (
            .O(N__83292),
            .I(N__83252));
    Span4Mux_h I__19446 (
            .O(N__83289),
            .I(N__83249));
    Span4Mux_v I__19445 (
            .O(N__83286),
            .I(N__83246));
    Span4Mux_h I__19444 (
            .O(N__83283),
            .I(N__83239));
    Span4Mux_h I__19443 (
            .O(N__83280),
            .I(N__83239));
    LocalMux I__19442 (
            .O(N__83275),
            .I(N__83239));
    Span4Mux_v I__19441 (
            .O(N__83272),
            .I(N__83236));
    Span12Mux_h I__19440 (
            .O(N__83269),
            .I(N__83233));
    InMux I__19439 (
            .O(N__83268),
            .I(N__83226));
    InMux I__19438 (
            .O(N__83267),
            .I(N__83226));
    InMux I__19437 (
            .O(N__83264),
            .I(N__83226));
    Span4Mux_v I__19436 (
            .O(N__83261),
            .I(N__83221));
    Span4Mux_v I__19435 (
            .O(N__83252),
            .I(N__83221));
    Span4Mux_v I__19434 (
            .O(N__83249),
            .I(N__83214));
    Span4Mux_h I__19433 (
            .O(N__83246),
            .I(N__83214));
    Span4Mux_v I__19432 (
            .O(N__83239),
            .I(N__83214));
    Odrv4 I__19431 (
            .O(N__83236),
            .I(pid_side_N_490));
    Odrv12 I__19430 (
            .O(N__83233),
            .I(pid_side_N_490));
    LocalMux I__19429 (
            .O(N__83226),
            .I(pid_side_N_490));
    Odrv4 I__19428 (
            .O(N__83221),
            .I(pid_side_N_490));
    Odrv4 I__19427 (
            .O(N__83214),
            .I(pid_side_N_490));
    CascadeMux I__19426 (
            .O(N__83203),
            .I(N__83200));
    InMux I__19425 (
            .O(N__83200),
            .I(N__83197));
    LocalMux I__19424 (
            .O(N__83197),
            .I(N__83194));
    Span4Mux_h I__19423 (
            .O(N__83194),
            .I(N__83191));
    Span4Mux_h I__19422 (
            .O(N__83191),
            .I(N__83188));
    Odrv4 I__19421 (
            .O(N__83188),
            .I(\pid_side.error_i_regZ0Z_4 ));
    CascadeMux I__19420 (
            .O(N__83185),
            .I(N__83179));
    CascadeMux I__19419 (
            .O(N__83184),
            .I(N__83171));
    InMux I__19418 (
            .O(N__83183),
            .I(N__83163));
    CascadeMux I__19417 (
            .O(N__83182),
            .I(N__83160));
    InMux I__19416 (
            .O(N__83179),
            .I(N__83157));
    InMux I__19415 (
            .O(N__83178),
            .I(N__83154));
    InMux I__19414 (
            .O(N__83177),
            .I(N__83151));
    CascadeMux I__19413 (
            .O(N__83176),
            .I(N__83147));
    InMux I__19412 (
            .O(N__83175),
            .I(N__83143));
    InMux I__19411 (
            .O(N__83174),
            .I(N__83140));
    InMux I__19410 (
            .O(N__83171),
            .I(N__83133));
    InMux I__19409 (
            .O(N__83170),
            .I(N__83133));
    InMux I__19408 (
            .O(N__83169),
            .I(N__83133));
    InMux I__19407 (
            .O(N__83168),
            .I(N__83125));
    InMux I__19406 (
            .O(N__83167),
            .I(N__83125));
    InMux I__19405 (
            .O(N__83166),
            .I(N__83125));
    LocalMux I__19404 (
            .O(N__83163),
            .I(N__83122));
    InMux I__19403 (
            .O(N__83160),
            .I(N__83119));
    LocalMux I__19402 (
            .O(N__83157),
            .I(N__83114));
    LocalMux I__19401 (
            .O(N__83154),
            .I(N__83114));
    LocalMux I__19400 (
            .O(N__83151),
            .I(N__83111));
    InMux I__19399 (
            .O(N__83150),
            .I(N__83108));
    InMux I__19398 (
            .O(N__83147),
            .I(N__83105));
    InMux I__19397 (
            .O(N__83146),
            .I(N__83102));
    LocalMux I__19396 (
            .O(N__83143),
            .I(N__83099));
    LocalMux I__19395 (
            .O(N__83140),
            .I(N__83094));
    LocalMux I__19394 (
            .O(N__83133),
            .I(N__83094));
    CascadeMux I__19393 (
            .O(N__83132),
            .I(N__83091));
    LocalMux I__19392 (
            .O(N__83125),
            .I(N__83086));
    Span4Mux_v I__19391 (
            .O(N__83122),
            .I(N__83086));
    LocalMux I__19390 (
            .O(N__83119),
            .I(N__83080));
    Span4Mux_v I__19389 (
            .O(N__83114),
            .I(N__83077));
    Span4Mux_v I__19388 (
            .O(N__83111),
            .I(N__83072));
    LocalMux I__19387 (
            .O(N__83108),
            .I(N__83072));
    LocalMux I__19386 (
            .O(N__83105),
            .I(N__83069));
    LocalMux I__19385 (
            .O(N__83102),
            .I(N__83062));
    Span4Mux_v I__19384 (
            .O(N__83099),
            .I(N__83062));
    Span4Mux_v I__19383 (
            .O(N__83094),
            .I(N__83062));
    InMux I__19382 (
            .O(N__83091),
            .I(N__83059));
    Span4Mux_h I__19381 (
            .O(N__83086),
            .I(N__83056));
    InMux I__19380 (
            .O(N__83085),
            .I(N__83049));
    InMux I__19379 (
            .O(N__83084),
            .I(N__83049));
    InMux I__19378 (
            .O(N__83083),
            .I(N__83049));
    Span4Mux_v I__19377 (
            .O(N__83080),
            .I(N__83038));
    Span4Mux_v I__19376 (
            .O(N__83077),
            .I(N__83038));
    Span4Mux_h I__19375 (
            .O(N__83072),
            .I(N__83038));
    Span4Mux_v I__19374 (
            .O(N__83069),
            .I(N__83038));
    Span4Mux_h I__19373 (
            .O(N__83062),
            .I(N__83038));
    LocalMux I__19372 (
            .O(N__83059),
            .I(xy_ki_fast_1));
    Odrv4 I__19371 (
            .O(N__83056),
            .I(xy_ki_fast_1));
    LocalMux I__19370 (
            .O(N__83049),
            .I(xy_ki_fast_1));
    Odrv4 I__19369 (
            .O(N__83038),
            .I(xy_ki_fast_1));
    InMux I__19368 (
            .O(N__83029),
            .I(N__83023));
    InMux I__19367 (
            .O(N__83028),
            .I(N__83020));
    InMux I__19366 (
            .O(N__83027),
            .I(N__83016));
    InMux I__19365 (
            .O(N__83026),
            .I(N__83013));
    LocalMux I__19364 (
            .O(N__83023),
            .I(N__83003));
    LocalMux I__19363 (
            .O(N__83020),
            .I(N__83003));
    InMux I__19362 (
            .O(N__83019),
            .I(N__82993));
    LocalMux I__19361 (
            .O(N__83016),
            .I(N__82988));
    LocalMux I__19360 (
            .O(N__83013),
            .I(N__82988));
    InMux I__19359 (
            .O(N__83012),
            .I(N__82985));
    InMux I__19358 (
            .O(N__83011),
            .I(N__82982));
    InMux I__19357 (
            .O(N__83010),
            .I(N__82979));
    InMux I__19356 (
            .O(N__83009),
            .I(N__82976));
    InMux I__19355 (
            .O(N__83008),
            .I(N__82973));
    Span4Mux_v I__19354 (
            .O(N__83003),
            .I(N__82970));
    InMux I__19353 (
            .O(N__83002),
            .I(N__82967));
    InMux I__19352 (
            .O(N__83001),
            .I(N__82960));
    InMux I__19351 (
            .O(N__83000),
            .I(N__82960));
    InMux I__19350 (
            .O(N__82999),
            .I(N__82960));
    InMux I__19349 (
            .O(N__82998),
            .I(N__82957));
    InMux I__19348 (
            .O(N__82997),
            .I(N__82954));
    InMux I__19347 (
            .O(N__82996),
            .I(N__82951));
    LocalMux I__19346 (
            .O(N__82993),
            .I(N__82946));
    Span4Mux_v I__19345 (
            .O(N__82988),
            .I(N__82946));
    LocalMux I__19344 (
            .O(N__82985),
            .I(N__82940));
    LocalMux I__19343 (
            .O(N__82982),
            .I(N__82933));
    LocalMux I__19342 (
            .O(N__82979),
            .I(N__82933));
    LocalMux I__19341 (
            .O(N__82976),
            .I(N__82933));
    LocalMux I__19340 (
            .O(N__82973),
            .I(N__82930));
    Span4Mux_v I__19339 (
            .O(N__82970),
            .I(N__82925));
    LocalMux I__19338 (
            .O(N__82967),
            .I(N__82925));
    LocalMux I__19337 (
            .O(N__82960),
            .I(N__82920));
    LocalMux I__19336 (
            .O(N__82957),
            .I(N__82920));
    LocalMux I__19335 (
            .O(N__82954),
            .I(N__82915));
    LocalMux I__19334 (
            .O(N__82951),
            .I(N__82915));
    Span4Mux_h I__19333 (
            .O(N__82946),
            .I(N__82912));
    InMux I__19332 (
            .O(N__82945),
            .I(N__82905));
    InMux I__19331 (
            .O(N__82944),
            .I(N__82905));
    InMux I__19330 (
            .O(N__82943),
            .I(N__82905));
    Span4Mux_v I__19329 (
            .O(N__82940),
            .I(N__82894));
    Span4Mux_v I__19328 (
            .O(N__82933),
            .I(N__82894));
    Span4Mux_v I__19327 (
            .O(N__82930),
            .I(N__82894));
    Span4Mux_h I__19326 (
            .O(N__82925),
            .I(N__82894));
    Span4Mux_v I__19325 (
            .O(N__82920),
            .I(N__82894));
    Odrv12 I__19324 (
            .O(N__82915),
            .I(xy_ki_0_rep1));
    Odrv4 I__19323 (
            .O(N__82912),
            .I(xy_ki_0_rep1));
    LocalMux I__19322 (
            .O(N__82905),
            .I(xy_ki_0_rep1));
    Odrv4 I__19321 (
            .O(N__82894),
            .I(xy_ki_0_rep1));
    InMux I__19320 (
            .O(N__82885),
            .I(N__82882));
    LocalMux I__19319 (
            .O(N__82882),
            .I(N__82879));
    Span4Mux_h I__19318 (
            .O(N__82879),
            .I(N__82875));
    InMux I__19317 (
            .O(N__82878),
            .I(N__82872));
    Span4Mux_h I__19316 (
            .O(N__82875),
            .I(N__82867));
    LocalMux I__19315 (
            .O(N__82872),
            .I(N__82867));
    Odrv4 I__19314 (
            .O(N__82867),
            .I(\pid_side.N_183 ));
    CascadeMux I__19313 (
            .O(N__82864),
            .I(\pid_side.N_538_cascade_ ));
    InMux I__19312 (
            .O(N__82861),
            .I(N__82856));
    InMux I__19311 (
            .O(N__82860),
            .I(N__82853));
    InMux I__19310 (
            .O(N__82859),
            .I(N__82847));
    LocalMux I__19309 (
            .O(N__82856),
            .I(N__82844));
    LocalMux I__19308 (
            .O(N__82853),
            .I(N__82841));
    InMux I__19307 (
            .O(N__82852),
            .I(N__82838));
    InMux I__19306 (
            .O(N__82851),
            .I(N__82835));
    InMux I__19305 (
            .O(N__82850),
            .I(N__82832));
    LocalMux I__19304 (
            .O(N__82847),
            .I(N__82829));
    Span4Mux_v I__19303 (
            .O(N__82844),
            .I(N__82824));
    Span4Mux_s0_h I__19302 (
            .O(N__82841),
            .I(N__82821));
    LocalMux I__19301 (
            .O(N__82838),
            .I(N__82815));
    LocalMux I__19300 (
            .O(N__82835),
            .I(N__82815));
    LocalMux I__19299 (
            .O(N__82832),
            .I(N__82812));
    Span4Mux_v I__19298 (
            .O(N__82829),
            .I(N__82809));
    InMux I__19297 (
            .O(N__82828),
            .I(N__82804));
    InMux I__19296 (
            .O(N__82827),
            .I(N__82804));
    Span4Mux_h I__19295 (
            .O(N__82824),
            .I(N__82798));
    Span4Mux_h I__19294 (
            .O(N__82821),
            .I(N__82798));
    InMux I__19293 (
            .O(N__82820),
            .I(N__82795));
    Span4Mux_v I__19292 (
            .O(N__82815),
            .I(N__82786));
    Span4Mux_v I__19291 (
            .O(N__82812),
            .I(N__82786));
    Span4Mux_h I__19290 (
            .O(N__82809),
            .I(N__82786));
    LocalMux I__19289 (
            .O(N__82804),
            .I(N__82786));
    InMux I__19288 (
            .O(N__82803),
            .I(N__82783));
    Odrv4 I__19287 (
            .O(N__82798),
            .I(\pid_side.error_6 ));
    LocalMux I__19286 (
            .O(N__82795),
            .I(\pid_side.error_6 ));
    Odrv4 I__19285 (
            .O(N__82786),
            .I(\pid_side.error_6 ));
    LocalMux I__19284 (
            .O(N__82783),
            .I(\pid_side.error_6 ));
    InMux I__19283 (
            .O(N__82774),
            .I(N__82768));
    InMux I__19282 (
            .O(N__82773),
            .I(N__82768));
    LocalMux I__19281 (
            .O(N__82768),
            .I(\pid_side.m58_0_o2_0 ));
    InMux I__19280 (
            .O(N__82765),
            .I(N__82760));
    InMux I__19279 (
            .O(N__82764),
            .I(N__82753));
    CascadeMux I__19278 (
            .O(N__82763),
            .I(N__82748));
    LocalMux I__19277 (
            .O(N__82760),
            .I(N__82745));
    InMux I__19276 (
            .O(N__82759),
            .I(N__82734));
    InMux I__19275 (
            .O(N__82758),
            .I(N__82731));
    InMux I__19274 (
            .O(N__82757),
            .I(N__82728));
    InMux I__19273 (
            .O(N__82756),
            .I(N__82725));
    LocalMux I__19272 (
            .O(N__82753),
            .I(N__82722));
    InMux I__19271 (
            .O(N__82752),
            .I(N__82719));
    InMux I__19270 (
            .O(N__82751),
            .I(N__82716));
    InMux I__19269 (
            .O(N__82748),
            .I(N__82713));
    Span4Mux_v I__19268 (
            .O(N__82745),
            .I(N__82710));
    InMux I__19267 (
            .O(N__82744),
            .I(N__82707));
    InMux I__19266 (
            .O(N__82743),
            .I(N__82702));
    InMux I__19265 (
            .O(N__82742),
            .I(N__82702));
    InMux I__19264 (
            .O(N__82741),
            .I(N__82697));
    InMux I__19263 (
            .O(N__82740),
            .I(N__82697));
    InMux I__19262 (
            .O(N__82739),
            .I(N__82690));
    InMux I__19261 (
            .O(N__82738),
            .I(N__82690));
    InMux I__19260 (
            .O(N__82737),
            .I(N__82690));
    LocalMux I__19259 (
            .O(N__82734),
            .I(N__82682));
    LocalMux I__19258 (
            .O(N__82731),
            .I(N__82679));
    LocalMux I__19257 (
            .O(N__82728),
            .I(N__82676));
    LocalMux I__19256 (
            .O(N__82725),
            .I(N__82671));
    Span4Mux_h I__19255 (
            .O(N__82722),
            .I(N__82671));
    LocalMux I__19254 (
            .O(N__82719),
            .I(N__82664));
    LocalMux I__19253 (
            .O(N__82716),
            .I(N__82664));
    LocalMux I__19252 (
            .O(N__82713),
            .I(N__82664));
    Span4Mux_h I__19251 (
            .O(N__82710),
            .I(N__82653));
    LocalMux I__19250 (
            .O(N__82707),
            .I(N__82653));
    LocalMux I__19249 (
            .O(N__82702),
            .I(N__82653));
    LocalMux I__19248 (
            .O(N__82697),
            .I(N__82653));
    LocalMux I__19247 (
            .O(N__82690),
            .I(N__82653));
    InMux I__19246 (
            .O(N__82689),
            .I(N__82650));
    InMux I__19245 (
            .O(N__82688),
            .I(N__82647));
    InMux I__19244 (
            .O(N__82687),
            .I(N__82644));
    InMux I__19243 (
            .O(N__82686),
            .I(N__82641));
    InMux I__19242 (
            .O(N__82685),
            .I(N__82632));
    Span4Mux_v I__19241 (
            .O(N__82682),
            .I(N__82627));
    Span4Mux_h I__19240 (
            .O(N__82679),
            .I(N__82627));
    Span4Mux_v I__19239 (
            .O(N__82676),
            .I(N__82620));
    Span4Mux_v I__19238 (
            .O(N__82671),
            .I(N__82620));
    Span4Mux_h I__19237 (
            .O(N__82664),
            .I(N__82620));
    Sp12to4 I__19236 (
            .O(N__82653),
            .I(N__82615));
    LocalMux I__19235 (
            .O(N__82650),
            .I(N__82615));
    LocalMux I__19234 (
            .O(N__82647),
            .I(N__82608));
    LocalMux I__19233 (
            .O(N__82644),
            .I(N__82608));
    LocalMux I__19232 (
            .O(N__82641),
            .I(N__82608));
    InMux I__19231 (
            .O(N__82640),
            .I(N__82605));
    InMux I__19230 (
            .O(N__82639),
            .I(N__82602));
    InMux I__19229 (
            .O(N__82638),
            .I(N__82597));
    InMux I__19228 (
            .O(N__82637),
            .I(N__82597));
    InMux I__19227 (
            .O(N__82636),
            .I(N__82594));
    InMux I__19226 (
            .O(N__82635),
            .I(N__82591));
    LocalMux I__19225 (
            .O(N__82632),
            .I(N__82586));
    Span4Mux_h I__19224 (
            .O(N__82627),
            .I(N__82586));
    Span4Mux_h I__19223 (
            .O(N__82620),
            .I(N__82583));
    Span12Mux_s9_h I__19222 (
            .O(N__82615),
            .I(N__82580));
    Span4Mux_v I__19221 (
            .O(N__82608),
            .I(N__82577));
    LocalMux I__19220 (
            .O(N__82605),
            .I(xy_ki_0_rep2));
    LocalMux I__19219 (
            .O(N__82602),
            .I(xy_ki_0_rep2));
    LocalMux I__19218 (
            .O(N__82597),
            .I(xy_ki_0_rep2));
    LocalMux I__19217 (
            .O(N__82594),
            .I(xy_ki_0_rep2));
    LocalMux I__19216 (
            .O(N__82591),
            .I(xy_ki_0_rep2));
    Odrv4 I__19215 (
            .O(N__82586),
            .I(xy_ki_0_rep2));
    Odrv4 I__19214 (
            .O(N__82583),
            .I(xy_ki_0_rep2));
    Odrv12 I__19213 (
            .O(N__82580),
            .I(xy_ki_0_rep2));
    Odrv4 I__19212 (
            .O(N__82577),
            .I(xy_ki_0_rep2));
    InMux I__19211 (
            .O(N__82558),
            .I(N__82555));
    LocalMux I__19210 (
            .O(N__82555),
            .I(N__82552));
    Span4Mux_h I__19209 (
            .O(N__82552),
            .I(N__82549));
    Odrv4 I__19208 (
            .O(N__82549),
            .I(\pid_side.O_2_8 ));
    InMux I__19207 (
            .O(N__82546),
            .I(N__82540));
    InMux I__19206 (
            .O(N__82545),
            .I(N__82540));
    LocalMux I__19205 (
            .O(N__82540),
            .I(N__82537));
    Odrv4 I__19204 (
            .O(N__82537),
            .I(\pid_side.error_p_regZ0Z_4 ));
    InMux I__19203 (
            .O(N__82534),
            .I(N__82528));
    InMux I__19202 (
            .O(N__82533),
            .I(N__82523));
    InMux I__19201 (
            .O(N__82532),
            .I(N__82523));
    InMux I__19200 (
            .O(N__82531),
            .I(N__82520));
    LocalMux I__19199 (
            .O(N__82528),
            .I(N__82517));
    LocalMux I__19198 (
            .O(N__82523),
            .I(N__82514));
    LocalMux I__19197 (
            .O(N__82520),
            .I(N__82511));
    Span4Mux_h I__19196 (
            .O(N__82517),
            .I(N__82508));
    Span4Mux_v I__19195 (
            .O(N__82514),
            .I(N__82503));
    Span4Mux_h I__19194 (
            .O(N__82511),
            .I(N__82503));
    Odrv4 I__19193 (
            .O(N__82508),
            .I(\pid_side.error_d_reg_prevZ0Z_1 ));
    Odrv4 I__19192 (
            .O(N__82503),
            .I(\pid_side.error_d_reg_prevZ0Z_1 ));
    InMux I__19191 (
            .O(N__82498),
            .I(N__82494));
    InMux I__19190 (
            .O(N__82497),
            .I(N__82491));
    LocalMux I__19189 (
            .O(N__82494),
            .I(N__82487));
    LocalMux I__19188 (
            .O(N__82491),
            .I(N__82484));
    InMux I__19187 (
            .O(N__82490),
            .I(N__82481));
    Span4Mux_v I__19186 (
            .O(N__82487),
            .I(N__82473));
    Span4Mux_h I__19185 (
            .O(N__82484),
            .I(N__82473));
    LocalMux I__19184 (
            .O(N__82481),
            .I(N__82470));
    InMux I__19183 (
            .O(N__82480),
            .I(N__82463));
    InMux I__19182 (
            .O(N__82479),
            .I(N__82463));
    InMux I__19181 (
            .O(N__82478),
            .I(N__82463));
    Odrv4 I__19180 (
            .O(N__82473),
            .I(\pid_side.error_d_regZ0Z_1 ));
    Odrv4 I__19179 (
            .O(N__82470),
            .I(\pid_side.error_d_regZ0Z_1 ));
    LocalMux I__19178 (
            .O(N__82463),
            .I(\pid_side.error_d_regZ0Z_1 ));
    InMux I__19177 (
            .O(N__82456),
            .I(N__82453));
    LocalMux I__19176 (
            .O(N__82453),
            .I(N__82450));
    Span4Mux_v I__19175 (
            .O(N__82450),
            .I(N__82447));
    Odrv4 I__19174 (
            .O(N__82447),
            .I(\pid_side.error_d_reg_prev_esr_RNIIFEIZ0Z_1 ));
    CascadeMux I__19173 (
            .O(N__82444),
            .I(N__82441));
    InMux I__19172 (
            .O(N__82441),
            .I(N__82435));
    InMux I__19171 (
            .O(N__82440),
            .I(N__82435));
    LocalMux I__19170 (
            .O(N__82435),
            .I(N__82432));
    Span4Mux_v I__19169 (
            .O(N__82432),
            .I(N__82429));
    Span4Mux_h I__19168 (
            .O(N__82429),
            .I(N__82426));
    Odrv4 I__19167 (
            .O(N__82426),
            .I(\pid_side.error_d_reg_prev_esr_RNIH7JOZ0Z_18 ));
    CascadeMux I__19166 (
            .O(N__82423),
            .I(N__82420));
    InMux I__19165 (
            .O(N__82420),
            .I(N__82414));
    InMux I__19164 (
            .O(N__82419),
            .I(N__82414));
    LocalMux I__19163 (
            .O(N__82414),
            .I(N__82411));
    Span4Mux_h I__19162 (
            .O(N__82411),
            .I(N__82408));
    Odrv4 I__19161 (
            .O(N__82408),
            .I(\pid_side.error_d_reg_prevZ0Z_19 ));
    InMux I__19160 (
            .O(N__82405),
            .I(N__82397));
    InMux I__19159 (
            .O(N__82404),
            .I(N__82397));
    InMux I__19158 (
            .O(N__82403),
            .I(N__82392));
    InMux I__19157 (
            .O(N__82402),
            .I(N__82392));
    LocalMux I__19156 (
            .O(N__82397),
            .I(N__82387));
    LocalMux I__19155 (
            .O(N__82392),
            .I(N__82387));
    Span4Mux_h I__19154 (
            .O(N__82387),
            .I(N__82384));
    Odrv4 I__19153 (
            .O(N__82384),
            .I(\pid_side.un1_pid_prereg_135_0 ));
    InMux I__19152 (
            .O(N__82381),
            .I(N__82378));
    LocalMux I__19151 (
            .O(N__82378),
            .I(N__82375));
    Odrv4 I__19150 (
            .O(N__82375),
            .I(\pid_side.g0_1_0 ));
    InMux I__19149 (
            .O(N__82372),
            .I(N__82365));
    InMux I__19148 (
            .O(N__82371),
            .I(N__82362));
    InMux I__19147 (
            .O(N__82370),
            .I(N__82355));
    InMux I__19146 (
            .O(N__82369),
            .I(N__82355));
    InMux I__19145 (
            .O(N__82368),
            .I(N__82355));
    LocalMux I__19144 (
            .O(N__82365),
            .I(N__82352));
    LocalMux I__19143 (
            .O(N__82362),
            .I(N__82345));
    LocalMux I__19142 (
            .O(N__82355),
            .I(N__82345));
    Span4Mux_h I__19141 (
            .O(N__82352),
            .I(N__82345));
    Odrv4 I__19140 (
            .O(N__82345),
            .I(\pid_side.error_d_reg_prevZ0Z_11 ));
    InMux I__19139 (
            .O(N__82342),
            .I(N__82336));
    InMux I__19138 (
            .O(N__82341),
            .I(N__82336));
    LocalMux I__19137 (
            .O(N__82336),
            .I(N__82333));
    Span4Mux_h I__19136 (
            .O(N__82333),
            .I(N__82330));
    Span4Mux_h I__19135 (
            .O(N__82330),
            .I(N__82327));
    Odrv4 I__19134 (
            .O(N__82327),
            .I(\pid_side.error_d_reg_prev_esr_RNISHIO_1Z0Z_11 ));
    InMux I__19133 (
            .O(N__82324),
            .I(N__82321));
    LocalMux I__19132 (
            .O(N__82321),
            .I(N__82318));
    Span4Mux_v I__19131 (
            .O(N__82318),
            .I(N__82314));
    InMux I__19130 (
            .O(N__82317),
            .I(N__82311));
    Span4Mux_h I__19129 (
            .O(N__82314),
            .I(N__82308));
    LocalMux I__19128 (
            .O(N__82311),
            .I(N__82305));
    Span4Mux_h I__19127 (
            .O(N__82308),
            .I(N__82302));
    Odrv4 I__19126 (
            .O(N__82305),
            .I(\pid_side.error_d_reg_fastZ0Z_13 ));
    Odrv4 I__19125 (
            .O(N__82302),
            .I(\pid_side.error_d_reg_fastZ0Z_13 ));
    InMux I__19124 (
            .O(N__82297),
            .I(N__82293));
    InMux I__19123 (
            .O(N__82296),
            .I(N__82290));
    LocalMux I__19122 (
            .O(N__82293),
            .I(N__82285));
    LocalMux I__19121 (
            .O(N__82290),
            .I(N__82285));
    Span4Mux_h I__19120 (
            .O(N__82285),
            .I(N__82282));
    Odrv4 I__19119 (
            .O(N__82282),
            .I(\pid_front.m0_0_03 ));
    InMux I__19118 (
            .O(N__82279),
            .I(N__82271));
    InMux I__19117 (
            .O(N__82278),
            .I(N__82271));
    InMux I__19116 (
            .O(N__82277),
            .I(N__82266));
    InMux I__19115 (
            .O(N__82276),
            .I(N__82266));
    LocalMux I__19114 (
            .O(N__82271),
            .I(N__82260));
    LocalMux I__19113 (
            .O(N__82266),
            .I(N__82260));
    InMux I__19112 (
            .O(N__82265),
            .I(N__82249));
    Span4Mux_v I__19111 (
            .O(N__82260),
            .I(N__82246));
    InMux I__19110 (
            .O(N__82259),
            .I(N__82241));
    InMux I__19109 (
            .O(N__82258),
            .I(N__82241));
    InMux I__19108 (
            .O(N__82257),
            .I(N__82237));
    InMux I__19107 (
            .O(N__82256),
            .I(N__82230));
    InMux I__19106 (
            .O(N__82255),
            .I(N__82230));
    InMux I__19105 (
            .O(N__82254),
            .I(N__82230));
    InMux I__19104 (
            .O(N__82253),
            .I(N__82227));
    InMux I__19103 (
            .O(N__82252),
            .I(N__82224));
    LocalMux I__19102 (
            .O(N__82249),
            .I(N__82217));
    Span4Mux_v I__19101 (
            .O(N__82246),
            .I(N__82217));
    LocalMux I__19100 (
            .O(N__82241),
            .I(N__82217));
    InMux I__19099 (
            .O(N__82240),
            .I(N__82213));
    LocalMux I__19098 (
            .O(N__82237),
            .I(N__82208));
    LocalMux I__19097 (
            .O(N__82230),
            .I(N__82205));
    LocalMux I__19096 (
            .O(N__82227),
            .I(N__82202));
    LocalMux I__19095 (
            .O(N__82224),
            .I(N__82197));
    Span4Mux_h I__19094 (
            .O(N__82217),
            .I(N__82197));
    InMux I__19093 (
            .O(N__82216),
            .I(N__82194));
    LocalMux I__19092 (
            .O(N__82213),
            .I(N__82191));
    InMux I__19091 (
            .O(N__82212),
            .I(N__82188));
    InMux I__19090 (
            .O(N__82211),
            .I(N__82183));
    Span12Mux_h I__19089 (
            .O(N__82208),
            .I(N__82180));
    Span12Mux_h I__19088 (
            .O(N__82205),
            .I(N__82177));
    Span4Mux_h I__19087 (
            .O(N__82202),
            .I(N__82170));
    Span4Mux_h I__19086 (
            .O(N__82197),
            .I(N__82170));
    LocalMux I__19085 (
            .O(N__82194),
            .I(N__82170));
    Span4Mux_h I__19084 (
            .O(N__82191),
            .I(N__82165));
    LocalMux I__19083 (
            .O(N__82188),
            .I(N__82165));
    InMux I__19082 (
            .O(N__82187),
            .I(N__82160));
    InMux I__19081 (
            .O(N__82186),
            .I(N__82160));
    LocalMux I__19080 (
            .O(N__82183),
            .I(xy_ki_fast_0));
    Odrv12 I__19079 (
            .O(N__82180),
            .I(xy_ki_fast_0));
    Odrv12 I__19078 (
            .O(N__82177),
            .I(xy_ki_fast_0));
    Odrv4 I__19077 (
            .O(N__82170),
            .I(xy_ki_fast_0));
    Odrv4 I__19076 (
            .O(N__82165),
            .I(xy_ki_fast_0));
    LocalMux I__19075 (
            .O(N__82160),
            .I(xy_ki_fast_0));
    InMux I__19074 (
            .O(N__82147),
            .I(N__82144));
    LocalMux I__19073 (
            .O(N__82144),
            .I(N__82141));
    Odrv4 I__19072 (
            .O(N__82141),
            .I(\pid_front.N_574 ));
    InMux I__19071 (
            .O(N__82138),
            .I(N__82135));
    LocalMux I__19070 (
            .O(N__82135),
            .I(N__82132));
    Span4Mux_v I__19069 (
            .O(N__82132),
            .I(N__82126));
    InMux I__19068 (
            .O(N__82131),
            .I(N__82123));
    InMux I__19067 (
            .O(N__82130),
            .I(N__82120));
    InMux I__19066 (
            .O(N__82129),
            .I(N__82117));
    Span4Mux_h I__19065 (
            .O(N__82126),
            .I(N__82112));
    LocalMux I__19064 (
            .O(N__82123),
            .I(N__82112));
    LocalMux I__19063 (
            .O(N__82120),
            .I(N__82109));
    LocalMux I__19062 (
            .O(N__82117),
            .I(N__82106));
    Span4Mux_v I__19061 (
            .O(N__82112),
            .I(N__82103));
    Span4Mux_v I__19060 (
            .O(N__82109),
            .I(N__82098));
    Span4Mux_h I__19059 (
            .O(N__82106),
            .I(N__82098));
    Span4Mux_h I__19058 (
            .O(N__82103),
            .I(N__82095));
    Span4Mux_v I__19057 (
            .O(N__82098),
            .I(N__82092));
    Odrv4 I__19056 (
            .O(N__82095),
            .I(\pid_front.state_ns_0 ));
    Odrv4 I__19055 (
            .O(N__82092),
            .I(\pid_front.state_ns_0 ));
    InMux I__19054 (
            .O(N__82087),
            .I(N__82083));
    InMux I__19053 (
            .O(N__82086),
            .I(N__82079));
    LocalMux I__19052 (
            .O(N__82083),
            .I(N__82074));
    InMux I__19051 (
            .O(N__82082),
            .I(N__82071));
    LocalMux I__19050 (
            .O(N__82079),
            .I(N__82068));
    InMux I__19049 (
            .O(N__82078),
            .I(N__82065));
    InMux I__19048 (
            .O(N__82077),
            .I(N__82061));
    Span4Mux_v I__19047 (
            .O(N__82074),
            .I(N__82058));
    LocalMux I__19046 (
            .O(N__82071),
            .I(N__82055));
    Span4Mux_h I__19045 (
            .O(N__82068),
            .I(N__82052));
    LocalMux I__19044 (
            .O(N__82065),
            .I(N__82048));
    CascadeMux I__19043 (
            .O(N__82064),
            .I(N__82045));
    LocalMux I__19042 (
            .O(N__82061),
            .I(N__82042));
    Span4Mux_h I__19041 (
            .O(N__82058),
            .I(N__82037));
    Span4Mux_h I__19040 (
            .O(N__82055),
            .I(N__82037));
    Span4Mux_v I__19039 (
            .O(N__82052),
            .I(N__82034));
    CascadeMux I__19038 (
            .O(N__82051),
            .I(N__82031));
    Span4Mux_h I__19037 (
            .O(N__82048),
            .I(N__82028));
    InMux I__19036 (
            .O(N__82045),
            .I(N__82025));
    Span4Mux_v I__19035 (
            .O(N__82042),
            .I(N__82022));
    Span4Mux_v I__19034 (
            .O(N__82037),
            .I(N__82017));
    Span4Mux_v I__19033 (
            .O(N__82034),
            .I(N__82017));
    InMux I__19032 (
            .O(N__82031),
            .I(N__82014));
    Sp12to4 I__19031 (
            .O(N__82028),
            .I(N__82011));
    LocalMux I__19030 (
            .O(N__82025),
            .I(N__82004));
    Span4Mux_h I__19029 (
            .O(N__82022),
            .I(N__82004));
    Span4Mux_h I__19028 (
            .O(N__82017),
            .I(N__82004));
    LocalMux I__19027 (
            .O(N__82014),
            .I(pid_side_N_607));
    Odrv12 I__19026 (
            .O(N__82011),
            .I(pid_side_N_607));
    Odrv4 I__19025 (
            .O(N__82004),
            .I(pid_side_N_607));
    InMux I__19024 (
            .O(N__81997),
            .I(N__81994));
    LocalMux I__19023 (
            .O(N__81994),
            .I(\pid_front.m7_2_01 ));
    InMux I__19022 (
            .O(N__81991),
            .I(N__81987));
    CascadeMux I__19021 (
            .O(N__81990),
            .I(N__81984));
    LocalMux I__19020 (
            .O(N__81987),
            .I(N__81981));
    InMux I__19019 (
            .O(N__81984),
            .I(N__81978));
    Span4Mux_h I__19018 (
            .O(N__81981),
            .I(N__81975));
    LocalMux I__19017 (
            .O(N__81978),
            .I(\pid_front.error_i_regZ0Z_3 ));
    Odrv4 I__19016 (
            .O(N__81975),
            .I(\pid_front.error_i_regZ0Z_3 ));
    InMux I__19015 (
            .O(N__81970),
            .I(N__81967));
    LocalMux I__19014 (
            .O(N__81967),
            .I(N__81964));
    Span4Mux_v I__19013 (
            .O(N__81964),
            .I(N__81961));
    Odrv4 I__19012 (
            .O(N__81961),
            .I(\pid_front.O_21 ));
    InMux I__19011 (
            .O(N__81958),
            .I(N__81953));
    InMux I__19010 (
            .O(N__81957),
            .I(N__81948));
    InMux I__19009 (
            .O(N__81956),
            .I(N__81948));
    LocalMux I__19008 (
            .O(N__81953),
            .I(N__81945));
    LocalMux I__19007 (
            .O(N__81948),
            .I(N__81942));
    Span4Mux_v I__19006 (
            .O(N__81945),
            .I(N__81937));
    Span4Mux_h I__19005 (
            .O(N__81942),
            .I(N__81937));
    Odrv4 I__19004 (
            .O(N__81937),
            .I(\pid_front.error_d_regZ0Z_18 ));
    InMux I__19003 (
            .O(N__81934),
            .I(N__81931));
    LocalMux I__19002 (
            .O(N__81931),
            .I(N__81928));
    Odrv12 I__19001 (
            .O(N__81928),
            .I(\pid_front.O_5 ));
    InMux I__19000 (
            .O(N__81925),
            .I(N__81916));
    InMux I__18999 (
            .O(N__81924),
            .I(N__81916));
    InMux I__18998 (
            .O(N__81923),
            .I(N__81916));
    LocalMux I__18997 (
            .O(N__81916),
            .I(N__81913));
    Span4Mux_h I__18996 (
            .O(N__81913),
            .I(N__81910));
    Odrv4 I__18995 (
            .O(N__81910),
            .I(\pid_front.error_d_regZ0Z_2 ));
    InMux I__18994 (
            .O(N__81907),
            .I(N__81904));
    LocalMux I__18993 (
            .O(N__81904),
            .I(N__81901));
    Odrv12 I__18992 (
            .O(N__81901),
            .I(\pid_front.O_13 ));
    CascadeMux I__18991 (
            .O(N__81898),
            .I(N__81891));
    InMux I__18990 (
            .O(N__81897),
            .I(N__81885));
    InMux I__18989 (
            .O(N__81896),
            .I(N__81885));
    InMux I__18988 (
            .O(N__81895),
            .I(N__81876));
    InMux I__18987 (
            .O(N__81894),
            .I(N__81876));
    InMux I__18986 (
            .O(N__81891),
            .I(N__81876));
    InMux I__18985 (
            .O(N__81890),
            .I(N__81876));
    LocalMux I__18984 (
            .O(N__81885),
            .I(N__81873));
    LocalMux I__18983 (
            .O(N__81876),
            .I(N__81870));
    Span4Mux_h I__18982 (
            .O(N__81873),
            .I(N__81867));
    Span4Mux_h I__18981 (
            .O(N__81870),
            .I(N__81864));
    Odrv4 I__18980 (
            .O(N__81867),
            .I(\pid_front.error_d_regZ0Z_10 ));
    Odrv4 I__18979 (
            .O(N__81864),
            .I(\pid_front.error_d_regZ0Z_10 ));
    InMux I__18978 (
            .O(N__81859),
            .I(N__81856));
    LocalMux I__18977 (
            .O(N__81856),
            .I(N__81853));
    Span4Mux_v I__18976 (
            .O(N__81853),
            .I(N__81849));
    InMux I__18975 (
            .O(N__81852),
            .I(N__81846));
    Span4Mux_h I__18974 (
            .O(N__81849),
            .I(N__81841));
    LocalMux I__18973 (
            .O(N__81846),
            .I(N__81841));
    Span4Mux_h I__18972 (
            .O(N__81841),
            .I(N__81838));
    Odrv4 I__18971 (
            .O(N__81838),
            .I(\pid_front.O_15 ));
    InMux I__18970 (
            .O(N__81835),
            .I(N__81828));
    InMux I__18969 (
            .O(N__81834),
            .I(N__81828));
    InMux I__18968 (
            .O(N__81833),
            .I(N__81820));
    LocalMux I__18967 (
            .O(N__81828),
            .I(N__81816));
    InMux I__18966 (
            .O(N__81827),
            .I(N__81811));
    InMux I__18965 (
            .O(N__81826),
            .I(N__81811));
    InMux I__18964 (
            .O(N__81825),
            .I(N__81804));
    InMux I__18963 (
            .O(N__81824),
            .I(N__81804));
    InMux I__18962 (
            .O(N__81823),
            .I(N__81804));
    LocalMux I__18961 (
            .O(N__81820),
            .I(N__81801));
    InMux I__18960 (
            .O(N__81819),
            .I(N__81798));
    Span4Mux_v I__18959 (
            .O(N__81816),
            .I(N__81793));
    LocalMux I__18958 (
            .O(N__81811),
            .I(N__81793));
    LocalMux I__18957 (
            .O(N__81804),
            .I(N__81790));
    Span4Mux_h I__18956 (
            .O(N__81801),
            .I(N__81787));
    LocalMux I__18955 (
            .O(N__81798),
            .I(N__81784));
    Span4Mux_v I__18954 (
            .O(N__81793),
            .I(N__81779));
    Span4Mux_h I__18953 (
            .O(N__81790),
            .I(N__81779));
    Span4Mux_h I__18952 (
            .O(N__81787),
            .I(N__81776));
    Span4Mux_v I__18951 (
            .O(N__81784),
            .I(N__81771));
    Span4Mux_h I__18950 (
            .O(N__81779),
            .I(N__81771));
    Odrv4 I__18949 (
            .O(N__81776),
            .I(\pid_front.error_d_regZ0Z_12 ));
    Odrv4 I__18948 (
            .O(N__81771),
            .I(\pid_front.error_d_regZ0Z_12 ));
    InMux I__18947 (
            .O(N__81766),
            .I(N__81763));
    LocalMux I__18946 (
            .O(N__81763),
            .I(N__81760));
    Span4Mux_v I__18945 (
            .O(N__81760),
            .I(N__81757));
    Span4Mux_h I__18944 (
            .O(N__81757),
            .I(N__81754));
    Odrv4 I__18943 (
            .O(N__81754),
            .I(\pid_front.O_9 ));
    InMux I__18942 (
            .O(N__81751),
            .I(N__81748));
    LocalMux I__18941 (
            .O(N__81748),
            .I(N__81745));
    Span4Mux_h I__18940 (
            .O(N__81745),
            .I(N__81739));
    InMux I__18939 (
            .O(N__81744),
            .I(N__81732));
    InMux I__18938 (
            .O(N__81743),
            .I(N__81732));
    InMux I__18937 (
            .O(N__81742),
            .I(N__81732));
    Span4Mux_v I__18936 (
            .O(N__81739),
            .I(N__81727));
    LocalMux I__18935 (
            .O(N__81732),
            .I(N__81727));
    Span4Mux_h I__18934 (
            .O(N__81727),
            .I(N__81722));
    InMux I__18933 (
            .O(N__81726),
            .I(N__81719));
    InMux I__18932 (
            .O(N__81725),
            .I(N__81716));
    Span4Mux_h I__18931 (
            .O(N__81722),
            .I(N__81713));
    LocalMux I__18930 (
            .O(N__81719),
            .I(N__81708));
    LocalMux I__18929 (
            .O(N__81716),
            .I(N__81708));
    Odrv4 I__18928 (
            .O(N__81713),
            .I(\pid_front.error_d_regZ0Z_6 ));
    Odrv12 I__18927 (
            .O(N__81708),
            .I(\pid_front.error_d_regZ0Z_6 ));
    InMux I__18926 (
            .O(N__81703),
            .I(N__81700));
    LocalMux I__18925 (
            .O(N__81700),
            .I(N__81697));
    Span4Mux_h I__18924 (
            .O(N__81697),
            .I(N__81694));
    Span4Mux_v I__18923 (
            .O(N__81694),
            .I(N__81691));
    Odrv4 I__18922 (
            .O(N__81691),
            .I(\pid_side.O_1_11 ));
    InMux I__18921 (
            .O(N__81688),
            .I(N__81685));
    LocalMux I__18920 (
            .O(N__81685),
            .I(N__81679));
    InMux I__18919 (
            .O(N__81684),
            .I(N__81674));
    InMux I__18918 (
            .O(N__81683),
            .I(N__81674));
    InMux I__18917 (
            .O(N__81682),
            .I(N__81671));
    Span4Mux_v I__18916 (
            .O(N__81679),
            .I(N__81666));
    LocalMux I__18915 (
            .O(N__81674),
            .I(N__81666));
    LocalMux I__18914 (
            .O(N__81671),
            .I(N__81663));
    Span4Mux_h I__18913 (
            .O(N__81666),
            .I(N__81660));
    Odrv12 I__18912 (
            .O(N__81663),
            .I(\pid_side.error_d_regZ0Z_8 ));
    Odrv4 I__18911 (
            .O(N__81660),
            .I(\pid_side.error_d_regZ0Z_8 ));
    InMux I__18910 (
            .O(N__81655),
            .I(N__81650));
    InMux I__18909 (
            .O(N__81654),
            .I(N__81644));
    InMux I__18908 (
            .O(N__81653),
            .I(N__81641));
    LocalMux I__18907 (
            .O(N__81650),
            .I(N__81637));
    InMux I__18906 (
            .O(N__81649),
            .I(N__81634));
    InMux I__18905 (
            .O(N__81648),
            .I(N__81631));
    InMux I__18904 (
            .O(N__81647),
            .I(N__81627));
    LocalMux I__18903 (
            .O(N__81644),
            .I(N__81624));
    LocalMux I__18902 (
            .O(N__81641),
            .I(N__81621));
    InMux I__18901 (
            .O(N__81640),
            .I(N__81618));
    Span4Mux_v I__18900 (
            .O(N__81637),
            .I(N__81615));
    LocalMux I__18899 (
            .O(N__81634),
            .I(N__81612));
    LocalMux I__18898 (
            .O(N__81631),
            .I(N__81609));
    InMux I__18897 (
            .O(N__81630),
            .I(N__81606));
    LocalMux I__18896 (
            .O(N__81627),
            .I(N__81603));
    Span4Mux_h I__18895 (
            .O(N__81624),
            .I(N__81599));
    Span4Mux_v I__18894 (
            .O(N__81621),
            .I(N__81594));
    LocalMux I__18893 (
            .O(N__81618),
            .I(N__81594));
    Span4Mux_v I__18892 (
            .O(N__81615),
            .I(N__81589));
    Span4Mux_s0_h I__18891 (
            .O(N__81612),
            .I(N__81589));
    Span4Mux_v I__18890 (
            .O(N__81609),
            .I(N__81584));
    LocalMux I__18889 (
            .O(N__81606),
            .I(N__81584));
    Span4Mux_h I__18888 (
            .O(N__81603),
            .I(N__81581));
    CascadeMux I__18887 (
            .O(N__81602),
            .I(N__81578));
    Span4Mux_v I__18886 (
            .O(N__81599),
            .I(N__81569));
    Span4Mux_h I__18885 (
            .O(N__81594),
            .I(N__81569));
    Span4Mux_h I__18884 (
            .O(N__81589),
            .I(N__81564));
    Span4Mux_h I__18883 (
            .O(N__81584),
            .I(N__81564));
    Span4Mux_h I__18882 (
            .O(N__81581),
            .I(N__81561));
    InMux I__18881 (
            .O(N__81578),
            .I(N__81556));
    InMux I__18880 (
            .O(N__81577),
            .I(N__81556));
    InMux I__18879 (
            .O(N__81576),
            .I(N__81553));
    InMux I__18878 (
            .O(N__81575),
            .I(N__81548));
    InMux I__18877 (
            .O(N__81574),
            .I(N__81548));
    Odrv4 I__18876 (
            .O(N__81569),
            .I(\pid_side.error_14 ));
    Odrv4 I__18875 (
            .O(N__81564),
            .I(\pid_side.error_14 ));
    Odrv4 I__18874 (
            .O(N__81561),
            .I(\pid_side.error_14 ));
    LocalMux I__18873 (
            .O(N__81556),
            .I(\pid_side.error_14 ));
    LocalMux I__18872 (
            .O(N__81553),
            .I(\pid_side.error_14 ));
    LocalMux I__18871 (
            .O(N__81548),
            .I(\pid_side.error_14 ));
    InMux I__18870 (
            .O(N__81535),
            .I(N__81530));
    InMux I__18869 (
            .O(N__81534),
            .I(N__81527));
    InMux I__18868 (
            .O(N__81533),
            .I(N__81521));
    LocalMux I__18867 (
            .O(N__81530),
            .I(N__81517));
    LocalMux I__18866 (
            .O(N__81527),
            .I(N__81514));
    InMux I__18865 (
            .O(N__81526),
            .I(N__81511));
    InMux I__18864 (
            .O(N__81525),
            .I(N__81506));
    InMux I__18863 (
            .O(N__81524),
            .I(N__81506));
    LocalMux I__18862 (
            .O(N__81521),
            .I(N__81503));
    InMux I__18861 (
            .O(N__81520),
            .I(N__81500));
    Span4Mux_s0_h I__18860 (
            .O(N__81517),
            .I(N__81496));
    Span4Mux_v I__18859 (
            .O(N__81514),
            .I(N__81493));
    LocalMux I__18858 (
            .O(N__81511),
            .I(N__81488));
    LocalMux I__18857 (
            .O(N__81506),
            .I(N__81488));
    Span4Mux_s1_h I__18856 (
            .O(N__81503),
            .I(N__81484));
    LocalMux I__18855 (
            .O(N__81500),
            .I(N__81481));
    InMux I__18854 (
            .O(N__81499),
            .I(N__81478));
    Span4Mux_h I__18853 (
            .O(N__81496),
            .I(N__81475));
    Span4Mux_h I__18852 (
            .O(N__81493),
            .I(N__81472));
    Span4Mux_h I__18851 (
            .O(N__81488),
            .I(N__81469));
    InMux I__18850 (
            .O(N__81487),
            .I(N__81466));
    Span4Mux_h I__18849 (
            .O(N__81484),
            .I(N__81459));
    Span4Mux_v I__18848 (
            .O(N__81481),
            .I(N__81459));
    LocalMux I__18847 (
            .O(N__81478),
            .I(N__81459));
    Odrv4 I__18846 (
            .O(N__81475),
            .I(\pid_side.error_10 ));
    Odrv4 I__18845 (
            .O(N__81472),
            .I(\pid_side.error_10 ));
    Odrv4 I__18844 (
            .O(N__81469),
            .I(\pid_side.error_10 ));
    LocalMux I__18843 (
            .O(N__81466),
            .I(\pid_side.error_10 ));
    Odrv4 I__18842 (
            .O(N__81459),
            .I(\pid_side.error_10 ));
    CascadeMux I__18841 (
            .O(N__81448),
            .I(\pid_side.N_225_cascade_ ));
    InMux I__18840 (
            .O(N__81445),
            .I(N__81438));
    InMux I__18839 (
            .O(N__81444),
            .I(N__81435));
    InMux I__18838 (
            .O(N__81443),
            .I(N__81432));
    InMux I__18837 (
            .O(N__81442),
            .I(N__81429));
    InMux I__18836 (
            .O(N__81441),
            .I(N__81426));
    LocalMux I__18835 (
            .O(N__81438),
            .I(N__81420));
    LocalMux I__18834 (
            .O(N__81435),
            .I(N__81420));
    LocalMux I__18833 (
            .O(N__81432),
            .I(N__81416));
    LocalMux I__18832 (
            .O(N__81429),
            .I(N__81411));
    LocalMux I__18831 (
            .O(N__81426),
            .I(N__81411));
    InMux I__18830 (
            .O(N__81425),
            .I(N__81408));
    Span4Mux_h I__18829 (
            .O(N__81420),
            .I(N__81405));
    InMux I__18828 (
            .O(N__81419),
            .I(N__81400));
    Span4Mux_v I__18827 (
            .O(N__81416),
            .I(N__81395));
    Span4Mux_v I__18826 (
            .O(N__81411),
            .I(N__81395));
    LocalMux I__18825 (
            .O(N__81408),
            .I(N__81390));
    Span4Mux_v I__18824 (
            .O(N__81405),
            .I(N__81390));
    InMux I__18823 (
            .O(N__81404),
            .I(N__81387));
    InMux I__18822 (
            .O(N__81403),
            .I(N__81384));
    LocalMux I__18821 (
            .O(N__81400),
            .I(pid_side_N_174));
    Odrv4 I__18820 (
            .O(N__81395),
            .I(pid_side_N_174));
    Odrv4 I__18819 (
            .O(N__81390),
            .I(pid_side_N_174));
    LocalMux I__18818 (
            .O(N__81387),
            .I(pid_side_N_174));
    LocalMux I__18817 (
            .O(N__81384),
            .I(pid_side_N_174));
    CascadeMux I__18816 (
            .O(N__81373),
            .I(\pid_side.m25_2_03_0_2_cascade_ ));
    InMux I__18815 (
            .O(N__81370),
            .I(N__81367));
    LocalMux I__18814 (
            .O(N__81367),
            .I(\pid_side.un4_error_i_reg_31_am_1 ));
    CascadeMux I__18813 (
            .O(N__81364),
            .I(\pid_side.error_i_reg_esr_RNO_0_0_21_cascade_ ));
    InMux I__18812 (
            .O(N__81361),
            .I(N__81358));
    LocalMux I__18811 (
            .O(N__81358),
            .I(\pid_side.error_i_reg_esr_RNO_1Z0Z_21 ));
    InMux I__18810 (
            .O(N__81355),
            .I(N__81352));
    LocalMux I__18809 (
            .O(N__81352),
            .I(N__81349));
    Span4Mux_v I__18808 (
            .O(N__81349),
            .I(N__81346));
    Span4Mux_v I__18807 (
            .O(N__81346),
            .I(N__81343));
    Span4Mux_h I__18806 (
            .O(N__81343),
            .I(N__81340));
    Odrv4 I__18805 (
            .O(N__81340),
            .I(\pid_side.error_i_regZ0Z_21 ));
    CascadeMux I__18804 (
            .O(N__81337),
            .I(\pid_side.N_254_cascade_ ));
    InMux I__18803 (
            .O(N__81334),
            .I(N__81329));
    InMux I__18802 (
            .O(N__81333),
            .I(N__81319));
    InMux I__18801 (
            .O(N__81332),
            .I(N__81315));
    LocalMux I__18800 (
            .O(N__81329),
            .I(N__81306));
    InMux I__18799 (
            .O(N__81328),
            .I(N__81301));
    InMux I__18798 (
            .O(N__81327),
            .I(N__81301));
    InMux I__18797 (
            .O(N__81326),
            .I(N__81298));
    InMux I__18796 (
            .O(N__81325),
            .I(N__81293));
    InMux I__18795 (
            .O(N__81324),
            .I(N__81293));
    InMux I__18794 (
            .O(N__81323),
            .I(N__81287));
    InMux I__18793 (
            .O(N__81322),
            .I(N__81287));
    LocalMux I__18792 (
            .O(N__81319),
            .I(N__81283));
    InMux I__18791 (
            .O(N__81318),
            .I(N__81280));
    LocalMux I__18790 (
            .O(N__81315),
            .I(N__81277));
    InMux I__18789 (
            .O(N__81314),
            .I(N__81274));
    InMux I__18788 (
            .O(N__81313),
            .I(N__81269));
    InMux I__18787 (
            .O(N__81312),
            .I(N__81269));
    InMux I__18786 (
            .O(N__81311),
            .I(N__81264));
    InMux I__18785 (
            .O(N__81310),
            .I(N__81264));
    InMux I__18784 (
            .O(N__81309),
            .I(N__81261));
    Span4Mux_v I__18783 (
            .O(N__81306),
            .I(N__81256));
    LocalMux I__18782 (
            .O(N__81301),
            .I(N__81253));
    LocalMux I__18781 (
            .O(N__81298),
            .I(N__81248));
    LocalMux I__18780 (
            .O(N__81293),
            .I(N__81248));
    InMux I__18779 (
            .O(N__81292),
            .I(N__81245));
    LocalMux I__18778 (
            .O(N__81287),
            .I(N__81240));
    InMux I__18777 (
            .O(N__81286),
            .I(N__81237));
    Span4Mux_h I__18776 (
            .O(N__81283),
            .I(N__81228));
    LocalMux I__18775 (
            .O(N__81280),
            .I(N__81228));
    Span4Mux_v I__18774 (
            .O(N__81277),
            .I(N__81228));
    LocalMux I__18773 (
            .O(N__81274),
            .I(N__81228));
    LocalMux I__18772 (
            .O(N__81269),
            .I(N__81221));
    LocalMux I__18771 (
            .O(N__81264),
            .I(N__81221));
    LocalMux I__18770 (
            .O(N__81261),
            .I(N__81221));
    InMux I__18769 (
            .O(N__81260),
            .I(N__81218));
    InMux I__18768 (
            .O(N__81259),
            .I(N__81215));
    Span4Mux_h I__18767 (
            .O(N__81256),
            .I(N__81212));
    Span4Mux_v I__18766 (
            .O(N__81253),
            .I(N__81205));
    Span4Mux_v I__18765 (
            .O(N__81248),
            .I(N__81205));
    LocalMux I__18764 (
            .O(N__81245),
            .I(N__81205));
    InMux I__18763 (
            .O(N__81244),
            .I(N__81202));
    InMux I__18762 (
            .O(N__81243),
            .I(N__81198));
    Span4Mux_h I__18761 (
            .O(N__81240),
            .I(N__81195));
    LocalMux I__18760 (
            .O(N__81237),
            .I(N__81188));
    Span4Mux_v I__18759 (
            .O(N__81228),
            .I(N__81188));
    Span4Mux_h I__18758 (
            .O(N__81221),
            .I(N__81188));
    LocalMux I__18757 (
            .O(N__81218),
            .I(N__81184));
    LocalMux I__18756 (
            .O(N__81215),
            .I(N__81175));
    Span4Mux_h I__18755 (
            .O(N__81212),
            .I(N__81175));
    Span4Mux_h I__18754 (
            .O(N__81205),
            .I(N__81175));
    LocalMux I__18753 (
            .O(N__81202),
            .I(N__81175));
    InMux I__18752 (
            .O(N__81201),
            .I(N__81172));
    LocalMux I__18751 (
            .O(N__81198),
            .I(N__81165));
    Span4Mux_h I__18750 (
            .O(N__81195),
            .I(N__81165));
    Span4Mux_h I__18749 (
            .O(N__81188),
            .I(N__81165));
    InMux I__18748 (
            .O(N__81187),
            .I(N__81162));
    Span4Mux_v I__18747 (
            .O(N__81184),
            .I(N__81157));
    Span4Mux_v I__18746 (
            .O(N__81175),
            .I(N__81157));
    LocalMux I__18745 (
            .O(N__81172),
            .I(N__81152));
    Sp12to4 I__18744 (
            .O(N__81165),
            .I(N__81152));
    LocalMux I__18743 (
            .O(N__81162),
            .I(pid_side_N_491));
    Odrv4 I__18742 (
            .O(N__81157),
            .I(pid_side_N_491));
    Odrv12 I__18741 (
            .O(N__81152),
            .I(pid_side_N_491));
    InMux I__18740 (
            .O(N__81145),
            .I(N__81142));
    LocalMux I__18739 (
            .O(N__81142),
            .I(N__81139));
    Span4Mux_h I__18738 (
            .O(N__81139),
            .I(N__81136));
    Span4Mux_h I__18737 (
            .O(N__81136),
            .I(N__81133));
    Odrv4 I__18736 (
            .O(N__81133),
            .I(\pid_side.m20_2_03_0_0 ));
    InMux I__18735 (
            .O(N__81130),
            .I(N__81127));
    LocalMux I__18734 (
            .O(N__81127),
            .I(N__81123));
    InMux I__18733 (
            .O(N__81126),
            .I(N__81120));
    Span4Mux_v I__18732 (
            .O(N__81123),
            .I(N__81117));
    LocalMux I__18731 (
            .O(N__81120),
            .I(pid_side_m20_2_03_0_a2_0_0));
    Odrv4 I__18730 (
            .O(N__81117),
            .I(pid_side_m20_2_03_0_a2_0_0));
    InMux I__18729 (
            .O(N__81112),
            .I(N__81107));
    InMux I__18728 (
            .O(N__81111),
            .I(N__81104));
    InMux I__18727 (
            .O(N__81110),
            .I(N__81100));
    LocalMux I__18726 (
            .O(N__81107),
            .I(N__81094));
    LocalMux I__18725 (
            .O(N__81104),
            .I(N__81091));
    InMux I__18724 (
            .O(N__81103),
            .I(N__81088));
    LocalMux I__18723 (
            .O(N__81100),
            .I(N__81085));
    InMux I__18722 (
            .O(N__81099),
            .I(N__81082));
    InMux I__18721 (
            .O(N__81098),
            .I(N__81076));
    InMux I__18720 (
            .O(N__81097),
            .I(N__81076));
    Span4Mux_h I__18719 (
            .O(N__81094),
            .I(N__81073));
    Span4Mux_h I__18718 (
            .O(N__81091),
            .I(N__81068));
    LocalMux I__18717 (
            .O(N__81088),
            .I(N__81068));
    Span4Mux_s0_h I__18716 (
            .O(N__81085),
            .I(N__81064));
    LocalMux I__18715 (
            .O(N__81082),
            .I(N__81061));
    CascadeMux I__18714 (
            .O(N__81081),
            .I(N__81058));
    LocalMux I__18713 (
            .O(N__81076),
            .I(N__81055));
    Span4Mux_h I__18712 (
            .O(N__81073),
            .I(N__81050));
    Span4Mux_h I__18711 (
            .O(N__81068),
            .I(N__81050));
    InMux I__18710 (
            .O(N__81067),
            .I(N__81047));
    Span4Mux_h I__18709 (
            .O(N__81064),
            .I(N__81044));
    Span12Mux_s5_h I__18708 (
            .O(N__81061),
            .I(N__81041));
    InMux I__18707 (
            .O(N__81058),
            .I(N__81038));
    Odrv12 I__18706 (
            .O(N__81055),
            .I(\pid_side.error_2 ));
    Odrv4 I__18705 (
            .O(N__81050),
            .I(\pid_side.error_2 ));
    LocalMux I__18704 (
            .O(N__81047),
            .I(\pid_side.error_2 ));
    Odrv4 I__18703 (
            .O(N__81044),
            .I(\pid_side.error_2 ));
    Odrv12 I__18702 (
            .O(N__81041),
            .I(\pid_side.error_2 ));
    LocalMux I__18701 (
            .O(N__81038),
            .I(\pid_side.error_2 ));
    InMux I__18700 (
            .O(N__81025),
            .I(N__81019));
    InMux I__18699 (
            .O(N__81024),
            .I(N__81014));
    InMux I__18698 (
            .O(N__81023),
            .I(N__81014));
    InMux I__18697 (
            .O(N__81022),
            .I(N__81010));
    LocalMux I__18696 (
            .O(N__81019),
            .I(N__81006));
    LocalMux I__18695 (
            .O(N__81014),
            .I(N__81003));
    InMux I__18694 (
            .O(N__81013),
            .I(N__81000));
    LocalMux I__18693 (
            .O(N__81010),
            .I(N__80997));
    InMux I__18692 (
            .O(N__81009),
            .I(N__80994));
    Span4Mux_s1_h I__18691 (
            .O(N__81006),
            .I(N__80991));
    Span4Mux_v I__18690 (
            .O(N__81003),
            .I(N__80986));
    LocalMux I__18689 (
            .O(N__81000),
            .I(N__80986));
    Span4Mux_s1_h I__18688 (
            .O(N__80997),
            .I(N__80983));
    LocalMux I__18687 (
            .O(N__80994),
            .I(N__80980));
    Span4Mux_h I__18686 (
            .O(N__80991),
            .I(N__80972));
    Span4Mux_h I__18685 (
            .O(N__80986),
            .I(N__80972));
    Span4Mux_h I__18684 (
            .O(N__80983),
            .I(N__80967));
    Span4Mux_h I__18683 (
            .O(N__80980),
            .I(N__80967));
    InMux I__18682 (
            .O(N__80979),
            .I(N__80962));
    InMux I__18681 (
            .O(N__80978),
            .I(N__80962));
    InMux I__18680 (
            .O(N__80977),
            .I(N__80959));
    Odrv4 I__18679 (
            .O(N__80972),
            .I(\pid_side.error_1 ));
    Odrv4 I__18678 (
            .O(N__80967),
            .I(\pid_side.error_1 ));
    LocalMux I__18677 (
            .O(N__80962),
            .I(\pid_side.error_1 ));
    LocalMux I__18676 (
            .O(N__80959),
            .I(\pid_side.error_1 ));
    InMux I__18675 (
            .O(N__80950),
            .I(N__80944));
    CascadeMux I__18674 (
            .O(N__80949),
            .I(N__80941));
    InMux I__18673 (
            .O(N__80948),
            .I(N__80937));
    CascadeMux I__18672 (
            .O(N__80947),
            .I(N__80931));
    LocalMux I__18671 (
            .O(N__80944),
            .I(N__80928));
    InMux I__18670 (
            .O(N__80941),
            .I(N__80923));
    InMux I__18669 (
            .O(N__80940),
            .I(N__80923));
    LocalMux I__18668 (
            .O(N__80937),
            .I(N__80920));
    InMux I__18667 (
            .O(N__80936),
            .I(N__80915));
    InMux I__18666 (
            .O(N__80935),
            .I(N__80915));
    InMux I__18665 (
            .O(N__80934),
            .I(N__80912));
    InMux I__18664 (
            .O(N__80931),
            .I(N__80909));
    Span12Mux_v I__18663 (
            .O(N__80928),
            .I(N__80906));
    LocalMux I__18662 (
            .O(N__80923),
            .I(N__80903));
    Span4Mux_v I__18661 (
            .O(N__80920),
            .I(N__80898));
    LocalMux I__18660 (
            .O(N__80915),
            .I(N__80898));
    LocalMux I__18659 (
            .O(N__80912),
            .I(N__80895));
    LocalMux I__18658 (
            .O(N__80909),
            .I(N__80892));
    Span12Mux_h I__18657 (
            .O(N__80906),
            .I(N__80889));
    Span4Mux_h I__18656 (
            .O(N__80903),
            .I(N__80886));
    Span4Mux_h I__18655 (
            .O(N__80898),
            .I(N__80883));
    Span12Mux_s4_h I__18654 (
            .O(N__80895),
            .I(N__80878));
    Span12Mux_v I__18653 (
            .O(N__80892),
            .I(N__80878));
    Odrv12 I__18652 (
            .O(N__80889),
            .I(drone_H_disp_side_0));
    Odrv4 I__18651 (
            .O(N__80886),
            .I(drone_H_disp_side_0));
    Odrv4 I__18650 (
            .O(N__80883),
            .I(drone_H_disp_side_0));
    Odrv12 I__18649 (
            .O(N__80878),
            .I(drone_H_disp_side_0));
    InMux I__18648 (
            .O(N__80869),
            .I(N__80860));
    InMux I__18647 (
            .O(N__80868),
            .I(N__80857));
    InMux I__18646 (
            .O(N__80867),
            .I(N__80854));
    InMux I__18645 (
            .O(N__80866),
            .I(N__80850));
    InMux I__18644 (
            .O(N__80865),
            .I(N__80845));
    InMux I__18643 (
            .O(N__80864),
            .I(N__80845));
    InMux I__18642 (
            .O(N__80863),
            .I(N__80842));
    LocalMux I__18641 (
            .O(N__80860),
            .I(N__80839));
    LocalMux I__18640 (
            .O(N__80857),
            .I(N__80836));
    LocalMux I__18639 (
            .O(N__80854),
            .I(N__80833));
    CascadeMux I__18638 (
            .O(N__80853),
            .I(N__80829));
    LocalMux I__18637 (
            .O(N__80850),
            .I(N__80822));
    LocalMux I__18636 (
            .O(N__80845),
            .I(N__80822));
    LocalMux I__18635 (
            .O(N__80842),
            .I(N__80822));
    Span4Mux_v I__18634 (
            .O(N__80839),
            .I(N__80817));
    Span4Mux_v I__18633 (
            .O(N__80836),
            .I(N__80817));
    Span4Mux_h I__18632 (
            .O(N__80833),
            .I(N__80813));
    InMux I__18631 (
            .O(N__80832),
            .I(N__80810));
    InMux I__18630 (
            .O(N__80829),
            .I(N__80807));
    Span4Mux_v I__18629 (
            .O(N__80822),
            .I(N__80802));
    Span4Mux_h I__18628 (
            .O(N__80817),
            .I(N__80802));
    InMux I__18627 (
            .O(N__80816),
            .I(N__80799));
    Odrv4 I__18626 (
            .O(N__80813),
            .I(\pid_side.error_3 ));
    LocalMux I__18625 (
            .O(N__80810),
            .I(\pid_side.error_3 ));
    LocalMux I__18624 (
            .O(N__80807),
            .I(\pid_side.error_3 ));
    Odrv4 I__18623 (
            .O(N__80802),
            .I(\pid_side.error_3 ));
    LocalMux I__18622 (
            .O(N__80799),
            .I(\pid_side.error_3 ));
    InMux I__18621 (
            .O(N__80788),
            .I(N__80785));
    LocalMux I__18620 (
            .O(N__80785),
            .I(N__80782));
    Span4Mux_v I__18619 (
            .O(N__80782),
            .I(N__80779));
    Odrv4 I__18618 (
            .O(N__80779),
            .I(\pid_side.N_40_0_i_i_o2_1 ));
    CascadeMux I__18617 (
            .O(N__80776),
            .I(\pid_side.N_40_0_i_i_o2_1_cascade_ ));
    InMux I__18616 (
            .O(N__80773),
            .I(N__80770));
    LocalMux I__18615 (
            .O(N__80770),
            .I(N__80766));
    InMux I__18614 (
            .O(N__80769),
            .I(N__80763));
    Span4Mux_v I__18613 (
            .O(N__80766),
            .I(N__80760));
    LocalMux I__18612 (
            .O(N__80763),
            .I(\pid_side.N_40_0_i_i_o2_0 ));
    Odrv4 I__18611 (
            .O(N__80760),
            .I(\pid_side.N_40_0_i_i_o2_0 ));
    InMux I__18610 (
            .O(N__80755),
            .I(N__80752));
    LocalMux I__18609 (
            .O(N__80752),
            .I(N__80749));
    Span4Mux_v I__18608 (
            .O(N__80749),
            .I(N__80746));
    Span4Mux_h I__18607 (
            .O(N__80746),
            .I(N__80743));
    Odrv4 I__18606 (
            .O(N__80743),
            .I(\pid_side.N_27_0_i_i_0 ));
    CascadeMux I__18605 (
            .O(N__80740),
            .I(\pid_side.m7_2_01_ns_1_cascade_ ));
    InMux I__18604 (
            .O(N__80737),
            .I(N__80734));
    LocalMux I__18603 (
            .O(N__80734),
            .I(N__80730));
    InMux I__18602 (
            .O(N__80733),
            .I(N__80727));
    Odrv4 I__18601 (
            .O(N__80730),
            .I(\pid_side.N_162 ));
    LocalMux I__18600 (
            .O(N__80727),
            .I(\pid_side.N_162 ));
    InMux I__18599 (
            .O(N__80722),
            .I(N__80719));
    LocalMux I__18598 (
            .O(N__80719),
            .I(N__80716));
    Sp12to4 I__18597 (
            .O(N__80716),
            .I(N__80713));
    Span12Mux_v I__18596 (
            .O(N__80713),
            .I(N__80710));
    Odrv12 I__18595 (
            .O(N__80710),
            .I(\pid_side.m7_2_01 ));
    CascadeMux I__18594 (
            .O(N__80707),
            .I(\pid_side.m7_2_01_cascade_ ));
    InMux I__18593 (
            .O(N__80704),
            .I(N__80701));
    LocalMux I__18592 (
            .O(N__80701),
            .I(N__80692));
    InMux I__18591 (
            .O(N__80700),
            .I(N__80685));
    InMux I__18590 (
            .O(N__80699),
            .I(N__80685));
    InMux I__18589 (
            .O(N__80698),
            .I(N__80682));
    InMux I__18588 (
            .O(N__80697),
            .I(N__80678));
    InMux I__18587 (
            .O(N__80696),
            .I(N__80674));
    InMux I__18586 (
            .O(N__80695),
            .I(N__80671));
    Span4Mux_v I__18585 (
            .O(N__80692),
            .I(N__80666));
    InMux I__18584 (
            .O(N__80691),
            .I(N__80663));
    InMux I__18583 (
            .O(N__80690),
            .I(N__80660));
    LocalMux I__18582 (
            .O(N__80685),
            .I(N__80656));
    LocalMux I__18581 (
            .O(N__80682),
            .I(N__80653));
    InMux I__18580 (
            .O(N__80681),
            .I(N__80650));
    LocalMux I__18579 (
            .O(N__80678),
            .I(N__80645));
    InMux I__18578 (
            .O(N__80677),
            .I(N__80642));
    LocalMux I__18577 (
            .O(N__80674),
            .I(N__80639));
    LocalMux I__18576 (
            .O(N__80671),
            .I(N__80636));
    InMux I__18575 (
            .O(N__80670),
            .I(N__80631));
    InMux I__18574 (
            .O(N__80669),
            .I(N__80631));
    Span4Mux_h I__18573 (
            .O(N__80666),
            .I(N__80624));
    LocalMux I__18572 (
            .O(N__80663),
            .I(N__80624));
    LocalMux I__18571 (
            .O(N__80660),
            .I(N__80621));
    InMux I__18570 (
            .O(N__80659),
            .I(N__80616));
    Span4Mux_v I__18569 (
            .O(N__80656),
            .I(N__80613));
    Span4Mux_v I__18568 (
            .O(N__80653),
            .I(N__80610));
    LocalMux I__18567 (
            .O(N__80650),
            .I(N__80607));
    InMux I__18566 (
            .O(N__80649),
            .I(N__80602));
    InMux I__18565 (
            .O(N__80648),
            .I(N__80602));
    Span4Mux_v I__18564 (
            .O(N__80645),
            .I(N__80599));
    LocalMux I__18563 (
            .O(N__80642),
            .I(N__80596));
    Span4Mux_h I__18562 (
            .O(N__80639),
            .I(N__80593));
    Span4Mux_v I__18561 (
            .O(N__80636),
            .I(N__80588));
    LocalMux I__18560 (
            .O(N__80631),
            .I(N__80588));
    InMux I__18559 (
            .O(N__80630),
            .I(N__80583));
    InMux I__18558 (
            .O(N__80629),
            .I(N__80583));
    Span4Mux_v I__18557 (
            .O(N__80624),
            .I(N__80578));
    Span4Mux_v I__18556 (
            .O(N__80621),
            .I(N__80578));
    InMux I__18555 (
            .O(N__80620),
            .I(N__80573));
    InMux I__18554 (
            .O(N__80619),
            .I(N__80573));
    LocalMux I__18553 (
            .O(N__80616),
            .I(N__80570));
    Span4Mux_v I__18552 (
            .O(N__80613),
            .I(N__80561));
    Span4Mux_h I__18551 (
            .O(N__80610),
            .I(N__80561));
    Span4Mux_v I__18550 (
            .O(N__80607),
            .I(N__80561));
    LocalMux I__18549 (
            .O(N__80602),
            .I(N__80561));
    Sp12to4 I__18548 (
            .O(N__80599),
            .I(N__80558));
    Span4Mux_h I__18547 (
            .O(N__80596),
            .I(N__80555));
    Span4Mux_v I__18546 (
            .O(N__80593),
            .I(N__80550));
    Span4Mux_h I__18545 (
            .O(N__80588),
            .I(N__80550));
    LocalMux I__18544 (
            .O(N__80583),
            .I(N__80543));
    Sp12to4 I__18543 (
            .O(N__80578),
            .I(N__80543));
    LocalMux I__18542 (
            .O(N__80573),
            .I(N__80543));
    Span4Mux_v I__18541 (
            .O(N__80570),
            .I(N__80538));
    Span4Mux_h I__18540 (
            .O(N__80561),
            .I(N__80538));
    Odrv12 I__18539 (
            .O(N__80558),
            .I(\pid_front.error_15 ));
    Odrv4 I__18538 (
            .O(N__80555),
            .I(\pid_front.error_15 ));
    Odrv4 I__18537 (
            .O(N__80550),
            .I(\pid_front.error_15 ));
    Odrv12 I__18536 (
            .O(N__80543),
            .I(\pid_front.error_15 ));
    Odrv4 I__18535 (
            .O(N__80538),
            .I(\pid_front.error_15 ));
    InMux I__18534 (
            .O(N__80527),
            .I(N__80524));
    LocalMux I__18533 (
            .O(N__80524),
            .I(N__80521));
    Span4Mux_h I__18532 (
            .O(N__80521),
            .I(N__80518));
    Span4Mux_h I__18531 (
            .O(N__80518),
            .I(N__80515));
    Odrv4 I__18530 (
            .O(N__80515),
            .I(\pid_front.error_i_reg_9_N_5L8_0_sx ));
    InMux I__18529 (
            .O(N__80512),
            .I(N__80509));
    LocalMux I__18528 (
            .O(N__80509),
            .I(N__80506));
    Span4Mux_h I__18527 (
            .O(N__80506),
            .I(N__80503));
    Span4Mux_h I__18526 (
            .O(N__80503),
            .I(N__80500));
    Odrv4 I__18525 (
            .O(N__80500),
            .I(\pid_side.N_186_0 ));
    InMux I__18524 (
            .O(N__80497),
            .I(N__80494));
    LocalMux I__18523 (
            .O(N__80494),
            .I(\pid_side.error_i_reg_esr_RNO_5Z0Z_12 ));
    InMux I__18522 (
            .O(N__80491),
            .I(N__80486));
    InMux I__18521 (
            .O(N__80490),
            .I(N__80483));
    InMux I__18520 (
            .O(N__80489),
            .I(N__80480));
    LocalMux I__18519 (
            .O(N__80486),
            .I(N__80476));
    LocalMux I__18518 (
            .O(N__80483),
            .I(N__80473));
    LocalMux I__18517 (
            .O(N__80480),
            .I(N__80469));
    CascadeMux I__18516 (
            .O(N__80479),
            .I(N__80466));
    Span4Mux_s1_h I__18515 (
            .O(N__80476),
            .I(N__80462));
    Span4Mux_s3_h I__18514 (
            .O(N__80473),
            .I(N__80459));
    InMux I__18513 (
            .O(N__80472),
            .I(N__80456));
    Span4Mux_v I__18512 (
            .O(N__80469),
            .I(N__80451));
    InMux I__18511 (
            .O(N__80466),
            .I(N__80446));
    InMux I__18510 (
            .O(N__80465),
            .I(N__80446));
    Span4Mux_h I__18509 (
            .O(N__80462),
            .I(N__80443));
    Span4Mux_v I__18508 (
            .O(N__80459),
            .I(N__80438));
    LocalMux I__18507 (
            .O(N__80456),
            .I(N__80438));
    InMux I__18506 (
            .O(N__80455),
            .I(N__80433));
    InMux I__18505 (
            .O(N__80454),
            .I(N__80433));
    Span4Mux_h I__18504 (
            .O(N__80451),
            .I(N__80428));
    LocalMux I__18503 (
            .O(N__80446),
            .I(N__80428));
    Odrv4 I__18502 (
            .O(N__80443),
            .I(\pid_side.error_9 ));
    Odrv4 I__18501 (
            .O(N__80438),
            .I(\pid_side.error_9 ));
    LocalMux I__18500 (
            .O(N__80433),
            .I(\pid_side.error_9 ));
    Odrv4 I__18499 (
            .O(N__80428),
            .I(\pid_side.error_9 ));
    InMux I__18498 (
            .O(N__80419),
            .I(N__80414));
    InMux I__18497 (
            .O(N__80418),
            .I(N__80411));
    InMux I__18496 (
            .O(N__80417),
            .I(N__80404));
    LocalMux I__18495 (
            .O(N__80414),
            .I(N__80401));
    LocalMux I__18494 (
            .O(N__80411),
            .I(N__80398));
    InMux I__18493 (
            .O(N__80410),
            .I(N__80395));
    InMux I__18492 (
            .O(N__80409),
            .I(N__80388));
    InMux I__18491 (
            .O(N__80408),
            .I(N__80388));
    InMux I__18490 (
            .O(N__80407),
            .I(N__80388));
    LocalMux I__18489 (
            .O(N__80404),
            .I(N__80385));
    Span4Mux_v I__18488 (
            .O(N__80401),
            .I(N__80380));
    Span4Mux_v I__18487 (
            .O(N__80398),
            .I(N__80380));
    LocalMux I__18486 (
            .O(N__80395),
            .I(N__80377));
    LocalMux I__18485 (
            .O(N__80388),
            .I(N__80371));
    Span4Mux_h I__18484 (
            .O(N__80385),
            .I(N__80371));
    Span4Mux_h I__18483 (
            .O(N__80380),
            .I(N__80366));
    Span4Mux_v I__18482 (
            .O(N__80377),
            .I(N__80363));
    InMux I__18481 (
            .O(N__80376),
            .I(N__80360));
    Span4Mux_v I__18480 (
            .O(N__80371),
            .I(N__80357));
    InMux I__18479 (
            .O(N__80370),
            .I(N__80352));
    InMux I__18478 (
            .O(N__80369),
            .I(N__80352));
    Odrv4 I__18477 (
            .O(N__80366),
            .I(\pid_side.error_13 ));
    Odrv4 I__18476 (
            .O(N__80363),
            .I(\pid_side.error_13 ));
    LocalMux I__18475 (
            .O(N__80360),
            .I(\pid_side.error_13 ));
    Odrv4 I__18474 (
            .O(N__80357),
            .I(\pid_side.error_13 ));
    LocalMux I__18473 (
            .O(N__80352),
            .I(\pid_side.error_13 ));
    InMux I__18472 (
            .O(N__80341),
            .I(N__80336));
    InMux I__18471 (
            .O(N__80340),
            .I(N__80333));
    InMux I__18470 (
            .O(N__80339),
            .I(N__80330));
    LocalMux I__18469 (
            .O(N__80336),
            .I(N__80325));
    LocalMux I__18468 (
            .O(N__80333),
            .I(N__80325));
    LocalMux I__18467 (
            .O(N__80330),
            .I(N__80320));
    Span4Mux_h I__18466 (
            .O(N__80325),
            .I(N__80320));
    Odrv4 I__18465 (
            .O(N__80320),
            .I(\pid_side.N_606 ));
    CascadeMux I__18464 (
            .O(N__80317),
            .I(\pid_side.N_606_cascade_ ));
    InMux I__18463 (
            .O(N__80314),
            .I(N__80307));
    InMux I__18462 (
            .O(N__80313),
            .I(N__80304));
    InMux I__18461 (
            .O(N__80312),
            .I(N__80300));
    InMux I__18460 (
            .O(N__80311),
            .I(N__80297));
    InMux I__18459 (
            .O(N__80310),
            .I(N__80294));
    LocalMux I__18458 (
            .O(N__80307),
            .I(N__80291));
    LocalMux I__18457 (
            .O(N__80304),
            .I(N__80288));
    InMux I__18456 (
            .O(N__80303),
            .I(N__80284));
    LocalMux I__18455 (
            .O(N__80300),
            .I(N__80278));
    LocalMux I__18454 (
            .O(N__80297),
            .I(N__80273));
    LocalMux I__18453 (
            .O(N__80294),
            .I(N__80273));
    Span4Mux_v I__18452 (
            .O(N__80291),
            .I(N__80268));
    Span4Mux_v I__18451 (
            .O(N__80288),
            .I(N__80268));
    InMux I__18450 (
            .O(N__80287),
            .I(N__80265));
    LocalMux I__18449 (
            .O(N__80284),
            .I(N__80262));
    InMux I__18448 (
            .O(N__80283),
            .I(N__80257));
    InMux I__18447 (
            .O(N__80282),
            .I(N__80257));
    CascadeMux I__18446 (
            .O(N__80281),
            .I(N__80254));
    Span4Mux_v I__18445 (
            .O(N__80278),
            .I(N__80248));
    Span4Mux_v I__18444 (
            .O(N__80273),
            .I(N__80248));
    Span4Mux_h I__18443 (
            .O(N__80268),
            .I(N__80243));
    LocalMux I__18442 (
            .O(N__80265),
            .I(N__80243));
    Span4Mux_v I__18441 (
            .O(N__80262),
            .I(N__80240));
    LocalMux I__18440 (
            .O(N__80257),
            .I(N__80237));
    InMux I__18439 (
            .O(N__80254),
            .I(N__80232));
    InMux I__18438 (
            .O(N__80253),
            .I(N__80232));
    Span4Mux_h I__18437 (
            .O(N__80248),
            .I(N__80229));
    Odrv4 I__18436 (
            .O(N__80243),
            .I(\pid_side.error_5 ));
    Odrv4 I__18435 (
            .O(N__80240),
            .I(\pid_side.error_5 ));
    Odrv4 I__18434 (
            .O(N__80237),
            .I(\pid_side.error_5 ));
    LocalMux I__18433 (
            .O(N__80232),
            .I(\pid_side.error_5 ));
    Odrv4 I__18432 (
            .O(N__80229),
            .I(\pid_side.error_5 ));
    InMux I__18431 (
            .O(N__80218),
            .I(N__80208));
    InMux I__18430 (
            .O(N__80217),
            .I(N__80208));
    InMux I__18429 (
            .O(N__80216),
            .I(N__80199));
    InMux I__18428 (
            .O(N__80215),
            .I(N__80199));
    CascadeMux I__18427 (
            .O(N__80214),
            .I(N__80195));
    InMux I__18426 (
            .O(N__80213),
            .I(N__80189));
    LocalMux I__18425 (
            .O(N__80208),
            .I(N__80184));
    InMux I__18424 (
            .O(N__80207),
            .I(N__80179));
    InMux I__18423 (
            .O(N__80206),
            .I(N__80179));
    InMux I__18422 (
            .O(N__80205),
            .I(N__80176));
    InMux I__18421 (
            .O(N__80204),
            .I(N__80173));
    LocalMux I__18420 (
            .O(N__80199),
            .I(N__80170));
    InMux I__18419 (
            .O(N__80198),
            .I(N__80167));
    InMux I__18418 (
            .O(N__80195),
            .I(N__80158));
    InMux I__18417 (
            .O(N__80194),
            .I(N__80158));
    InMux I__18416 (
            .O(N__80193),
            .I(N__80158));
    InMux I__18415 (
            .O(N__80192),
            .I(N__80158));
    LocalMux I__18414 (
            .O(N__80189),
            .I(N__80155));
    InMux I__18413 (
            .O(N__80188),
            .I(N__80152));
    InMux I__18412 (
            .O(N__80187),
            .I(N__80149));
    Span4Mux_h I__18411 (
            .O(N__80184),
            .I(N__80142));
    LocalMux I__18410 (
            .O(N__80179),
            .I(N__80142));
    LocalMux I__18409 (
            .O(N__80176),
            .I(N__80142));
    LocalMux I__18408 (
            .O(N__80173),
            .I(N__80139));
    Span4Mux_v I__18407 (
            .O(N__80170),
            .I(N__80136));
    LocalMux I__18406 (
            .O(N__80167),
            .I(N__80130));
    LocalMux I__18405 (
            .O(N__80158),
            .I(N__80130));
    Span4Mux_v I__18404 (
            .O(N__80155),
            .I(N__80121));
    LocalMux I__18403 (
            .O(N__80152),
            .I(N__80121));
    LocalMux I__18402 (
            .O(N__80149),
            .I(N__80121));
    Span4Mux_v I__18401 (
            .O(N__80142),
            .I(N__80121));
    Span4Mux_h I__18400 (
            .O(N__80139),
            .I(N__80114));
    Span4Mux_h I__18399 (
            .O(N__80136),
            .I(N__80114));
    InMux I__18398 (
            .O(N__80135),
            .I(N__80111));
    Span4Mux_h I__18397 (
            .O(N__80130),
            .I(N__80108));
    Span4Mux_h I__18396 (
            .O(N__80121),
            .I(N__80105));
    InMux I__18395 (
            .O(N__80120),
            .I(N__80100));
    InMux I__18394 (
            .O(N__80119),
            .I(N__80100));
    Odrv4 I__18393 (
            .O(N__80114),
            .I(xy_ki_fast_2));
    LocalMux I__18392 (
            .O(N__80111),
            .I(xy_ki_fast_2));
    Odrv4 I__18391 (
            .O(N__80108),
            .I(xy_ki_fast_2));
    Odrv4 I__18390 (
            .O(N__80105),
            .I(xy_ki_fast_2));
    LocalMux I__18389 (
            .O(N__80100),
            .I(xy_ki_fast_2));
    InMux I__18388 (
            .O(N__80089),
            .I(N__80086));
    LocalMux I__18387 (
            .O(N__80086),
            .I(N__80083));
    Odrv12 I__18386 (
            .O(N__80083),
            .I(\pid_side.N_188 ));
    InMux I__18385 (
            .O(N__80080),
            .I(N__80074));
    InMux I__18384 (
            .O(N__80079),
            .I(N__80074));
    LocalMux I__18383 (
            .O(N__80074),
            .I(N__80070));
    InMux I__18382 (
            .O(N__80073),
            .I(N__80067));
    Span4Mux_h I__18381 (
            .O(N__80070),
            .I(N__80064));
    LocalMux I__18380 (
            .O(N__80067),
            .I(\pid_side.N_231 ));
    Odrv4 I__18379 (
            .O(N__80064),
            .I(\pid_side.N_231 ));
    CascadeMux I__18378 (
            .O(N__80059),
            .I(\pid_side.N_231_cascade_ ));
    InMux I__18377 (
            .O(N__80056),
            .I(N__80053));
    LocalMux I__18376 (
            .O(N__80053),
            .I(N__80048));
    InMux I__18375 (
            .O(N__80052),
            .I(N__80045));
    InMux I__18374 (
            .O(N__80051),
            .I(N__80042));
    Span4Mux_h I__18373 (
            .O(N__80048),
            .I(N__80039));
    LocalMux I__18372 (
            .O(N__80045),
            .I(\pid_side.N_184 ));
    LocalMux I__18371 (
            .O(N__80042),
            .I(\pid_side.N_184 ));
    Odrv4 I__18370 (
            .O(N__80039),
            .I(\pid_side.N_184 ));
    InMux I__18369 (
            .O(N__80032),
            .I(N__80029));
    LocalMux I__18368 (
            .O(N__80029),
            .I(N__80026));
    Span4Mux_h I__18367 (
            .O(N__80026),
            .I(N__80023));
    Span4Mux_h I__18366 (
            .O(N__80023),
            .I(N__80020));
    Odrv4 I__18365 (
            .O(N__80020),
            .I(\pid_side.N_339 ));
    InMux I__18364 (
            .O(N__80017),
            .I(N__80014));
    LocalMux I__18363 (
            .O(N__80014),
            .I(N__80008));
    InMux I__18362 (
            .O(N__80013),
            .I(N__80005));
    InMux I__18361 (
            .O(N__80012),
            .I(N__79999));
    InMux I__18360 (
            .O(N__80011),
            .I(N__79995));
    Span4Mux_v I__18359 (
            .O(N__80008),
            .I(N__79992));
    LocalMux I__18358 (
            .O(N__80005),
            .I(N__79989));
    InMux I__18357 (
            .O(N__80004),
            .I(N__79986));
    InMux I__18356 (
            .O(N__80003),
            .I(N__79983));
    InMux I__18355 (
            .O(N__80002),
            .I(N__79980));
    LocalMux I__18354 (
            .O(N__79999),
            .I(N__79977));
    InMux I__18353 (
            .O(N__79998),
            .I(N__79974));
    LocalMux I__18352 (
            .O(N__79995),
            .I(N__79968));
    Sp12to4 I__18351 (
            .O(N__79992),
            .I(N__79965));
    Span12Mux_v I__18350 (
            .O(N__79989),
            .I(N__79962));
    LocalMux I__18349 (
            .O(N__79986),
            .I(N__79957));
    LocalMux I__18348 (
            .O(N__79983),
            .I(N__79957));
    LocalMux I__18347 (
            .O(N__79980),
            .I(N__79954));
    Span4Mux_h I__18346 (
            .O(N__79977),
            .I(N__79949));
    LocalMux I__18345 (
            .O(N__79974),
            .I(N__79949));
    InMux I__18344 (
            .O(N__79973),
            .I(N__79942));
    InMux I__18343 (
            .O(N__79972),
            .I(N__79942));
    InMux I__18342 (
            .O(N__79971),
            .I(N__79942));
    Span4Mux_h I__18341 (
            .O(N__79968),
            .I(N__79939));
    Span12Mux_h I__18340 (
            .O(N__79965),
            .I(N__79932));
    Span12Mux_h I__18339 (
            .O(N__79962),
            .I(N__79932));
    Span12Mux_h I__18338 (
            .O(N__79957),
            .I(N__79932));
    Span4Mux_v I__18337 (
            .O(N__79954),
            .I(N__79927));
    Span4Mux_h I__18336 (
            .O(N__79949),
            .I(N__79927));
    LocalMux I__18335 (
            .O(N__79942),
            .I(N__79922));
    Span4Mux_h I__18334 (
            .O(N__79939),
            .I(N__79922));
    Odrv12 I__18333 (
            .O(N__79932),
            .I(\pid_front.error_2 ));
    Odrv4 I__18332 (
            .O(N__79927),
            .I(\pid_front.error_2 ));
    Odrv4 I__18331 (
            .O(N__79922),
            .I(\pid_front.error_2 ));
    InMux I__18330 (
            .O(N__79915),
            .I(N__79909));
    InMux I__18329 (
            .O(N__79914),
            .I(N__79906));
    InMux I__18328 (
            .O(N__79913),
            .I(N__79900));
    InMux I__18327 (
            .O(N__79912),
            .I(N__79897));
    LocalMux I__18326 (
            .O(N__79909),
            .I(N__79894));
    LocalMux I__18325 (
            .O(N__79906),
            .I(N__79891));
    InMux I__18324 (
            .O(N__79905),
            .I(N__79885));
    InMux I__18323 (
            .O(N__79904),
            .I(N__79885));
    InMux I__18322 (
            .O(N__79903),
            .I(N__79880));
    LocalMux I__18321 (
            .O(N__79900),
            .I(N__79877));
    LocalMux I__18320 (
            .O(N__79897),
            .I(N__79874));
    Span4Mux_v I__18319 (
            .O(N__79894),
            .I(N__79871));
    Span4Mux_s1_h I__18318 (
            .O(N__79891),
            .I(N__79868));
    CascadeMux I__18317 (
            .O(N__79890),
            .I(N__79865));
    LocalMux I__18316 (
            .O(N__79885),
            .I(N__79862));
    InMux I__18315 (
            .O(N__79884),
            .I(N__79857));
    InMux I__18314 (
            .O(N__79883),
            .I(N__79857));
    LocalMux I__18313 (
            .O(N__79880),
            .I(N__79852));
    Span4Mux_v I__18312 (
            .O(N__79877),
            .I(N__79847));
    Span4Mux_v I__18311 (
            .O(N__79874),
            .I(N__79847));
    Span4Mux_h I__18310 (
            .O(N__79871),
            .I(N__79844));
    Span4Mux_h I__18309 (
            .O(N__79868),
            .I(N__79841));
    InMux I__18308 (
            .O(N__79865),
            .I(N__79838));
    Span4Mux_h I__18307 (
            .O(N__79862),
            .I(N__79835));
    LocalMux I__18306 (
            .O(N__79857),
            .I(N__79832));
    InMux I__18305 (
            .O(N__79856),
            .I(N__79829));
    InMux I__18304 (
            .O(N__79855),
            .I(N__79826));
    Span4Mux_v I__18303 (
            .O(N__79852),
            .I(N__79821));
    Span4Mux_h I__18302 (
            .O(N__79847),
            .I(N__79821));
    Span4Mux_h I__18301 (
            .O(N__79844),
            .I(N__79818));
    Span4Mux_h I__18300 (
            .O(N__79841),
            .I(N__79815));
    LocalMux I__18299 (
            .O(N__79838),
            .I(N__79812));
    Span4Mux_h I__18298 (
            .O(N__79835),
            .I(N__79809));
    Span4Mux_v I__18297 (
            .O(N__79832),
            .I(N__79806));
    LocalMux I__18296 (
            .O(N__79829),
            .I(N__79803));
    LocalMux I__18295 (
            .O(N__79826),
            .I(N__79794));
    Span4Mux_h I__18294 (
            .O(N__79821),
            .I(N__79794));
    Span4Mux_h I__18293 (
            .O(N__79818),
            .I(N__79794));
    Span4Mux_h I__18292 (
            .O(N__79815),
            .I(N__79794));
    Odrv4 I__18291 (
            .O(N__79812),
            .I(\pid_front.error_4 ));
    Odrv4 I__18290 (
            .O(N__79809),
            .I(\pid_front.error_4 ));
    Odrv4 I__18289 (
            .O(N__79806),
            .I(\pid_front.error_4 ));
    Odrv12 I__18288 (
            .O(N__79803),
            .I(\pid_front.error_4 ));
    Odrv4 I__18287 (
            .O(N__79794),
            .I(\pid_front.error_4 ));
    InMux I__18286 (
            .O(N__79783),
            .I(N__79779));
    InMux I__18285 (
            .O(N__79782),
            .I(N__79776));
    LocalMux I__18284 (
            .O(N__79779),
            .I(N__79773));
    LocalMux I__18283 (
            .O(N__79776),
            .I(N__79770));
    Span4Mux_h I__18282 (
            .O(N__79773),
            .I(N__79767));
    Span4Mux_h I__18281 (
            .O(N__79770),
            .I(N__79764));
    Odrv4 I__18280 (
            .O(N__79767),
            .I(\pid_front.N_525 ));
    Odrv4 I__18279 (
            .O(N__79764),
            .I(\pid_front.N_525 ));
    CascadeMux I__18278 (
            .O(N__79759),
            .I(\pid_side.m24_2_03_0_0_cascade_ ));
    CascadeMux I__18277 (
            .O(N__79756),
            .I(\pid_side.error_i_reg_esr_RNO_6Z0Z_20_cascade_ ));
    InMux I__18276 (
            .O(N__79753),
            .I(N__79750));
    LocalMux I__18275 (
            .O(N__79750),
            .I(\pid_side.error_i_reg_esr_RNO_5Z0Z_20 ));
    InMux I__18274 (
            .O(N__79747),
            .I(N__79744));
    LocalMux I__18273 (
            .O(N__79744),
            .I(\pid_side.m24_2_03_0_1 ));
    CascadeMux I__18272 (
            .O(N__79741),
            .I(\pid_side.N_162_cascade_ ));
    InMux I__18271 (
            .O(N__79738),
            .I(N__79734));
    InMux I__18270 (
            .O(N__79737),
            .I(N__79731));
    LocalMux I__18269 (
            .O(N__79734),
            .I(N__79728));
    LocalMux I__18268 (
            .O(N__79731),
            .I(N__79725));
    Span4Mux_v I__18267 (
            .O(N__79728),
            .I(N__79722));
    Span4Mux_v I__18266 (
            .O(N__79725),
            .I(N__79717));
    Span4Mux_h I__18265 (
            .O(N__79722),
            .I(N__79717));
    Odrv4 I__18264 (
            .O(N__79717),
            .I(\pid_side.N_206 ));
    CascadeMux I__18263 (
            .O(N__79714),
            .I(\pid_side.N_206_cascade_ ));
    InMux I__18262 (
            .O(N__79711),
            .I(N__79707));
    InMux I__18261 (
            .O(N__79710),
            .I(N__79704));
    LocalMux I__18260 (
            .O(N__79707),
            .I(N__79701));
    LocalMux I__18259 (
            .O(N__79704),
            .I(\pid_side.N_629 ));
    Odrv12 I__18258 (
            .O(N__79701),
            .I(\pid_side.N_629 ));
    InMux I__18257 (
            .O(N__79696),
            .I(N__79693));
    LocalMux I__18256 (
            .O(N__79693),
            .I(N__79690));
    Span4Mux_h I__18255 (
            .O(N__79690),
            .I(N__79687));
    Odrv4 I__18254 (
            .O(N__79687),
            .I(\pid_side.m9_2_03_3_i_0_o2_0 ));
    CascadeMux I__18253 (
            .O(N__79684),
            .I(\pid_side.m9_2_03_3_i_0_o2_2_cascade_ ));
    CascadeMux I__18252 (
            .O(N__79681),
            .I(N__79678));
    InMux I__18251 (
            .O(N__79678),
            .I(N__79675));
    LocalMux I__18250 (
            .O(N__79675),
            .I(N__79672));
    Span4Mux_h I__18249 (
            .O(N__79672),
            .I(N__79669));
    Span4Mux_v I__18248 (
            .O(N__79669),
            .I(N__79666));
    Span4Mux_h I__18247 (
            .O(N__79666),
            .I(N__79663));
    Odrv4 I__18246 (
            .O(N__79663),
            .I(\pid_side.error_i_regZ0Z_5 ));
    CascadeMux I__18245 (
            .O(N__79660),
            .I(N__79656));
    CascadeMux I__18244 (
            .O(N__79659),
            .I(N__79651));
    InMux I__18243 (
            .O(N__79656),
            .I(N__79647));
    InMux I__18242 (
            .O(N__79655),
            .I(N__79644));
    CascadeMux I__18241 (
            .O(N__79654),
            .I(N__79641));
    InMux I__18240 (
            .O(N__79651),
            .I(N__79638));
    CascadeMux I__18239 (
            .O(N__79650),
            .I(N__79635));
    LocalMux I__18238 (
            .O(N__79647),
            .I(N__79630));
    LocalMux I__18237 (
            .O(N__79644),
            .I(N__79630));
    InMux I__18236 (
            .O(N__79641),
            .I(N__79627));
    LocalMux I__18235 (
            .O(N__79638),
            .I(N__79622));
    InMux I__18234 (
            .O(N__79635),
            .I(N__79619));
    Span4Mux_h I__18233 (
            .O(N__79630),
            .I(N__79616));
    LocalMux I__18232 (
            .O(N__79627),
            .I(N__79613));
    CascadeMux I__18231 (
            .O(N__79626),
            .I(N__79609));
    InMux I__18230 (
            .O(N__79625),
            .I(N__79606));
    Span4Mux_v I__18229 (
            .O(N__79622),
            .I(N__79603));
    LocalMux I__18228 (
            .O(N__79619),
            .I(N__79596));
    Span4Mux_v I__18227 (
            .O(N__79616),
            .I(N__79596));
    Span4Mux_h I__18226 (
            .O(N__79613),
            .I(N__79596));
    InMux I__18225 (
            .O(N__79612),
            .I(N__79591));
    InMux I__18224 (
            .O(N__79609),
            .I(N__79591));
    LocalMux I__18223 (
            .O(N__79606),
            .I(N__79588));
    Odrv4 I__18222 (
            .O(N__79603),
            .I(xy_ki_fast_3_rep1));
    Odrv4 I__18221 (
            .O(N__79596),
            .I(xy_ki_fast_3_rep1));
    LocalMux I__18220 (
            .O(N__79591),
            .I(xy_ki_fast_3_rep1));
    Odrv12 I__18219 (
            .O(N__79588),
            .I(xy_ki_fast_3_rep1));
    CascadeMux I__18218 (
            .O(N__79579),
            .I(pid_side_N_496_cascade_));
    InMux I__18217 (
            .O(N__79576),
            .I(N__79572));
    InMux I__18216 (
            .O(N__79575),
            .I(N__79569));
    LocalMux I__18215 (
            .O(N__79572),
            .I(N__79566));
    LocalMux I__18214 (
            .O(N__79569),
            .I(N__79561));
    Span4Mux_v I__18213 (
            .O(N__79566),
            .I(N__79561));
    Odrv4 I__18212 (
            .O(N__79561),
            .I(\pid_side.N_536 ));
    CascadeMux I__18211 (
            .O(N__79558),
            .I(\pid_side.N_8_cascade_ ));
    CascadeMux I__18210 (
            .O(N__79555),
            .I(\pid_side.error_i_reg_esr_RNO_0Z0Z_18_cascade_ ));
    CascadeMux I__18209 (
            .O(N__79552),
            .I(N__79549));
    InMux I__18208 (
            .O(N__79549),
            .I(N__79546));
    LocalMux I__18207 (
            .O(N__79546),
            .I(N__79543));
    Span4Mux_v I__18206 (
            .O(N__79543),
            .I(N__79540));
    Span4Mux_h I__18205 (
            .O(N__79540),
            .I(N__79537));
    Odrv4 I__18204 (
            .O(N__79537),
            .I(\pid_side.error_i_regZ0Z_18 ));
    InMux I__18203 (
            .O(N__79534),
            .I(N__79531));
    LocalMux I__18202 (
            .O(N__79531),
            .I(\pid_side.m22_2_03_0_2 ));
    InMux I__18201 (
            .O(N__79528),
            .I(N__79522));
    InMux I__18200 (
            .O(N__79527),
            .I(N__79522));
    LocalMux I__18199 (
            .O(N__79522),
            .I(N__79519));
    Span4Mux_v I__18198 (
            .O(N__79519),
            .I(N__79516));
    Span4Mux_h I__18197 (
            .O(N__79516),
            .I(N__79513));
    Odrv4 I__18196 (
            .O(N__79513),
            .I(\pid_side.error_cry_1_c_RNI6K4BZ0Z1 ));
    InMux I__18195 (
            .O(N__79510),
            .I(N__79507));
    LocalMux I__18194 (
            .O(N__79507),
            .I(\pid_side.N_8 ));
    CascadeMux I__18193 (
            .O(N__79504),
            .I(N__79501));
    InMux I__18192 (
            .O(N__79501),
            .I(N__79498));
    LocalMux I__18191 (
            .O(N__79498),
            .I(N__79495));
    Span4Mux_h I__18190 (
            .O(N__79495),
            .I(N__79492));
    Span4Mux_h I__18189 (
            .O(N__79492),
            .I(N__79489));
    Odrv4 I__18188 (
            .O(N__79489),
            .I(\pid_side.error_i_regZ0Z_2 ));
    InMux I__18187 (
            .O(N__79486),
            .I(N__79483));
    LocalMux I__18186 (
            .O(N__79483),
            .I(N__79480));
    Span4Mux_v I__18185 (
            .O(N__79480),
            .I(N__79477));
    Span4Mux_v I__18184 (
            .O(N__79477),
            .I(N__79474));
    Odrv4 I__18183 (
            .O(N__79474),
            .I(\pid_front.error_i_reg_9_sn_sn_15 ));
    CascadeMux I__18182 (
            .O(N__79471),
            .I(\pid_side.N_314_cascade_ ));
    InMux I__18181 (
            .O(N__79468),
            .I(N__79463));
    InMux I__18180 (
            .O(N__79467),
            .I(N__79460));
    InMux I__18179 (
            .O(N__79466),
            .I(N__79457));
    LocalMux I__18178 (
            .O(N__79463),
            .I(N__79454));
    LocalMux I__18177 (
            .O(N__79460),
            .I(N__79447));
    LocalMux I__18176 (
            .O(N__79457),
            .I(N__79447));
    Span4Mux_v I__18175 (
            .O(N__79454),
            .I(N__79442));
    InMux I__18174 (
            .O(N__79453),
            .I(N__79437));
    InMux I__18173 (
            .O(N__79452),
            .I(N__79437));
    Span4Mux_h I__18172 (
            .O(N__79447),
            .I(N__79434));
    InMux I__18171 (
            .O(N__79446),
            .I(N__79429));
    InMux I__18170 (
            .O(N__79445),
            .I(N__79429));
    Odrv4 I__18169 (
            .O(N__79442),
            .I(\pid_side.error_d_reg_prevZ0Z_12 ));
    LocalMux I__18168 (
            .O(N__79437),
            .I(\pid_side.error_d_reg_prevZ0Z_12 ));
    Odrv4 I__18167 (
            .O(N__79434),
            .I(\pid_side.error_d_reg_prevZ0Z_12 ));
    LocalMux I__18166 (
            .O(N__79429),
            .I(\pid_side.error_d_reg_prevZ0Z_12 ));
    CascadeMux I__18165 (
            .O(N__79420),
            .I(\pid_side.g0_1_0_1_cascade_ ));
    InMux I__18164 (
            .O(N__79417),
            .I(N__79414));
    LocalMux I__18163 (
            .O(N__79414),
            .I(\pid_side.g0_1 ));
    InMux I__18162 (
            .O(N__79411),
            .I(N__79408));
    LocalMux I__18161 (
            .O(N__79408),
            .I(N__79405));
    Span4Mux_h I__18160 (
            .O(N__79405),
            .I(N__79402));
    Odrv4 I__18159 (
            .O(N__79402),
            .I(\pid_side.O_0_3 ));
    InMux I__18158 (
            .O(N__79399),
            .I(N__79395));
    InMux I__18157 (
            .O(N__79398),
            .I(N__79392));
    LocalMux I__18156 (
            .O(N__79395),
            .I(N__79387));
    LocalMux I__18155 (
            .O(N__79392),
            .I(N__79387));
    Span4Mux_h I__18154 (
            .O(N__79387),
            .I(N__79381));
    InMux I__18153 (
            .O(N__79386),
            .I(N__79374));
    InMux I__18152 (
            .O(N__79385),
            .I(N__79374));
    InMux I__18151 (
            .O(N__79384),
            .I(N__79374));
    Odrv4 I__18150 (
            .O(N__79381),
            .I(\pid_side.error_d_regZ0Z_0 ));
    LocalMux I__18149 (
            .O(N__79374),
            .I(\pid_side.error_d_regZ0Z_0 ));
    InMux I__18148 (
            .O(N__79369),
            .I(N__79366));
    LocalMux I__18147 (
            .O(N__79366),
            .I(N__79363));
    Span4Mux_h I__18146 (
            .O(N__79363),
            .I(N__79360));
    Odrv4 I__18145 (
            .O(N__79360),
            .I(\pid_side.O_1_4 ));
    InMux I__18144 (
            .O(N__79357),
            .I(N__79354));
    LocalMux I__18143 (
            .O(N__79354),
            .I(N__79351));
    Span4Mux_v I__18142 (
            .O(N__79351),
            .I(N__79348));
    Odrv4 I__18141 (
            .O(N__79348),
            .I(\pid_side.O_2_6 ));
    InMux I__18140 (
            .O(N__79345),
            .I(N__79341));
    InMux I__18139 (
            .O(N__79344),
            .I(N__79338));
    LocalMux I__18138 (
            .O(N__79341),
            .I(N__79335));
    LocalMux I__18137 (
            .O(N__79338),
            .I(N__79332));
    Odrv4 I__18136 (
            .O(N__79335),
            .I(\pid_side.error_p_regZ0Z_2 ));
    Odrv4 I__18135 (
            .O(N__79332),
            .I(\pid_side.error_p_regZ0Z_2 ));
    InMux I__18134 (
            .O(N__79327),
            .I(N__79322));
    InMux I__18133 (
            .O(N__79326),
            .I(N__79317));
    InMux I__18132 (
            .O(N__79325),
            .I(N__79317));
    LocalMux I__18131 (
            .O(N__79322),
            .I(N__79313));
    LocalMux I__18130 (
            .O(N__79317),
            .I(N__79310));
    InMux I__18129 (
            .O(N__79316),
            .I(N__79307));
    Span4Mux_v I__18128 (
            .O(N__79313),
            .I(N__79302));
    Span4Mux_v I__18127 (
            .O(N__79310),
            .I(N__79302));
    LocalMux I__18126 (
            .O(N__79307),
            .I(\pid_side.error_d_reg_fastZ0Z_12 ));
    Odrv4 I__18125 (
            .O(N__79302),
            .I(\pid_side.error_d_reg_fastZ0Z_12 ));
    InMux I__18124 (
            .O(N__79297),
            .I(N__79294));
    LocalMux I__18123 (
            .O(N__79294),
            .I(N__79291));
    Span4Mux_h I__18122 (
            .O(N__79291),
            .I(N__79288));
    Odrv4 I__18121 (
            .O(N__79288),
            .I(\pid_side.O_1_5 ));
    InMux I__18120 (
            .O(N__79285),
            .I(N__79279));
    InMux I__18119 (
            .O(N__79284),
            .I(N__79279));
    LocalMux I__18118 (
            .O(N__79279),
            .I(N__79276));
    Span4Mux_h I__18117 (
            .O(N__79276),
            .I(N__79272));
    InMux I__18116 (
            .O(N__79275),
            .I(N__79269));
    Odrv4 I__18115 (
            .O(N__79272),
            .I(\pid_side.error_d_regZ0Z_2 ));
    LocalMux I__18114 (
            .O(N__79269),
            .I(\pid_side.error_d_regZ0Z_2 ));
    InMux I__18113 (
            .O(N__79264),
            .I(N__79261));
    LocalMux I__18112 (
            .O(N__79261),
            .I(N__79258));
    Span4Mux_h I__18111 (
            .O(N__79258),
            .I(N__79255));
    Odrv4 I__18110 (
            .O(N__79255),
            .I(\pid_side.N_232 ));
    CascadeMux I__18109 (
            .O(N__79252),
            .I(\pid_side.N_45_i_i_0_cascade_ ));
    InMux I__18108 (
            .O(N__79249),
            .I(N__79243));
    InMux I__18107 (
            .O(N__79248),
            .I(N__79243));
    LocalMux I__18106 (
            .O(N__79243),
            .I(\pid_side.error_p_reg_esr_RNIFEEQZ0Z_3 ));
    InMux I__18105 (
            .O(N__79240),
            .I(N__79237));
    LocalMux I__18104 (
            .O(N__79237),
            .I(N__79234));
    Span4Mux_v I__18103 (
            .O(N__79234),
            .I(N__79231));
    Span4Mux_h I__18102 (
            .O(N__79231),
            .I(N__79228));
    Odrv4 I__18101 (
            .O(N__79228),
            .I(\pid_side.O_1_12 ));
    InMux I__18100 (
            .O(N__79225),
            .I(N__79214));
    InMux I__18099 (
            .O(N__79224),
            .I(N__79214));
    InMux I__18098 (
            .O(N__79223),
            .I(N__79214));
    InMux I__18097 (
            .O(N__79222),
            .I(N__79209));
    InMux I__18096 (
            .O(N__79221),
            .I(N__79209));
    LocalMux I__18095 (
            .O(N__79214),
            .I(N__79206));
    LocalMux I__18094 (
            .O(N__79209),
            .I(N__79203));
    Odrv4 I__18093 (
            .O(N__79206),
            .I(\pid_side.error_d_regZ0Z_9 ));
    Odrv12 I__18092 (
            .O(N__79203),
            .I(\pid_side.error_d_regZ0Z_9 ));
    InMux I__18091 (
            .O(N__79198),
            .I(N__79195));
    LocalMux I__18090 (
            .O(N__79195),
            .I(N__79192));
    Span12Mux_h I__18089 (
            .O(N__79192),
            .I(N__79189));
    Odrv12 I__18088 (
            .O(N__79189),
            .I(\pid_side.O_1_6 ));
    InMux I__18087 (
            .O(N__79186),
            .I(N__79177));
    InMux I__18086 (
            .O(N__79185),
            .I(N__79177));
    InMux I__18085 (
            .O(N__79184),
            .I(N__79177));
    LocalMux I__18084 (
            .O(N__79177),
            .I(\pid_side.error_d_regZ0Z_3 ));
    InMux I__18083 (
            .O(N__79174),
            .I(N__79170));
    InMux I__18082 (
            .O(N__79173),
            .I(N__79165));
    LocalMux I__18081 (
            .O(N__79170),
            .I(N__79162));
    InMux I__18080 (
            .O(N__79169),
            .I(N__79157));
    InMux I__18079 (
            .O(N__79168),
            .I(N__79157));
    LocalMux I__18078 (
            .O(N__79165),
            .I(N__79154));
    Span4Mux_h I__18077 (
            .O(N__79162),
            .I(N__79149));
    LocalMux I__18076 (
            .O(N__79157),
            .I(N__79149));
    Span4Mux_h I__18075 (
            .O(N__79154),
            .I(N__79144));
    Span4Mux_h I__18074 (
            .O(N__79149),
            .I(N__79144));
    Odrv4 I__18073 (
            .O(N__79144),
            .I(\pid_side.error_d_reg_prevZ0Z_14 ));
    CascadeMux I__18072 (
            .O(N__79141),
            .I(\pid_side.N_2608_0_0_0_cascade_ ));
    InMux I__18071 (
            .O(N__79138),
            .I(N__79135));
    LocalMux I__18070 (
            .O(N__79135),
            .I(\pid_side.N_5_1 ));
    CascadeMux I__18069 (
            .O(N__79132),
            .I(\pid_side.g0_2_0_cascade_ ));
    InMux I__18068 (
            .O(N__79129),
            .I(N__79126));
    LocalMux I__18067 (
            .O(N__79126),
            .I(\pid_side.error_d_reg_prev_esr_RNI7PM14Z0Z_12 ));
    InMux I__18066 (
            .O(N__79123),
            .I(N__79113));
    InMux I__18065 (
            .O(N__79122),
            .I(N__79113));
    InMux I__18064 (
            .O(N__79121),
            .I(N__79110));
    CascadeMux I__18063 (
            .O(N__79120),
            .I(N__79107));
    InMux I__18062 (
            .O(N__79119),
            .I(N__79100));
    InMux I__18061 (
            .O(N__79118),
            .I(N__79100));
    LocalMux I__18060 (
            .O(N__79113),
            .I(N__79095));
    LocalMux I__18059 (
            .O(N__79110),
            .I(N__79095));
    InMux I__18058 (
            .O(N__79107),
            .I(N__79088));
    InMux I__18057 (
            .O(N__79106),
            .I(N__79088));
    InMux I__18056 (
            .O(N__79105),
            .I(N__79088));
    LocalMux I__18055 (
            .O(N__79100),
            .I(\pid_side.error_d_reg_prevZ0Z_13 ));
    Odrv12 I__18054 (
            .O(N__79095),
            .I(\pid_side.error_d_reg_prevZ0Z_13 ));
    LocalMux I__18053 (
            .O(N__79088),
            .I(\pid_side.error_d_reg_prevZ0Z_13 ));
    InMux I__18052 (
            .O(N__79081),
            .I(N__79078));
    LocalMux I__18051 (
            .O(N__79078),
            .I(N__79075));
    Odrv4 I__18050 (
            .O(N__79075),
            .I(\pid_side.N_4_1_0_1 ));
    InMux I__18049 (
            .O(N__79072),
            .I(N__79069));
    LocalMux I__18048 (
            .O(N__79069),
            .I(N__79066));
    Span4Mux_h I__18047 (
            .O(N__79066),
            .I(N__79063));
    Span4Mux_v I__18046 (
            .O(N__79063),
            .I(N__79060));
    Span4Mux_v I__18045 (
            .O(N__79060),
            .I(N__79057));
    Odrv4 I__18044 (
            .O(N__79057),
            .I(\pid_side.O_1_10 ));
    InMux I__18043 (
            .O(N__79054),
            .I(N__79048));
    InMux I__18042 (
            .O(N__79053),
            .I(N__79048));
    LocalMux I__18041 (
            .O(N__79048),
            .I(N__79043));
    InMux I__18040 (
            .O(N__79047),
            .I(N__79038));
    InMux I__18039 (
            .O(N__79046),
            .I(N__79038));
    Span4Mux_v I__18038 (
            .O(N__79043),
            .I(N__79033));
    LocalMux I__18037 (
            .O(N__79038),
            .I(N__79033));
    Span4Mux_v I__18036 (
            .O(N__79033),
            .I(N__79030));
    Odrv4 I__18035 (
            .O(N__79030),
            .I(\pid_side.error_d_regZ0Z_7 ));
    InMux I__18034 (
            .O(N__79027),
            .I(N__79024));
    LocalMux I__18033 (
            .O(N__79024),
            .I(N__79021));
    Span4Mux_h I__18032 (
            .O(N__79021),
            .I(N__79018));
    Odrv4 I__18031 (
            .O(N__79018),
            .I(\pid_side.O_2_7 ));
    InMux I__18030 (
            .O(N__79015),
            .I(N__79011));
    CascadeMux I__18029 (
            .O(N__79014),
            .I(N__79008));
    LocalMux I__18028 (
            .O(N__79011),
            .I(N__79005));
    InMux I__18027 (
            .O(N__79008),
            .I(N__79002));
    Span4Mux_h I__18026 (
            .O(N__79005),
            .I(N__78999));
    LocalMux I__18025 (
            .O(N__79002),
            .I(N__78996));
    Span4Mux_v I__18024 (
            .O(N__78999),
            .I(N__78993));
    Odrv4 I__18023 (
            .O(N__78996),
            .I(\pid_side.error_d_reg_prev_esr_RNI9BFR3Z0Z_1 ));
    Odrv4 I__18022 (
            .O(N__78993),
            .I(\pid_side.error_d_reg_prev_esr_RNI9BFR3Z0Z_1 ));
    CascadeMux I__18021 (
            .O(N__78988),
            .I(N__78985));
    InMux I__18020 (
            .O(N__78985),
            .I(N__78982));
    LocalMux I__18019 (
            .O(N__78982),
            .I(N__78979));
    Span4Mux_h I__18018 (
            .O(N__78979),
            .I(N__78976));
    Span4Mux_h I__18017 (
            .O(N__78976),
            .I(N__78973));
    Odrv4 I__18016 (
            .O(N__78973),
            .I(\pid_side.error_p_reg_esr_RNIU3T36Z0Z_2 ));
    InMux I__18015 (
            .O(N__78970),
            .I(N__78967));
    LocalMux I__18014 (
            .O(N__78967),
            .I(\pid_side.error_p_reg_esr_RNICBEQZ0Z_2 ));
    CascadeMux I__18013 (
            .O(N__78964),
            .I(\pid_side.error_p_reg_esr_RNICBEQZ0Z_2_cascade_ ));
    InMux I__18012 (
            .O(N__78961),
            .I(N__78954));
    InMux I__18011 (
            .O(N__78960),
            .I(N__78954));
    InMux I__18010 (
            .O(N__78959),
            .I(N__78951));
    LocalMux I__18009 (
            .O(N__78954),
            .I(N__78948));
    LocalMux I__18008 (
            .O(N__78951),
            .I(N__78945));
    Span12Mux_s5_h I__18007 (
            .O(N__78948),
            .I(N__78942));
    Odrv4 I__18006 (
            .O(N__78945),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_2_c_RNIQUGJ ));
    Odrv12 I__18005 (
            .O(N__78942),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_2_c_RNIQUGJ ));
    CascadeMux I__18004 (
            .O(N__78937),
            .I(N__78934));
    InMux I__18003 (
            .O(N__78934),
            .I(N__78931));
    LocalMux I__18002 (
            .O(N__78931),
            .I(N__78928));
    Span4Mux_h I__18001 (
            .O(N__78928),
            .I(N__78924));
    InMux I__18000 (
            .O(N__78927),
            .I(N__78921));
    Span4Mux_h I__17999 (
            .O(N__78924),
            .I(N__78918));
    LocalMux I__17998 (
            .O(N__78921),
            .I(\pid_side.error_p_reg_esr_RNILOD82Z0Z_2 ));
    Odrv4 I__17997 (
            .O(N__78918),
            .I(\pid_side.error_p_reg_esr_RNILOD82Z0Z_2 ));
    InMux I__17996 (
            .O(N__78913),
            .I(N__78907));
    InMux I__17995 (
            .O(N__78912),
            .I(N__78907));
    LocalMux I__17994 (
            .O(N__78907),
            .I(\pid_side.error_p_reg_esr_RNIFEEQ_0Z0Z_3 ));
    InMux I__17993 (
            .O(N__78904),
            .I(N__78900));
    InMux I__17992 (
            .O(N__78903),
            .I(N__78897));
    LocalMux I__17991 (
            .O(N__78900),
            .I(N__78894));
    LocalMux I__17990 (
            .O(N__78897),
            .I(\pid_side.error_d_reg_prevZ0Z_2 ));
    Odrv4 I__17989 (
            .O(N__78894),
            .I(\pid_side.error_d_reg_prevZ0Z_2 ));
    CascadeMux I__17988 (
            .O(N__78889),
            .I(N__78886));
    InMux I__17987 (
            .O(N__78886),
            .I(N__78880));
    InMux I__17986 (
            .O(N__78885),
            .I(N__78880));
    LocalMux I__17985 (
            .O(N__78880),
            .I(\pid_side.error_d_reg_prevZ0Z_3 ));
    InMux I__17984 (
            .O(N__78877),
            .I(N__78871));
    InMux I__17983 (
            .O(N__78876),
            .I(N__78871));
    LocalMux I__17982 (
            .O(N__78871),
            .I(\pid_side.error_p_regZ0Z_3 ));
    InMux I__17981 (
            .O(N__78868),
            .I(N__78865));
    LocalMux I__17980 (
            .O(N__78865),
            .I(\pid_front.N_27_0_i_i_0 ));
    CascadeMux I__17979 (
            .O(N__78862),
            .I(\pid_front.N_426_cascade_ ));
    InMux I__17978 (
            .O(N__78859),
            .I(N__78856));
    LocalMux I__17977 (
            .O(N__78856),
            .I(N__78853));
    Span4Mux_h I__17976 (
            .O(N__78853),
            .I(N__78850));
    Odrv4 I__17975 (
            .O(N__78850),
            .I(\pid_front.error_cry_2_c_RNIKGVOZ0Z2 ));
    CascadeMux I__17974 (
            .O(N__78847),
            .I(\pid_front.m7_2_01_cascade_ ));
    InMux I__17973 (
            .O(N__78844),
            .I(N__78841));
    LocalMux I__17972 (
            .O(N__78841),
            .I(N__78838));
    Span4Mux_h I__17971 (
            .O(N__78838),
            .I(N__78835));
    Odrv4 I__17970 (
            .O(N__78835),
            .I(\pid_front.error_i_reg_esr_RNO_5Z0Z_19 ));
    InMux I__17969 (
            .O(N__78832),
            .I(N__78829));
    LocalMux I__17968 (
            .O(N__78829),
            .I(\pid_front.error_i_reg_esr_RNO_2_0_19 ));
    InMux I__17967 (
            .O(N__78826),
            .I(N__78823));
    LocalMux I__17966 (
            .O(N__78823),
            .I(\pid_front.error_i_reg_esr_RNO_3Z0Z_19 ));
    InMux I__17965 (
            .O(N__78820),
            .I(N__78817));
    LocalMux I__17964 (
            .O(N__78817),
            .I(N__78814));
    Span12Mux_h I__17963 (
            .O(N__78814),
            .I(N__78811));
    Odrv12 I__17962 (
            .O(N__78811),
            .I(\pid_front.O_11 ));
    InMux I__17961 (
            .O(N__78808),
            .I(N__78800));
    InMux I__17960 (
            .O(N__78807),
            .I(N__78800));
    InMux I__17959 (
            .O(N__78806),
            .I(N__78797));
    InMux I__17958 (
            .O(N__78805),
            .I(N__78794));
    LocalMux I__17957 (
            .O(N__78800),
            .I(N__78791));
    LocalMux I__17956 (
            .O(N__78797),
            .I(N__78786));
    LocalMux I__17955 (
            .O(N__78794),
            .I(N__78786));
    Span4Mux_v I__17954 (
            .O(N__78791),
            .I(N__78781));
    Span4Mux_h I__17953 (
            .O(N__78786),
            .I(N__78781));
    Odrv4 I__17952 (
            .O(N__78781),
            .I(\pid_front.error_d_regZ0Z_8 ));
    InMux I__17951 (
            .O(N__78778),
            .I(N__78775));
    LocalMux I__17950 (
            .O(N__78775),
            .I(N__78772));
    Odrv12 I__17949 (
            .O(N__78772),
            .I(\pid_front.O_6 ));
    InMux I__17948 (
            .O(N__78769),
            .I(N__78760));
    InMux I__17947 (
            .O(N__78768),
            .I(N__78760));
    InMux I__17946 (
            .O(N__78767),
            .I(N__78760));
    LocalMux I__17945 (
            .O(N__78760),
            .I(N__78757));
    Span4Mux_h I__17944 (
            .O(N__78757),
            .I(N__78754));
    Span4Mux_h I__17943 (
            .O(N__78754),
            .I(N__78751));
    Odrv4 I__17942 (
            .O(N__78751),
            .I(\pid_front.error_d_regZ0Z_3 ));
    InMux I__17941 (
            .O(N__78748),
            .I(N__78745));
    LocalMux I__17940 (
            .O(N__78745),
            .I(N__78742));
    Odrv12 I__17939 (
            .O(N__78742),
            .I(\pid_front.O_12 ));
    InMux I__17938 (
            .O(N__78739),
            .I(N__78733));
    InMux I__17937 (
            .O(N__78738),
            .I(N__78728));
    InMux I__17936 (
            .O(N__78737),
            .I(N__78728));
    CascadeMux I__17935 (
            .O(N__78736),
            .I(N__78724));
    LocalMux I__17934 (
            .O(N__78733),
            .I(N__78719));
    LocalMux I__17933 (
            .O(N__78728),
            .I(N__78719));
    InMux I__17932 (
            .O(N__78727),
            .I(N__78714));
    InMux I__17931 (
            .O(N__78724),
            .I(N__78714));
    Span4Mux_v I__17930 (
            .O(N__78719),
            .I(N__78711));
    LocalMux I__17929 (
            .O(N__78714),
            .I(N__78708));
    Odrv4 I__17928 (
            .O(N__78711),
            .I(\pid_front.error_d_regZ0Z_9 ));
    Odrv12 I__17927 (
            .O(N__78708),
            .I(\pid_front.error_d_regZ0Z_9 ));
    InMux I__17926 (
            .O(N__78703),
            .I(N__78699));
    InMux I__17925 (
            .O(N__78702),
            .I(N__78696));
    LocalMux I__17924 (
            .O(N__78699),
            .I(N__78691));
    LocalMux I__17923 (
            .O(N__78696),
            .I(N__78686));
    CascadeMux I__17922 (
            .O(N__78695),
            .I(N__78683));
    InMux I__17921 (
            .O(N__78694),
            .I(N__78679));
    Span4Mux_h I__17920 (
            .O(N__78691),
            .I(N__78676));
    InMux I__17919 (
            .O(N__78690),
            .I(N__78673));
    InMux I__17918 (
            .O(N__78689),
            .I(N__78670));
    Span4Mux_h I__17917 (
            .O(N__78686),
            .I(N__78667));
    InMux I__17916 (
            .O(N__78683),
            .I(N__78662));
    InMux I__17915 (
            .O(N__78682),
            .I(N__78662));
    LocalMux I__17914 (
            .O(N__78679),
            .I(\pid_front.error_d_reg_prevZ0Z_12 ));
    Odrv4 I__17913 (
            .O(N__78676),
            .I(\pid_front.error_d_reg_prevZ0Z_12 ));
    LocalMux I__17912 (
            .O(N__78673),
            .I(\pid_front.error_d_reg_prevZ0Z_12 ));
    LocalMux I__17911 (
            .O(N__78670),
            .I(\pid_front.error_d_reg_prevZ0Z_12 ));
    Odrv4 I__17910 (
            .O(N__78667),
            .I(\pid_front.error_d_reg_prevZ0Z_12 ));
    LocalMux I__17909 (
            .O(N__78662),
            .I(\pid_front.error_d_reg_prevZ0Z_12 ));
    CascadeMux I__17908 (
            .O(N__78649),
            .I(N__78646));
    InMux I__17907 (
            .O(N__78646),
            .I(N__78643));
    LocalMux I__17906 (
            .O(N__78643),
            .I(N__78640));
    Span4Mux_h I__17905 (
            .O(N__78640),
            .I(N__78637));
    Odrv4 I__17904 (
            .O(N__78637),
            .I(\pid_front.N_5_0_0 ));
    InMux I__17903 (
            .O(N__78634),
            .I(N__78631));
    LocalMux I__17902 (
            .O(N__78631),
            .I(N__78628));
    Span12Mux_v I__17901 (
            .O(N__78628),
            .I(N__78625));
    Odrv12 I__17900 (
            .O(N__78625),
            .I(\pid_side.O_1_8 ));
    InMux I__17899 (
            .O(N__78622),
            .I(N__78618));
    InMux I__17898 (
            .O(N__78621),
            .I(N__78615));
    LocalMux I__17897 (
            .O(N__78618),
            .I(N__78608));
    LocalMux I__17896 (
            .O(N__78615),
            .I(N__78608));
    InMux I__17895 (
            .O(N__78614),
            .I(N__78603));
    InMux I__17894 (
            .O(N__78613),
            .I(N__78600));
    Span4Mux_v I__17893 (
            .O(N__78608),
            .I(N__78597));
    InMux I__17892 (
            .O(N__78607),
            .I(N__78594));
    InMux I__17891 (
            .O(N__78606),
            .I(N__78591));
    LocalMux I__17890 (
            .O(N__78603),
            .I(N__78588));
    LocalMux I__17889 (
            .O(N__78600),
            .I(N__78585));
    Odrv4 I__17888 (
            .O(N__78597),
            .I(\pid_side.error_d_regZ0Z_5 ));
    LocalMux I__17887 (
            .O(N__78594),
            .I(\pid_side.error_d_regZ0Z_5 ));
    LocalMux I__17886 (
            .O(N__78591),
            .I(\pid_side.error_d_regZ0Z_5 ));
    Odrv4 I__17885 (
            .O(N__78588),
            .I(\pid_side.error_d_regZ0Z_5 ));
    Odrv4 I__17884 (
            .O(N__78585),
            .I(\pid_side.error_d_regZ0Z_5 ));
    InMux I__17883 (
            .O(N__78574),
            .I(N__78571));
    LocalMux I__17882 (
            .O(N__78571),
            .I(N__78568));
    Span4Mux_v I__17881 (
            .O(N__78568),
            .I(N__78565));
    Span4Mux_v I__17880 (
            .O(N__78565),
            .I(N__78562));
    Span4Mux_h I__17879 (
            .O(N__78562),
            .I(N__78559));
    Odrv4 I__17878 (
            .O(N__78559),
            .I(\pid_side.O_1_9 ));
    InMux I__17877 (
            .O(N__78556),
            .I(N__78544));
    InMux I__17876 (
            .O(N__78555),
            .I(N__78544));
    InMux I__17875 (
            .O(N__78554),
            .I(N__78544));
    InMux I__17874 (
            .O(N__78553),
            .I(N__78544));
    LocalMux I__17873 (
            .O(N__78544),
            .I(N__78539));
    InMux I__17872 (
            .O(N__78543),
            .I(N__78536));
    InMux I__17871 (
            .O(N__78542),
            .I(N__78533));
    Span4Mux_h I__17870 (
            .O(N__78539),
            .I(N__78530));
    LocalMux I__17869 (
            .O(N__78536),
            .I(N__78527));
    LocalMux I__17868 (
            .O(N__78533),
            .I(N__78524));
    Odrv4 I__17867 (
            .O(N__78530),
            .I(\pid_side.error_d_regZ0Z_6 ));
    Odrv4 I__17866 (
            .O(N__78527),
            .I(\pid_side.error_d_regZ0Z_6 ));
    Odrv4 I__17865 (
            .O(N__78524),
            .I(\pid_side.error_d_regZ0Z_6 ));
    CascadeMux I__17864 (
            .O(N__78517),
            .I(\pid_side.m9_2_03_3_i_0_o2_0_cascade_ ));
    InMux I__17863 (
            .O(N__78514),
            .I(N__78511));
    LocalMux I__17862 (
            .O(N__78511),
            .I(N__78507));
    InMux I__17861 (
            .O(N__78510),
            .I(N__78504));
    Span4Mux_v I__17860 (
            .O(N__78507),
            .I(N__78491));
    LocalMux I__17859 (
            .O(N__78504),
            .I(N__78491));
    InMux I__17858 (
            .O(N__78503),
            .I(N__78488));
    InMux I__17857 (
            .O(N__78502),
            .I(N__78485));
    InMux I__17856 (
            .O(N__78501),
            .I(N__78482));
    InMux I__17855 (
            .O(N__78500),
            .I(N__78477));
    InMux I__17854 (
            .O(N__78499),
            .I(N__78477));
    InMux I__17853 (
            .O(N__78498),
            .I(N__78474));
    InMux I__17852 (
            .O(N__78497),
            .I(N__78469));
    InMux I__17851 (
            .O(N__78496),
            .I(N__78469));
    Span4Mux_v I__17850 (
            .O(N__78491),
            .I(N__78465));
    LocalMux I__17849 (
            .O(N__78488),
            .I(N__78460));
    LocalMux I__17848 (
            .O(N__78485),
            .I(N__78460));
    LocalMux I__17847 (
            .O(N__78482),
            .I(N__78453));
    LocalMux I__17846 (
            .O(N__78477),
            .I(N__78453));
    LocalMux I__17845 (
            .O(N__78474),
            .I(N__78453));
    LocalMux I__17844 (
            .O(N__78469),
            .I(N__78450));
    InMux I__17843 (
            .O(N__78468),
            .I(N__78447));
    Span4Mux_h I__17842 (
            .O(N__78465),
            .I(N__78440));
    Span4Mux_v I__17841 (
            .O(N__78460),
            .I(N__78440));
    Span4Mux_v I__17840 (
            .O(N__78453),
            .I(N__78440));
    Span12Mux_s10_h I__17839 (
            .O(N__78450),
            .I(N__78436));
    LocalMux I__17838 (
            .O(N__78447),
            .I(N__78433));
    Sp12to4 I__17837 (
            .O(N__78440),
            .I(N__78430));
    InMux I__17836 (
            .O(N__78439),
            .I(N__78427));
    Odrv12 I__17835 (
            .O(N__78436),
            .I(xy_ki_fast_3));
    Odrv4 I__17834 (
            .O(N__78433),
            .I(xy_ki_fast_3));
    Odrv12 I__17833 (
            .O(N__78430),
            .I(xy_ki_fast_3));
    LocalMux I__17832 (
            .O(N__78427),
            .I(xy_ki_fast_3));
    InMux I__17831 (
            .O(N__78418),
            .I(N__78414));
    InMux I__17830 (
            .O(N__78417),
            .I(N__78409));
    LocalMux I__17829 (
            .O(N__78414),
            .I(N__78406));
    InMux I__17828 (
            .O(N__78413),
            .I(N__78403));
    InMux I__17827 (
            .O(N__78412),
            .I(N__78400));
    LocalMux I__17826 (
            .O(N__78409),
            .I(N__78397));
    Span4Mux_s0_h I__17825 (
            .O(N__78406),
            .I(N__78392));
    LocalMux I__17824 (
            .O(N__78403),
            .I(N__78388));
    LocalMux I__17823 (
            .O(N__78400),
            .I(N__78383));
    Span4Mux_h I__17822 (
            .O(N__78397),
            .I(N__78383));
    InMux I__17821 (
            .O(N__78396),
            .I(N__78380));
    CascadeMux I__17820 (
            .O(N__78395),
            .I(N__78377));
    Span4Mux_v I__17819 (
            .O(N__78392),
            .I(N__78373));
    InMux I__17818 (
            .O(N__78391),
            .I(N__78370));
    Span4Mux_v I__17817 (
            .O(N__78388),
            .I(N__78367));
    Span4Mux_h I__17816 (
            .O(N__78383),
            .I(N__78362));
    LocalMux I__17815 (
            .O(N__78380),
            .I(N__78362));
    InMux I__17814 (
            .O(N__78377),
            .I(N__78357));
    InMux I__17813 (
            .O(N__78376),
            .I(N__78357));
    Sp12to4 I__17812 (
            .O(N__78373),
            .I(N__78354));
    LocalMux I__17811 (
            .O(N__78370),
            .I(N__78351));
    Span4Mux_h I__17810 (
            .O(N__78367),
            .I(N__78348));
    Span4Mux_h I__17809 (
            .O(N__78362),
            .I(N__78345));
    LocalMux I__17808 (
            .O(N__78357),
            .I(N__78342));
    Span12Mux_h I__17807 (
            .O(N__78354),
            .I(N__78337));
    Span12Mux_h I__17806 (
            .O(N__78351),
            .I(N__78337));
    Odrv4 I__17805 (
            .O(N__78348),
            .I(\pid_front.error_10 ));
    Odrv4 I__17804 (
            .O(N__78345),
            .I(\pid_front.error_10 ));
    Odrv12 I__17803 (
            .O(N__78342),
            .I(\pid_front.error_10 ));
    Odrv12 I__17802 (
            .O(N__78337),
            .I(\pid_front.error_10 ));
    CascadeMux I__17801 (
            .O(N__78328),
            .I(\pid_front.error_i_reg_esr_RNO_6_0_12_cascade_ ));
    InMux I__17800 (
            .O(N__78325),
            .I(N__78320));
    InMux I__17799 (
            .O(N__78324),
            .I(N__78316));
    InMux I__17798 (
            .O(N__78323),
            .I(N__78313));
    LocalMux I__17797 (
            .O(N__78320),
            .I(N__78308));
    InMux I__17796 (
            .O(N__78319),
            .I(N__78301));
    LocalMux I__17795 (
            .O(N__78316),
            .I(N__78298));
    LocalMux I__17794 (
            .O(N__78313),
            .I(N__78295));
    InMux I__17793 (
            .O(N__78312),
            .I(N__78290));
    InMux I__17792 (
            .O(N__78311),
            .I(N__78290));
    Span4Mux_h I__17791 (
            .O(N__78308),
            .I(N__78287));
    InMux I__17790 (
            .O(N__78307),
            .I(N__78282));
    InMux I__17789 (
            .O(N__78306),
            .I(N__78282));
    InMux I__17788 (
            .O(N__78305),
            .I(N__78276));
    InMux I__17787 (
            .O(N__78304),
            .I(N__78276));
    LocalMux I__17786 (
            .O(N__78301),
            .I(N__78271));
    Span4Mux_h I__17785 (
            .O(N__78298),
            .I(N__78268));
    Span4Mux_h I__17784 (
            .O(N__78295),
            .I(N__78263));
    LocalMux I__17783 (
            .O(N__78290),
            .I(N__78263));
    Span4Mux_h I__17782 (
            .O(N__78287),
            .I(N__78260));
    LocalMux I__17781 (
            .O(N__78282),
            .I(N__78257));
    InMux I__17780 (
            .O(N__78281),
            .I(N__78254));
    LocalMux I__17779 (
            .O(N__78276),
            .I(N__78251));
    InMux I__17778 (
            .O(N__78275),
            .I(N__78246));
    InMux I__17777 (
            .O(N__78274),
            .I(N__78246));
    Span12Mux_s1_h I__17776 (
            .O(N__78271),
            .I(N__78243));
    Span4Mux_h I__17775 (
            .O(N__78268),
            .I(N__78240));
    Span4Mux_h I__17774 (
            .O(N__78263),
            .I(N__78237));
    Span4Mux_v I__17773 (
            .O(N__78260),
            .I(N__78234));
    Span4Mux_v I__17772 (
            .O(N__78257),
            .I(N__78231));
    LocalMux I__17771 (
            .O(N__78254),
            .I(N__78224));
    Span4Mux_v I__17770 (
            .O(N__78251),
            .I(N__78224));
    LocalMux I__17769 (
            .O(N__78246),
            .I(N__78224));
    Span12Mux_h I__17768 (
            .O(N__78243),
            .I(N__78221));
    Span4Mux_h I__17767 (
            .O(N__78240),
            .I(N__78218));
    Odrv4 I__17766 (
            .O(N__78237),
            .I(\pid_front.error_14 ));
    Odrv4 I__17765 (
            .O(N__78234),
            .I(\pid_front.error_14 ));
    Odrv4 I__17764 (
            .O(N__78231),
            .I(\pid_front.error_14 ));
    Odrv4 I__17763 (
            .O(N__78224),
            .I(\pid_front.error_14 ));
    Odrv12 I__17762 (
            .O(N__78221),
            .I(\pid_front.error_14 ));
    Odrv4 I__17761 (
            .O(N__78218),
            .I(\pid_front.error_14 ));
    InMux I__17760 (
            .O(N__78205),
            .I(N__78202));
    LocalMux I__17759 (
            .O(N__78202),
            .I(N__78199));
    Span4Mux_h I__17758 (
            .O(N__78199),
            .I(N__78196));
    Odrv4 I__17757 (
            .O(N__78196),
            .I(\pid_front.N_228_0 ));
    InMux I__17756 (
            .O(N__78193),
            .I(N__78190));
    LocalMux I__17755 (
            .O(N__78190),
            .I(\pid_side.un4_error_i_reg_31_bm_sx ));
    InMux I__17754 (
            .O(N__78187),
            .I(N__78184));
    LocalMux I__17753 (
            .O(N__78184),
            .I(N__78181));
    Odrv4 I__17752 (
            .O(N__78181),
            .I(\pid_front.error_i_reg_esr_RNO_4Z0Z_19 ));
    InMux I__17751 (
            .O(N__78178),
            .I(N__78175));
    LocalMux I__17750 (
            .O(N__78175),
            .I(N__78172));
    Span4Mux_h I__17749 (
            .O(N__78172),
            .I(N__78169));
    Odrv4 I__17748 (
            .O(N__78169),
            .I(\pid_front.error_i_reg_esr_RNO_0Z0Z_19 ));
    CascadeMux I__17747 (
            .O(N__78166),
            .I(\pid_front.error_i_reg_esr_RNO_1_0_19_cascade_ ));
    InMux I__17746 (
            .O(N__78163),
            .I(N__78160));
    LocalMux I__17745 (
            .O(N__78160),
            .I(N__78157));
    Span4Mux_h I__17744 (
            .O(N__78157),
            .I(N__78154));
    Span4Mux_h I__17743 (
            .O(N__78154),
            .I(N__78151));
    Odrv4 I__17742 (
            .O(N__78151),
            .I(\pid_front.error_i_regZ0Z_19 ));
    CEMux I__17741 (
            .O(N__78148),
            .I(N__78143));
    CEMux I__17740 (
            .O(N__78147),
            .I(N__78138));
    CEMux I__17739 (
            .O(N__78146),
            .I(N__78132));
    LocalMux I__17738 (
            .O(N__78143),
            .I(N__78126));
    CEMux I__17737 (
            .O(N__78142),
            .I(N__78123));
    CEMux I__17736 (
            .O(N__78141),
            .I(N__78120));
    LocalMux I__17735 (
            .O(N__78138),
            .I(N__78117));
    CEMux I__17734 (
            .O(N__78137),
            .I(N__78114));
    CEMux I__17733 (
            .O(N__78136),
            .I(N__78111));
    CEMux I__17732 (
            .O(N__78135),
            .I(N__78107));
    LocalMux I__17731 (
            .O(N__78132),
            .I(N__78102));
    CEMux I__17730 (
            .O(N__78131),
            .I(N__78099));
    CEMux I__17729 (
            .O(N__78130),
            .I(N__78096));
    CEMux I__17728 (
            .O(N__78129),
            .I(N__78093));
    Span4Mux_h I__17727 (
            .O(N__78126),
            .I(N__78088));
    LocalMux I__17726 (
            .O(N__78123),
            .I(N__78088));
    LocalMux I__17725 (
            .O(N__78120),
            .I(N__78085));
    Span4Mux_v I__17724 (
            .O(N__78117),
            .I(N__78080));
    LocalMux I__17723 (
            .O(N__78114),
            .I(N__78080));
    LocalMux I__17722 (
            .O(N__78111),
            .I(N__78077));
    CEMux I__17721 (
            .O(N__78110),
            .I(N__78074));
    LocalMux I__17720 (
            .O(N__78107),
            .I(N__78071));
    CEMux I__17719 (
            .O(N__78106),
            .I(N__78067));
    CEMux I__17718 (
            .O(N__78105),
            .I(N__78064));
    Span4Mux_h I__17717 (
            .O(N__78102),
            .I(N__78059));
    LocalMux I__17716 (
            .O(N__78099),
            .I(N__78059));
    LocalMux I__17715 (
            .O(N__78096),
            .I(N__78054));
    LocalMux I__17714 (
            .O(N__78093),
            .I(N__78054));
    Span4Mux_h I__17713 (
            .O(N__78088),
            .I(N__78051));
    Span4Mux_v I__17712 (
            .O(N__78085),
            .I(N__78048));
    Span4Mux_h I__17711 (
            .O(N__78080),
            .I(N__78043));
    Span4Mux_h I__17710 (
            .O(N__78077),
            .I(N__78043));
    LocalMux I__17709 (
            .O(N__78074),
            .I(N__78038));
    Span4Mux_h I__17708 (
            .O(N__78071),
            .I(N__78038));
    CEMux I__17707 (
            .O(N__78070),
            .I(N__78035));
    LocalMux I__17706 (
            .O(N__78067),
            .I(N__78030));
    LocalMux I__17705 (
            .O(N__78064),
            .I(N__78030));
    Span4Mux_h I__17704 (
            .O(N__78059),
            .I(N__78027));
    Span4Mux_h I__17703 (
            .O(N__78054),
            .I(N__78022));
    Span4Mux_h I__17702 (
            .O(N__78051),
            .I(N__78022));
    Span4Mux_h I__17701 (
            .O(N__78048),
            .I(N__78015));
    Span4Mux_h I__17700 (
            .O(N__78043),
            .I(N__78015));
    Span4Mux_h I__17699 (
            .O(N__78038),
            .I(N__78015));
    LocalMux I__17698 (
            .O(N__78035),
            .I(N__78011));
    Span4Mux_v I__17697 (
            .O(N__78030),
            .I(N__78006));
    Span4Mux_h I__17696 (
            .O(N__78027),
            .I(N__78006));
    Sp12to4 I__17695 (
            .O(N__78022),
            .I(N__78001));
    Sp12to4 I__17694 (
            .O(N__78015),
            .I(N__78001));
    CEMux I__17693 (
            .O(N__78014),
            .I(N__77998));
    Span4Mux_h I__17692 (
            .O(N__78011),
            .I(N__77993));
    Span4Mux_v I__17691 (
            .O(N__78006),
            .I(N__77993));
    Span12Mux_v I__17690 (
            .O(N__78001),
            .I(N__77990));
    LocalMux I__17689 (
            .O(N__77998),
            .I(\pid_front.state_ns_0_0 ));
    Odrv4 I__17688 (
            .O(N__77993),
            .I(\pid_front.state_ns_0_0 ));
    Odrv12 I__17687 (
            .O(N__77990),
            .I(\pid_front.state_ns_0_0 ));
    InMux I__17686 (
            .O(N__77983),
            .I(N__77978));
    InMux I__17685 (
            .O(N__77982),
            .I(N__77975));
    InMux I__17684 (
            .O(N__77981),
            .I(N__77969));
    LocalMux I__17683 (
            .O(N__77978),
            .I(N__77963));
    LocalMux I__17682 (
            .O(N__77975),
            .I(N__77960));
    InMux I__17681 (
            .O(N__77974),
            .I(N__77956));
    InMux I__17680 (
            .O(N__77973),
            .I(N__77953));
    InMux I__17679 (
            .O(N__77972),
            .I(N__77950));
    LocalMux I__17678 (
            .O(N__77969),
            .I(N__77947));
    InMux I__17677 (
            .O(N__77968),
            .I(N__77944));
    InMux I__17676 (
            .O(N__77967),
            .I(N__77939));
    InMux I__17675 (
            .O(N__77966),
            .I(N__77939));
    Span4Mux_v I__17674 (
            .O(N__77963),
            .I(N__77936));
    Span4Mux_h I__17673 (
            .O(N__77960),
            .I(N__77933));
    InMux I__17672 (
            .O(N__77959),
            .I(N__77930));
    LocalMux I__17671 (
            .O(N__77956),
            .I(N__77927));
    LocalMux I__17670 (
            .O(N__77953),
            .I(N__77924));
    LocalMux I__17669 (
            .O(N__77950),
            .I(N__77921));
    Span4Mux_v I__17668 (
            .O(N__77947),
            .I(N__77914));
    LocalMux I__17667 (
            .O(N__77944),
            .I(N__77914));
    LocalMux I__17666 (
            .O(N__77939),
            .I(N__77914));
    Span4Mux_v I__17665 (
            .O(N__77936),
            .I(N__77911));
    Span4Mux_h I__17664 (
            .O(N__77933),
            .I(N__77908));
    LocalMux I__17663 (
            .O(N__77930),
            .I(N__77905));
    Span4Mux_v I__17662 (
            .O(N__77927),
            .I(N__77902));
    Span4Mux_v I__17661 (
            .O(N__77924),
            .I(N__77895));
    Span4Mux_v I__17660 (
            .O(N__77921),
            .I(N__77895));
    Span4Mux_h I__17659 (
            .O(N__77914),
            .I(N__77895));
    Sp12to4 I__17658 (
            .O(N__77911),
            .I(N__77892));
    Span4Mux_h I__17657 (
            .O(N__77908),
            .I(N__77889));
    Span4Mux_v I__17656 (
            .O(N__77905),
            .I(N__77884));
    Span4Mux_h I__17655 (
            .O(N__77902),
            .I(N__77884));
    Span4Mux_h I__17654 (
            .O(N__77895),
            .I(N__77881));
    Odrv12 I__17653 (
            .O(N__77892),
            .I(\pid_front.error_5 ));
    Odrv4 I__17652 (
            .O(N__77889),
            .I(\pid_front.error_5 ));
    Odrv4 I__17651 (
            .O(N__77884),
            .I(\pid_front.error_5 ));
    Odrv4 I__17650 (
            .O(N__77881),
            .I(\pid_front.error_5 ));
    InMux I__17649 (
            .O(N__77872),
            .I(N__77868));
    InMux I__17648 (
            .O(N__77871),
            .I(N__77864));
    LocalMux I__17647 (
            .O(N__77868),
            .I(N__77861));
    InMux I__17646 (
            .O(N__77867),
            .I(N__77858));
    LocalMux I__17645 (
            .O(N__77864),
            .I(N__77850));
    Span4Mux_v I__17644 (
            .O(N__77861),
            .I(N__77845));
    LocalMux I__17643 (
            .O(N__77858),
            .I(N__77842));
    InMux I__17642 (
            .O(N__77857),
            .I(N__77839));
    InMux I__17641 (
            .O(N__77856),
            .I(N__77836));
    InMux I__17640 (
            .O(N__77855),
            .I(N__77831));
    InMux I__17639 (
            .O(N__77854),
            .I(N__77831));
    InMux I__17638 (
            .O(N__77853),
            .I(N__77828));
    Span4Mux_h I__17637 (
            .O(N__77850),
            .I(N__77825));
    InMux I__17636 (
            .O(N__77849),
            .I(N__77820));
    InMux I__17635 (
            .O(N__77848),
            .I(N__77820));
    Span4Mux_h I__17634 (
            .O(N__77845),
            .I(N__77817));
    Span4Mux_v I__17633 (
            .O(N__77842),
            .I(N__77814));
    LocalMux I__17632 (
            .O(N__77839),
            .I(N__77811));
    LocalMux I__17631 (
            .O(N__77836),
            .I(N__77807));
    LocalMux I__17630 (
            .O(N__77831),
            .I(N__77804));
    LocalMux I__17629 (
            .O(N__77828),
            .I(N__77801));
    Span4Mux_h I__17628 (
            .O(N__77825),
            .I(N__77796));
    LocalMux I__17627 (
            .O(N__77820),
            .I(N__77796));
    Span4Mux_v I__17626 (
            .O(N__77817),
            .I(N__77793));
    Sp12to4 I__17625 (
            .O(N__77814),
            .I(N__77790));
    Span4Mux_v I__17624 (
            .O(N__77811),
            .I(N__77787));
    InMux I__17623 (
            .O(N__77810),
            .I(N__77784));
    Span4Mux_h I__17622 (
            .O(N__77807),
            .I(N__77777));
    Span4Mux_h I__17621 (
            .O(N__77804),
            .I(N__77777));
    Span4Mux_h I__17620 (
            .O(N__77801),
            .I(N__77772));
    Span4Mux_h I__17619 (
            .O(N__77796),
            .I(N__77772));
    Sp12to4 I__17618 (
            .O(N__77793),
            .I(N__77763));
    Span12Mux_s10_h I__17617 (
            .O(N__77790),
            .I(N__77763));
    Sp12to4 I__17616 (
            .O(N__77787),
            .I(N__77763));
    LocalMux I__17615 (
            .O(N__77784),
            .I(N__77763));
    InMux I__17614 (
            .O(N__77783),
            .I(N__77758));
    InMux I__17613 (
            .O(N__77782),
            .I(N__77758));
    Odrv4 I__17612 (
            .O(N__77777),
            .I(\pid_front.error_6 ));
    Odrv4 I__17611 (
            .O(N__77772),
            .I(\pid_front.error_6 ));
    Odrv12 I__17610 (
            .O(N__77763),
            .I(\pid_front.error_6 ));
    LocalMux I__17609 (
            .O(N__77758),
            .I(\pid_front.error_6 ));
    InMux I__17608 (
            .O(N__77749),
            .I(N__77744));
    InMux I__17607 (
            .O(N__77748),
            .I(N__77740));
    InMux I__17606 (
            .O(N__77747),
            .I(N__77736));
    LocalMux I__17605 (
            .O(N__77744),
            .I(N__77733));
    InMux I__17604 (
            .O(N__77743),
            .I(N__77729));
    LocalMux I__17603 (
            .O(N__77740),
            .I(N__77726));
    InMux I__17602 (
            .O(N__77739),
            .I(N__77723));
    LocalMux I__17601 (
            .O(N__77736),
            .I(N__77719));
    Span4Mux_h I__17600 (
            .O(N__77733),
            .I(N__77716));
    InMux I__17599 (
            .O(N__77732),
            .I(N__77713));
    LocalMux I__17598 (
            .O(N__77729),
            .I(N__77710));
    Span4Mux_h I__17597 (
            .O(N__77726),
            .I(N__77705));
    LocalMux I__17596 (
            .O(N__77723),
            .I(N__77705));
    InMux I__17595 (
            .O(N__77722),
            .I(N__77702));
    Span12Mux_s1_h I__17594 (
            .O(N__77719),
            .I(N__77699));
    Span4Mux_h I__17593 (
            .O(N__77716),
            .I(N__77696));
    LocalMux I__17592 (
            .O(N__77713),
            .I(N__77691));
    Span4Mux_h I__17591 (
            .O(N__77710),
            .I(N__77691));
    Span4Mux_h I__17590 (
            .O(N__77705),
            .I(N__77688));
    LocalMux I__17589 (
            .O(N__77702),
            .I(N__77685));
    Span12Mux_h I__17588 (
            .O(N__77699),
            .I(N__77680));
    Span4Mux_h I__17587 (
            .O(N__77696),
            .I(N__77675));
    Span4Mux_h I__17586 (
            .O(N__77691),
            .I(N__77675));
    Span4Mux_h I__17585 (
            .O(N__77688),
            .I(N__77670));
    Span4Mux_h I__17584 (
            .O(N__77685),
            .I(N__77670));
    InMux I__17583 (
            .O(N__77684),
            .I(N__77665));
    InMux I__17582 (
            .O(N__77683),
            .I(N__77665));
    Odrv12 I__17581 (
            .O(N__77680),
            .I(\pid_front.error_7 ));
    Odrv4 I__17580 (
            .O(N__77675),
            .I(\pid_front.error_7 ));
    Odrv4 I__17579 (
            .O(N__77670),
            .I(\pid_front.error_7 ));
    LocalMux I__17578 (
            .O(N__77665),
            .I(\pid_front.error_7 ));
    CascadeMux I__17577 (
            .O(N__77656),
            .I(\pid_side.error_i_reg_esr_RNO_4Z0Z_22_cascade_ ));
    InMux I__17576 (
            .O(N__77653),
            .I(N__77650));
    LocalMux I__17575 (
            .O(N__77650),
            .I(\pid_side.error_i_reg_esr_RNO_3Z0Z_22 ));
    CascadeMux I__17574 (
            .O(N__77647),
            .I(\pid_side.N_297_cascade_ ));
    InMux I__17573 (
            .O(N__77644),
            .I(N__77641));
    LocalMux I__17572 (
            .O(N__77641),
            .I(N__77638));
    Span4Mux_h I__17571 (
            .O(N__77638),
            .I(N__77635));
    Odrv4 I__17570 (
            .O(N__77635),
            .I(\pid_side.N_301 ));
    InMux I__17569 (
            .O(N__77632),
            .I(N__77629));
    LocalMux I__17568 (
            .O(N__77629),
            .I(\pid_side.N_252 ));
    CascadeMux I__17567 (
            .O(N__77626),
            .I(\pid_side.N_252_cascade_ ));
    InMux I__17566 (
            .O(N__77623),
            .I(N__77619));
    InMux I__17565 (
            .O(N__77622),
            .I(N__77616));
    LocalMux I__17564 (
            .O(N__77619),
            .I(N__77613));
    LocalMux I__17563 (
            .O(N__77616),
            .I(N__77609));
    Span4Mux_v I__17562 (
            .O(N__77613),
            .I(N__77606));
    InMux I__17561 (
            .O(N__77612),
            .I(N__77602));
    Span4Mux_h I__17560 (
            .O(N__77609),
            .I(N__77597));
    Span4Mux_h I__17559 (
            .O(N__77606),
            .I(N__77597));
    InMux I__17558 (
            .O(N__77605),
            .I(N__77594));
    LocalMux I__17557 (
            .O(N__77602),
            .I(\pid_side.m1_0_03 ));
    Odrv4 I__17556 (
            .O(N__77597),
            .I(\pid_side.m1_0_03 ));
    LocalMux I__17555 (
            .O(N__77594),
            .I(\pid_side.m1_0_03 ));
    CascadeMux I__17554 (
            .O(N__77587),
            .I(\pid_side.N_537_cascade_ ));
    InMux I__17553 (
            .O(N__77584),
            .I(N__77581));
    LocalMux I__17552 (
            .O(N__77581),
            .I(N__77578));
    Span4Mux_h I__17551 (
            .O(N__77578),
            .I(N__77575));
    Span4Mux_v I__17550 (
            .O(N__77575),
            .I(N__77571));
    InMux I__17549 (
            .O(N__77574),
            .I(N__77568));
    Odrv4 I__17548 (
            .O(N__77571),
            .I(\pid_side.N_189 ));
    LocalMux I__17547 (
            .O(N__77568),
            .I(\pid_side.N_189 ));
    InMux I__17546 (
            .O(N__77563),
            .I(N__77560));
    LocalMux I__17545 (
            .O(N__77560),
            .I(N__77557));
    Span4Mux_h I__17544 (
            .O(N__77557),
            .I(N__77554));
    Span4Mux_h I__17543 (
            .O(N__77554),
            .I(N__77551));
    Odrv4 I__17542 (
            .O(N__77551),
            .I(drone_H_disp_side_i_8));
    InMux I__17541 (
            .O(N__77548),
            .I(bfn_20_16_0_));
    InMux I__17540 (
            .O(N__77545),
            .I(N__77542));
    LocalMux I__17539 (
            .O(N__77542),
            .I(N__77539));
    Span4Mux_h I__17538 (
            .O(N__77539),
            .I(N__77536));
    Span4Mux_h I__17537 (
            .O(N__77536),
            .I(N__77533));
    Odrv4 I__17536 (
            .O(N__77533),
            .I(drone_H_disp_side_i_9));
    InMux I__17535 (
            .O(N__77530),
            .I(\pid_side.error_cry_4 ));
    InMux I__17534 (
            .O(N__77527),
            .I(N__77524));
    LocalMux I__17533 (
            .O(N__77524),
            .I(N__77521));
    Odrv12 I__17532 (
            .O(N__77521),
            .I(drone_H_disp_side_i_10));
    InMux I__17531 (
            .O(N__77518),
            .I(\pid_side.error_cry_5 ));
    InMux I__17530 (
            .O(N__77515),
            .I(N__77512));
    LocalMux I__17529 (
            .O(N__77512),
            .I(N__77509));
    Span4Mux_h I__17528 (
            .O(N__77509),
            .I(N__77506));
    Span4Mux_h I__17527 (
            .O(N__77506),
            .I(N__77503));
    Odrv4 I__17526 (
            .O(N__77503),
            .I(\pid_side.error_axbZ0Z_7 ));
    InMux I__17525 (
            .O(N__77500),
            .I(\pid_side.error_cry_6 ));
    InMux I__17524 (
            .O(N__77497),
            .I(N__77494));
    LocalMux I__17523 (
            .O(N__77494),
            .I(N__77491));
    Span4Mux_h I__17522 (
            .O(N__77491),
            .I(N__77488));
    Span4Mux_h I__17521 (
            .O(N__77488),
            .I(N__77485));
    Odrv4 I__17520 (
            .O(N__77485),
            .I(\pid_side.error_axb_8_l_ofxZ0 ));
    CascadeMux I__17519 (
            .O(N__77482),
            .I(N__77478));
    InMux I__17518 (
            .O(N__77481),
            .I(N__77475));
    InMux I__17517 (
            .O(N__77478),
            .I(N__77472));
    LocalMux I__17516 (
            .O(N__77475),
            .I(N__77469));
    LocalMux I__17515 (
            .O(N__77472),
            .I(N__77466));
    Span4Mux_v I__17514 (
            .O(N__77469),
            .I(N__77462));
    Span12Mux_s8_h I__17513 (
            .O(N__77466),
            .I(N__77459));
    InMux I__17512 (
            .O(N__77465),
            .I(N__77456));
    Odrv4 I__17511 (
            .O(N__77462),
            .I(drone_H_disp_side_12));
    Odrv12 I__17510 (
            .O(N__77459),
            .I(drone_H_disp_side_12));
    LocalMux I__17509 (
            .O(N__77456),
            .I(drone_H_disp_side_12));
    InMux I__17508 (
            .O(N__77449),
            .I(\pid_side.error_cry_7 ));
    InMux I__17507 (
            .O(N__77446),
            .I(N__77443));
    LocalMux I__17506 (
            .O(N__77443),
            .I(N__77440));
    Odrv12 I__17505 (
            .O(N__77440),
            .I(drone_H_disp_side_i_12));
    CascadeMux I__17504 (
            .O(N__77437),
            .I(N__77434));
    InMux I__17503 (
            .O(N__77434),
            .I(N__77431));
    LocalMux I__17502 (
            .O(N__77431),
            .I(N__77428));
    Span4Mux_h I__17501 (
            .O(N__77428),
            .I(N__77424));
    InMux I__17500 (
            .O(N__77427),
            .I(N__77421));
    Span4Mux_h I__17499 (
            .O(N__77424),
            .I(N__77416));
    LocalMux I__17498 (
            .O(N__77421),
            .I(N__77416));
    Odrv4 I__17497 (
            .O(N__77416),
            .I(drone_H_disp_side_13));
    InMux I__17496 (
            .O(N__77413),
            .I(\pid_side.error_cry_8 ));
    InMux I__17495 (
            .O(N__77410),
            .I(N__77407));
    LocalMux I__17494 (
            .O(N__77407),
            .I(N__77404));
    Odrv12 I__17493 (
            .O(N__77404),
            .I(drone_H_disp_side_i_13));
    InMux I__17492 (
            .O(N__77401),
            .I(\pid_side.error_cry_9 ));
    InMux I__17491 (
            .O(N__77398),
            .I(N__77395));
    LocalMux I__17490 (
            .O(N__77395),
            .I(N__77392));
    Sp12to4 I__17489 (
            .O(N__77392),
            .I(N__77389));
    Odrv12 I__17488 (
            .O(N__77389),
            .I(drone_H_disp_side_15));
    CascadeMux I__17487 (
            .O(N__77386),
            .I(N__77382));
    InMux I__17486 (
            .O(N__77385),
            .I(N__77377));
    InMux I__17485 (
            .O(N__77382),
            .I(N__77377));
    LocalMux I__17484 (
            .O(N__77377),
            .I(N__77374));
    Odrv12 I__17483 (
            .O(N__77374),
            .I(drone_H_disp_side_14));
    InMux I__17482 (
            .O(N__77371),
            .I(\pid_side.error_cry_10 ));
    InMux I__17481 (
            .O(N__77368),
            .I(N__77364));
    InMux I__17480 (
            .O(N__77367),
            .I(N__77361));
    LocalMux I__17479 (
            .O(N__77364),
            .I(N__77358));
    LocalMux I__17478 (
            .O(N__77361),
            .I(N__77355));
    Span4Mux_v I__17477 (
            .O(N__77358),
            .I(N__77352));
    Span4Mux_v I__17476 (
            .O(N__77355),
            .I(N__77347));
    Span4Mux_h I__17475 (
            .O(N__77352),
            .I(N__77347));
    Odrv4 I__17474 (
            .O(N__77347),
            .I(\pid_side.N_224 ));
    InMux I__17473 (
            .O(N__77344),
            .I(N__77341));
    LocalMux I__17472 (
            .O(N__77341),
            .I(N__77338));
    Span4Mux_v I__17471 (
            .O(N__77338),
            .I(N__77335));
    Odrv4 I__17470 (
            .O(N__77335),
            .I(\pid_side.m19_2_03_0_1 ));
    InMux I__17469 (
            .O(N__77332),
            .I(N__77329));
    LocalMux I__17468 (
            .O(N__77329),
            .I(N__77326));
    Span4Mux_h I__17467 (
            .O(N__77326),
            .I(N__77323));
    Span4Mux_h I__17466 (
            .O(N__77323),
            .I(N__77320));
    Odrv4 I__17465 (
            .O(N__77320),
            .I(dron_frame_decoder_1_source_H_disp_side_fast_0));
    CascadeMux I__17464 (
            .O(N__77317),
            .I(N__77314));
    InMux I__17463 (
            .O(N__77314),
            .I(N__77311));
    LocalMux I__17462 (
            .O(N__77311),
            .I(\pid_side.error_axb_0 ));
    CascadeMux I__17461 (
            .O(N__77308),
            .I(N__77305));
    InMux I__17460 (
            .O(N__77305),
            .I(N__77302));
    LocalMux I__17459 (
            .O(N__77302),
            .I(N__77299));
    Span4Mux_v I__17458 (
            .O(N__77299),
            .I(N__77296));
    Span4Mux_h I__17457 (
            .O(N__77296),
            .I(N__77293));
    Odrv4 I__17456 (
            .O(N__77293),
            .I(\pid_side.error_axbZ0Z_1 ));
    InMux I__17455 (
            .O(N__77290),
            .I(\pid_side.error_cry_0 ));
    CascadeMux I__17454 (
            .O(N__77287),
            .I(N__77284));
    InMux I__17453 (
            .O(N__77284),
            .I(N__77281));
    LocalMux I__17452 (
            .O(N__77281),
            .I(N__77278));
    Span4Mux_v I__17451 (
            .O(N__77278),
            .I(N__77275));
    Span4Mux_h I__17450 (
            .O(N__77275),
            .I(N__77272));
    Odrv4 I__17449 (
            .O(N__77272),
            .I(\pid_side.error_axbZ0Z_2 ));
    InMux I__17448 (
            .O(N__77269),
            .I(\pid_side.error_cry_1 ));
    InMux I__17447 (
            .O(N__77266),
            .I(N__77263));
    LocalMux I__17446 (
            .O(N__77263),
            .I(N__77260));
    Span4Mux_v I__17445 (
            .O(N__77260),
            .I(N__77257));
    Span4Mux_h I__17444 (
            .O(N__77257),
            .I(N__77254));
    Odrv4 I__17443 (
            .O(N__77254),
            .I(\pid_side.error_axbZ0Z_3 ));
    InMux I__17442 (
            .O(N__77251),
            .I(\pid_side.error_cry_2 ));
    InMux I__17441 (
            .O(N__77248),
            .I(N__77245));
    LocalMux I__17440 (
            .O(N__77245),
            .I(N__77242));
    Span4Mux_h I__17439 (
            .O(N__77242),
            .I(N__77239));
    Span4Mux_h I__17438 (
            .O(N__77239),
            .I(N__77236));
    Odrv4 I__17437 (
            .O(N__77236),
            .I(drone_H_disp_side_i_4));
    InMux I__17436 (
            .O(N__77233),
            .I(N__77228));
    InMux I__17435 (
            .O(N__77232),
            .I(N__77225));
    InMux I__17434 (
            .O(N__77231),
            .I(N__77219));
    LocalMux I__17433 (
            .O(N__77228),
            .I(N__77215));
    LocalMux I__17432 (
            .O(N__77225),
            .I(N__77212));
    InMux I__17431 (
            .O(N__77224),
            .I(N__77207));
    InMux I__17430 (
            .O(N__77223),
            .I(N__77207));
    InMux I__17429 (
            .O(N__77222),
            .I(N__77204));
    LocalMux I__17428 (
            .O(N__77219),
            .I(N__77201));
    InMux I__17427 (
            .O(N__77218),
            .I(N__77198));
    Span4Mux_v I__17426 (
            .O(N__77215),
            .I(N__77195));
    Span4Mux_s0_h I__17425 (
            .O(N__77212),
            .I(N__77192));
    LocalMux I__17424 (
            .O(N__77207),
            .I(N__77189));
    LocalMux I__17423 (
            .O(N__77204),
            .I(N__77182));
    Span4Mux_v I__17422 (
            .O(N__77201),
            .I(N__77182));
    LocalMux I__17421 (
            .O(N__77198),
            .I(N__77182));
    Span4Mux_h I__17420 (
            .O(N__77195),
            .I(N__77177));
    Span4Mux_h I__17419 (
            .O(N__77192),
            .I(N__77177));
    Span4Mux_v I__17418 (
            .O(N__77189),
            .I(N__77174));
    Span4Mux_h I__17417 (
            .O(N__77182),
            .I(N__77171));
    Odrv4 I__17416 (
            .O(N__77177),
            .I(\pid_side.error_4 ));
    Odrv4 I__17415 (
            .O(N__77174),
            .I(\pid_side.error_4 ));
    Odrv4 I__17414 (
            .O(N__77171),
            .I(\pid_side.error_4 ));
    InMux I__17413 (
            .O(N__77164),
            .I(\pid_side.error_cry_3 ));
    InMux I__17412 (
            .O(N__77161),
            .I(N__77158));
    LocalMux I__17411 (
            .O(N__77158),
            .I(N__77155));
    Span4Mux_h I__17410 (
            .O(N__77155),
            .I(N__77152));
    Span4Mux_h I__17409 (
            .O(N__77152),
            .I(N__77149));
    Odrv4 I__17408 (
            .O(N__77149),
            .I(drone_H_disp_side_i_5));
    InMux I__17407 (
            .O(N__77146),
            .I(\pid_side.error_cry_0_0 ));
    InMux I__17406 (
            .O(N__77143),
            .I(N__77140));
    LocalMux I__17405 (
            .O(N__77140),
            .I(N__77137));
    Span4Mux_h I__17404 (
            .O(N__77137),
            .I(N__77134));
    Span4Mux_h I__17403 (
            .O(N__77134),
            .I(N__77131));
    Odrv4 I__17402 (
            .O(N__77131),
            .I(drone_H_disp_side_i_6));
    InMux I__17401 (
            .O(N__77128),
            .I(\pid_side.error_cry_1_0 ));
    InMux I__17400 (
            .O(N__77125),
            .I(N__77122));
    LocalMux I__17399 (
            .O(N__77122),
            .I(N__77119));
    Odrv12 I__17398 (
            .O(N__77119),
            .I(drone_H_disp_side_i_7));
    InMux I__17397 (
            .O(N__77116),
            .I(\pid_side.error_cry_2_0 ));
    CascadeMux I__17396 (
            .O(N__77113),
            .I(\pid_side.N_224_cascade_ ));
    InMux I__17395 (
            .O(N__77110),
            .I(N__77107));
    LocalMux I__17394 (
            .O(N__77107),
            .I(\pid_side.N_258 ));
    InMux I__17393 (
            .O(N__77104),
            .I(N__77101));
    LocalMux I__17392 (
            .O(N__77101),
            .I(N__77098));
    Odrv4 I__17391 (
            .O(N__77098),
            .I(\pid_side.m17_2_03_4_0 ));
    CascadeMux I__17390 (
            .O(N__77095),
            .I(pid_side_N_491_cascade_));
    CascadeMux I__17389 (
            .O(N__77092),
            .I(\pid_front.m21_2_03_0_1_1_cascade_ ));
    InMux I__17388 (
            .O(N__77089),
            .I(N__77085));
    InMux I__17387 (
            .O(N__77088),
            .I(N__77080));
    LocalMux I__17386 (
            .O(N__77085),
            .I(N__77076));
    InMux I__17385 (
            .O(N__77084),
            .I(N__77073));
    InMux I__17384 (
            .O(N__77083),
            .I(N__77070));
    LocalMux I__17383 (
            .O(N__77080),
            .I(N__77067));
    InMux I__17382 (
            .O(N__77079),
            .I(N__77064));
    Span4Mux_v I__17381 (
            .O(N__77076),
            .I(N__77059));
    LocalMux I__17380 (
            .O(N__77073),
            .I(N__77059));
    LocalMux I__17379 (
            .O(N__77070),
            .I(N__77054));
    Span4Mux_h I__17378 (
            .O(N__77067),
            .I(N__77054));
    LocalMux I__17377 (
            .O(N__77064),
            .I(\pid_front.N_163 ));
    Odrv4 I__17376 (
            .O(N__77059),
            .I(\pid_front.N_163 ));
    Odrv4 I__17375 (
            .O(N__77054),
            .I(\pid_front.N_163 ));
    InMux I__17374 (
            .O(N__77047),
            .I(N__77044));
    LocalMux I__17373 (
            .O(N__77044),
            .I(N__77041));
    Span4Mux_v I__17372 (
            .O(N__77041),
            .I(N__77038));
    Odrv4 I__17371 (
            .O(N__77038),
            .I(\pid_front.m21_2_03_0_1 ));
    CascadeMux I__17370 (
            .O(N__77035),
            .I(\pid_side.m78_0_m2_1_ns_1_cascade_ ));
    CascadeMux I__17369 (
            .O(N__77032),
            .I(\pid_side.N_184_cascade_ ));
    InMux I__17368 (
            .O(N__77029),
            .I(N__77025));
    InMux I__17367 (
            .O(N__77028),
            .I(N__77022));
    LocalMux I__17366 (
            .O(N__77025),
            .I(N__77017));
    LocalMux I__17365 (
            .O(N__77022),
            .I(N__77017));
    Span4Mux_v I__17364 (
            .O(N__77017),
            .I(N__77014));
    Odrv4 I__17363 (
            .O(N__77014),
            .I(\pid_side.N_229 ));
    InMux I__17362 (
            .O(N__77011),
            .I(N__77008));
    LocalMux I__17361 (
            .O(N__77008),
            .I(N__77005));
    Span4Mux_h I__17360 (
            .O(N__77005),
            .I(N__77002));
    Odrv4 I__17359 (
            .O(N__77002),
            .I(\pid_side.N_437 ));
    InMux I__17358 (
            .O(N__76999),
            .I(N__76996));
    LocalMux I__17357 (
            .O(N__76996),
            .I(\pid_side.N_245 ));
    CascadeMux I__17356 (
            .O(N__76993),
            .I(\pid_side.N_245_cascade_ ));
    InMux I__17355 (
            .O(N__76990),
            .I(N__76987));
    LocalMux I__17354 (
            .O(N__76987),
            .I(N__76984));
    Odrv4 I__17353 (
            .O(N__76984),
            .I(\pid_side.N_262 ));
    CascadeMux I__17352 (
            .O(N__76981),
            .I(N__76978));
    InMux I__17351 (
            .O(N__76978),
            .I(N__76975));
    LocalMux I__17350 (
            .O(N__76975),
            .I(N__76972));
    Span4Mux_v I__17349 (
            .O(N__76972),
            .I(N__76969));
    Span4Mux_h I__17348 (
            .O(N__76969),
            .I(N__76966));
    Odrv4 I__17347 (
            .O(N__76966),
            .I(pid_side_N_306));
    InMux I__17346 (
            .O(N__76963),
            .I(N__76960));
    LocalMux I__17345 (
            .O(N__76960),
            .I(N__76957));
    Span4Mux_v I__17344 (
            .O(N__76957),
            .I(N__76951));
    InMux I__17343 (
            .O(N__76956),
            .I(N__76948));
    InMux I__17342 (
            .O(N__76955),
            .I(N__76945));
    InMux I__17341 (
            .O(N__76954),
            .I(N__76942));
    Span4Mux_h I__17340 (
            .O(N__76951),
            .I(N__76939));
    LocalMux I__17339 (
            .O(N__76948),
            .I(N__76936));
    LocalMux I__17338 (
            .O(N__76945),
            .I(N__76933));
    LocalMux I__17337 (
            .O(N__76942),
            .I(N__76930));
    Span4Mux_h I__17336 (
            .O(N__76939),
            .I(N__76927));
    Span4Mux_v I__17335 (
            .O(N__76936),
            .I(N__76920));
    Span4Mux_h I__17334 (
            .O(N__76933),
            .I(N__76920));
    Span4Mux_v I__17333 (
            .O(N__76930),
            .I(N__76920));
    Odrv4 I__17332 (
            .O(N__76927),
            .I(pid_front_N_474_1));
    Odrv4 I__17331 (
            .O(N__76920),
            .I(pid_front_N_474_1));
    CascadeMux I__17330 (
            .O(N__76915),
            .I(pid_side_N_306_cascade_));
    InMux I__17329 (
            .O(N__76912),
            .I(N__76909));
    LocalMux I__17328 (
            .O(N__76909),
            .I(N__76906));
    Span4Mux_v I__17327 (
            .O(N__76906),
            .I(N__76903));
    Odrv4 I__17326 (
            .O(N__76903),
            .I(\pid_side.m27_2_03_0_0 ));
    InMux I__17325 (
            .O(N__76900),
            .I(N__76897));
    LocalMux I__17324 (
            .O(N__76897),
            .I(N__76892));
    InMux I__17323 (
            .O(N__76896),
            .I(N__76889));
    InMux I__17322 (
            .O(N__76895),
            .I(N__76886));
    Span4Mux_h I__17321 (
            .O(N__76892),
            .I(N__76881));
    LocalMux I__17320 (
            .O(N__76889),
            .I(N__76881));
    LocalMux I__17319 (
            .O(N__76886),
            .I(N__76878));
    Span4Mux_v I__17318 (
            .O(N__76881),
            .I(N__76870));
    Span4Mux_v I__17317 (
            .O(N__76878),
            .I(N__76870));
    InMux I__17316 (
            .O(N__76877),
            .I(N__76861));
    InMux I__17315 (
            .O(N__76876),
            .I(N__76856));
    InMux I__17314 (
            .O(N__76875),
            .I(N__76856));
    Span4Mux_h I__17313 (
            .O(N__76870),
            .I(N__76852));
    InMux I__17312 (
            .O(N__76869),
            .I(N__76849));
    CascadeMux I__17311 (
            .O(N__76868),
            .I(N__76846));
    InMux I__17310 (
            .O(N__76867),
            .I(N__76843));
    InMux I__17309 (
            .O(N__76866),
            .I(N__76840));
    InMux I__17308 (
            .O(N__76865),
            .I(N__76837));
    InMux I__17307 (
            .O(N__76864),
            .I(N__76834));
    LocalMux I__17306 (
            .O(N__76861),
            .I(N__76829));
    LocalMux I__17305 (
            .O(N__76856),
            .I(N__76829));
    InMux I__17304 (
            .O(N__76855),
            .I(N__76826));
    Span4Mux_h I__17303 (
            .O(N__76852),
            .I(N__76821));
    LocalMux I__17302 (
            .O(N__76849),
            .I(N__76821));
    InMux I__17301 (
            .O(N__76846),
            .I(N__76817));
    LocalMux I__17300 (
            .O(N__76843),
            .I(N__76814));
    LocalMux I__17299 (
            .O(N__76840),
            .I(N__76805));
    LocalMux I__17298 (
            .O(N__76837),
            .I(N__76805));
    LocalMux I__17297 (
            .O(N__76834),
            .I(N__76805));
    Span4Mux_v I__17296 (
            .O(N__76829),
            .I(N__76805));
    LocalMux I__17295 (
            .O(N__76826),
            .I(N__76802));
    Span4Mux_v I__17294 (
            .O(N__76821),
            .I(N__76799));
    InMux I__17293 (
            .O(N__76820),
            .I(N__76796));
    LocalMux I__17292 (
            .O(N__76817),
            .I(N__76793));
    Span4Mux_v I__17291 (
            .O(N__76814),
            .I(N__76790));
    Span4Mux_v I__17290 (
            .O(N__76805),
            .I(N__76787));
    Sp12to4 I__17289 (
            .O(N__76802),
            .I(N__76780));
    Sp12to4 I__17288 (
            .O(N__76799),
            .I(N__76780));
    LocalMux I__17287 (
            .O(N__76796),
            .I(N__76780));
    Span4Mux_v I__17286 (
            .O(N__76793),
            .I(N__76773));
    Span4Mux_v I__17285 (
            .O(N__76790),
            .I(N__76773));
    Span4Mux_h I__17284 (
            .O(N__76787),
            .I(N__76773));
    Span12Mux_s9_h I__17283 (
            .O(N__76780),
            .I(N__76770));
    Odrv4 I__17282 (
            .O(N__76773),
            .I(pid_side_N_492));
    Odrv12 I__17281 (
            .O(N__76770),
            .I(pid_side_N_492));
    CascadeMux I__17280 (
            .O(N__76765),
            .I(\pid_side.error_i_reg_esr_RNO_5Z0Z_14_cascade_ ));
    InMux I__17279 (
            .O(N__76762),
            .I(N__76759));
    LocalMux I__17278 (
            .O(N__76759),
            .I(N__76756));
    Odrv12 I__17277 (
            .O(N__76756),
            .I(\pid_side.error_i_reg_esr_RNO_4Z0Z_14 ));
    InMux I__17276 (
            .O(N__76753),
            .I(N__76750));
    LocalMux I__17275 (
            .O(N__76750),
            .I(\pid_side.N_160 ));
    CascadeMux I__17274 (
            .O(N__76747),
            .I(\pid_side.N_160_cascade_ ));
    CascadeMux I__17273 (
            .O(N__76744),
            .I(\pid_side.error_d_reg_prev_esr_RNIBGIE2Z0Z_1_cascade_ ));
    InMux I__17272 (
            .O(N__76741),
            .I(N__76738));
    LocalMux I__17271 (
            .O(N__76738),
            .I(\pid_side.error_p_reg_esr_RNIIQL11_0Z0Z_1 ));
    InMux I__17270 (
            .O(N__76735),
            .I(N__76729));
    InMux I__17269 (
            .O(N__76734),
            .I(N__76729));
    LocalMux I__17268 (
            .O(N__76729),
            .I(N__76726));
    Span12Mux_s10_v I__17267 (
            .O(N__76726),
            .I(N__76721));
    InMux I__17266 (
            .O(N__76725),
            .I(N__76716));
    InMux I__17265 (
            .O(N__76724),
            .I(N__76716));
    Odrv12 I__17264 (
            .O(N__76721),
            .I(\pid_side.error_d_reg_prevZ0Z_0 ));
    LocalMux I__17263 (
            .O(N__76716),
            .I(\pid_side.error_d_reg_prevZ0Z_0 ));
    InMux I__17262 (
            .O(N__76711),
            .I(N__76705));
    InMux I__17261 (
            .O(N__76710),
            .I(N__76705));
    LocalMux I__17260 (
            .O(N__76705),
            .I(\pid_side.error_p_reg_esr_RNICBEQ_0Z0Z_2 ));
    CascadeMux I__17259 (
            .O(N__76702),
            .I(N__76699));
    InMux I__17258 (
            .O(N__76699),
            .I(N__76695));
    CascadeMux I__17257 (
            .O(N__76698),
            .I(N__76692));
    LocalMux I__17256 (
            .O(N__76695),
            .I(N__76689));
    InMux I__17255 (
            .O(N__76692),
            .I(N__76686));
    Span4Mux_v I__17254 (
            .O(N__76689),
            .I(N__76683));
    LocalMux I__17253 (
            .O(N__76686),
            .I(N__76680));
    Span4Mux_v I__17252 (
            .O(N__76683),
            .I(N__76675));
    Span4Mux_h I__17251 (
            .O(N__76680),
            .I(N__76675));
    Span4Mux_v I__17250 (
            .O(N__76675),
            .I(N__76672));
    Odrv4 I__17249 (
            .O(N__76672),
            .I(pid_side_error_i_reg_9_sn_rn_1_15));
    CascadeMux I__17248 (
            .O(N__76669),
            .I(\pid_side.error_i_reg_9_sn_rn_0_15_cascade_ ));
    InMux I__17247 (
            .O(N__76666),
            .I(N__76663));
    LocalMux I__17246 (
            .O(N__76663),
            .I(N__76660));
    Odrv12 I__17245 (
            .O(N__76660),
            .I(\pid_side.error_i_reg_9_sn_sn_15 ));
    InMux I__17244 (
            .O(N__76657),
            .I(N__76652));
    InMux I__17243 (
            .O(N__76656),
            .I(N__76649));
    InMux I__17242 (
            .O(N__76655),
            .I(N__76644));
    LocalMux I__17241 (
            .O(N__76652),
            .I(N__76641));
    LocalMux I__17240 (
            .O(N__76649),
            .I(N__76638));
    InMux I__17239 (
            .O(N__76648),
            .I(N__76635));
    InMux I__17238 (
            .O(N__76647),
            .I(N__76632));
    LocalMux I__17237 (
            .O(N__76644),
            .I(N__76629));
    Odrv4 I__17236 (
            .O(N__76641),
            .I(\pid_side.N_161 ));
    Odrv4 I__17235 (
            .O(N__76638),
            .I(\pid_side.N_161 ));
    LocalMux I__17234 (
            .O(N__76635),
            .I(\pid_side.N_161 ));
    LocalMux I__17233 (
            .O(N__76632),
            .I(\pid_side.N_161 ));
    Odrv12 I__17232 (
            .O(N__76629),
            .I(\pid_side.N_161 ));
    CascadeMux I__17231 (
            .O(N__76618),
            .I(\pid_side.N_258_cascade_ ));
    InMux I__17230 (
            .O(N__76615),
            .I(N__76612));
    LocalMux I__17229 (
            .O(N__76612),
            .I(N__76609));
    Span4Mux_h I__17228 (
            .O(N__76609),
            .I(N__76606));
    Span4Mux_v I__17227 (
            .O(N__76606),
            .I(N__76603));
    Span4Mux_h I__17226 (
            .O(N__76603),
            .I(N__76600));
    Odrv4 I__17225 (
            .O(N__76600),
            .I(\pid_side.error_i_reg_9_rn_1_15 ));
    CascadeMux I__17224 (
            .O(N__76597),
            .I(\pid_side.m19_2_03_0_0_cascade_ ));
    InMux I__17223 (
            .O(N__76594),
            .I(N__76591));
    LocalMux I__17222 (
            .O(N__76591),
            .I(\pid_side.error_i_reg_9_sn_15 ));
    CascadeMux I__17221 (
            .O(N__76588),
            .I(N__76585));
    InMux I__17220 (
            .O(N__76585),
            .I(N__76582));
    LocalMux I__17219 (
            .O(N__76582),
            .I(N__76579));
    Span4Mux_v I__17218 (
            .O(N__76579),
            .I(N__76576));
    Span4Mux_h I__17217 (
            .O(N__76576),
            .I(N__76573));
    Odrv4 I__17216 (
            .O(N__76573),
            .I(\pid_side.error_i_regZ0Z_15 ));
    InMux I__17215 (
            .O(N__76570),
            .I(N__76567));
    LocalMux I__17214 (
            .O(N__76567),
            .I(N__76564));
    Span4Mux_h I__17213 (
            .O(N__76564),
            .I(N__76561));
    Span4Mux_v I__17212 (
            .O(N__76561),
            .I(N__76558));
    Odrv4 I__17211 (
            .O(N__76558),
            .I(\pid_side.g1_2_1 ));
    CascadeMux I__17210 (
            .O(N__76555),
            .I(\pid_side.g0_3_2_cascade_ ));
    InMux I__17209 (
            .O(N__76552),
            .I(N__76548));
    InMux I__17208 (
            .O(N__76551),
            .I(N__76545));
    LocalMux I__17207 (
            .O(N__76548),
            .I(N__76542));
    LocalMux I__17206 (
            .O(N__76545),
            .I(N__76539));
    Span4Mux_h I__17205 (
            .O(N__76542),
            .I(N__76536));
    Span4Mux_v I__17204 (
            .O(N__76539),
            .I(N__76530));
    Span4Mux_h I__17203 (
            .O(N__76536),
            .I(N__76530));
    InMux I__17202 (
            .O(N__76535),
            .I(N__76527));
    Odrv4 I__17201 (
            .O(N__76530),
            .I(\pid_side.error_i_reg_esr_RNIO6NRZ0Z_14 ));
    LocalMux I__17200 (
            .O(N__76527),
            .I(\pid_side.error_i_reg_esr_RNIO6NRZ0Z_14 ));
    CascadeMux I__17199 (
            .O(N__76522),
            .I(\pid_side.g1_3_cascade_ ));
    InMux I__17198 (
            .O(N__76519),
            .I(N__76516));
    LocalMux I__17197 (
            .O(N__76516),
            .I(N__76513));
    Span4Mux_v I__17196 (
            .O(N__76513),
            .I(N__76507));
    InMux I__17195 (
            .O(N__76512),
            .I(N__76504));
    InMux I__17194 (
            .O(N__76511),
            .I(N__76499));
    InMux I__17193 (
            .O(N__76510),
            .I(N__76499));
    Span4Mux_h I__17192 (
            .O(N__76507),
            .I(N__76494));
    LocalMux I__17191 (
            .O(N__76504),
            .I(N__76494));
    LocalMux I__17190 (
            .O(N__76499),
            .I(N__76491));
    Odrv4 I__17189 (
            .O(N__76494),
            .I(\pid_side.error_i_reg_esr_RNIM3MRZ0Z_13 ));
    Odrv4 I__17188 (
            .O(N__76491),
            .I(\pid_side.error_i_reg_esr_RNIM3MRZ0Z_13 ));
    CascadeMux I__17187 (
            .O(N__76486),
            .I(N__76482));
    InMux I__17186 (
            .O(N__76485),
            .I(N__76479));
    InMux I__17185 (
            .O(N__76482),
            .I(N__76476));
    LocalMux I__17184 (
            .O(N__76479),
            .I(N__76471));
    LocalMux I__17183 (
            .O(N__76476),
            .I(N__76471));
    Span4Mux_h I__17182 (
            .O(N__76471),
            .I(N__76468));
    Odrv4 I__17181 (
            .O(N__76468),
            .I(\pid_side.error_p_reg_esr_RNI46CB9Z0Z_12 ));
    CascadeMux I__17180 (
            .O(N__76465),
            .I(\pid_side.N_2608_0_cascade_ ));
    InMux I__17179 (
            .O(N__76462),
            .I(N__76459));
    LocalMux I__17178 (
            .O(N__76459),
            .I(N__76456));
    Odrv12 I__17177 (
            .O(N__76456),
            .I(\pid_side.g0_2 ));
    CascadeMux I__17176 (
            .O(N__76453),
            .I(N__76450));
    InMux I__17175 (
            .O(N__76450),
            .I(N__76446));
    CascadeMux I__17174 (
            .O(N__76449),
            .I(N__76443));
    LocalMux I__17173 (
            .O(N__76446),
            .I(N__76440));
    InMux I__17172 (
            .O(N__76443),
            .I(N__76436));
    Span4Mux_v I__17171 (
            .O(N__76440),
            .I(N__76433));
    InMux I__17170 (
            .O(N__76439),
            .I(N__76430));
    LocalMux I__17169 (
            .O(N__76436),
            .I(N__76427));
    Span4Mux_h I__17168 (
            .O(N__76433),
            .I(N__76424));
    LocalMux I__17167 (
            .O(N__76430),
            .I(N__76419));
    Span4Mux_h I__17166 (
            .O(N__76427),
            .I(N__76419));
    Odrv4 I__17165 (
            .O(N__76424),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_1_c_RNI0LLN ));
    Odrv4 I__17164 (
            .O(N__76419),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_1_c_RNI0LLN ));
    InMux I__17163 (
            .O(N__76414),
            .I(N__76411));
    LocalMux I__17162 (
            .O(N__76411),
            .I(N__76408));
    Span4Mux_h I__17161 (
            .O(N__76408),
            .I(N__76405));
    Span4Mux_v I__17160 (
            .O(N__76405),
            .I(N__76402));
    Odrv4 I__17159 (
            .O(N__76402),
            .I(\pid_side.error_d_reg_prev_esr_RNI905J4Z0Z_1 ));
    CascadeMux I__17158 (
            .O(N__76399),
            .I(\pid_side.error_p_reg_esr_RNIIQL11Z0Z_1_cascade_ ));
    InMux I__17157 (
            .O(N__76396),
            .I(N__76393));
    LocalMux I__17156 (
            .O(N__76393),
            .I(\pid_side.error_d_reg_prev_esr_RNIBGIE2Z0Z_1 ));
    CascadeMux I__17155 (
            .O(N__76390),
            .I(\pid_side.error_p_reg_esr_RNIG7MC2_0Z0Z_5_cascade_ ));
    CascadeMux I__17154 (
            .O(N__76387),
            .I(N__76384));
    InMux I__17153 (
            .O(N__76384),
            .I(N__76381));
    LocalMux I__17152 (
            .O(N__76381),
            .I(N__76378));
    Span4Mux_h I__17151 (
            .O(N__76378),
            .I(N__76375));
    Odrv4 I__17150 (
            .O(N__76375),
            .I(\pid_side.error_p_reg_esr_RNIN4BP4Z0Z_3 ));
    InMux I__17149 (
            .O(N__76372),
            .I(N__76366));
    InMux I__17148 (
            .O(N__76371),
            .I(N__76366));
    LocalMux I__17147 (
            .O(N__76366),
            .I(\pid_side.error_d_reg_prevZ0Z_4 ));
    InMux I__17146 (
            .O(N__76363),
            .I(N__76360));
    LocalMux I__17145 (
            .O(N__76360),
            .I(\pid_side.error_p_reg_esr_RNIIHEQ_0Z0Z_4 ));
    CascadeMux I__17144 (
            .O(N__76357),
            .I(\pid_side.error_p_reg_esr_RNIIHEQ_0Z0Z_4_cascade_ ));
    InMux I__17143 (
            .O(N__76354),
            .I(N__76349));
    InMux I__17142 (
            .O(N__76353),
            .I(N__76344));
    InMux I__17141 (
            .O(N__76352),
            .I(N__76344));
    LocalMux I__17140 (
            .O(N__76349),
            .I(N__76341));
    LocalMux I__17139 (
            .O(N__76344),
            .I(N__76338));
    Odrv4 I__17138 (
            .O(N__76341),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_3_c_RNI6TNN ));
    Odrv12 I__17137 (
            .O(N__76338),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_3_c_RNI6TNN ));
    InMux I__17136 (
            .O(N__76333),
            .I(N__76330));
    LocalMux I__17135 (
            .O(N__76330),
            .I(N__76327));
    Span4Mux_h I__17134 (
            .O(N__76327),
            .I(N__76324));
    Span4Mux_v I__17133 (
            .O(N__76324),
            .I(N__76321));
    Odrv4 I__17132 (
            .O(N__76321),
            .I(\pid_side.error_p_reg_esr_RNISL2L4Z0Z_3 ));
    InMux I__17131 (
            .O(N__76318),
            .I(N__76314));
    InMux I__17130 (
            .O(N__76317),
            .I(N__76311));
    LocalMux I__17129 (
            .O(N__76314),
            .I(N__76306));
    LocalMux I__17128 (
            .O(N__76311),
            .I(N__76306));
    Span4Mux_v I__17127 (
            .O(N__76306),
            .I(N__76303));
    Span4Mux_h I__17126 (
            .O(N__76303),
            .I(N__76300));
    Odrv4 I__17125 (
            .O(N__76300),
            .I(\pid_side.error_d_reg_prev_esr_RNIKAJOZ0Z_19 ));
    InMux I__17124 (
            .O(N__76297),
            .I(N__76291));
    InMux I__17123 (
            .O(N__76296),
            .I(N__76291));
    LocalMux I__17122 (
            .O(N__76291),
            .I(N__76288));
    Odrv12 I__17121 (
            .O(N__76288),
            .I(\pid_side.error_d_reg_prev_esr_RNIKAJO_0Z0Z_19 ));
    InMux I__17120 (
            .O(N__76285),
            .I(N__76280));
    InMux I__17119 (
            .O(N__76284),
            .I(N__76277));
    InMux I__17118 (
            .O(N__76283),
            .I(N__76274));
    LocalMux I__17117 (
            .O(N__76280),
            .I(N__76265));
    LocalMux I__17116 (
            .O(N__76277),
            .I(N__76265));
    LocalMux I__17115 (
            .O(N__76274),
            .I(N__76265));
    InMux I__17114 (
            .O(N__76273),
            .I(N__76262));
    InMux I__17113 (
            .O(N__76272),
            .I(N__76259));
    Span4Mux_v I__17112 (
            .O(N__76265),
            .I(N__76254));
    LocalMux I__17111 (
            .O(N__76262),
            .I(N__76254));
    LocalMux I__17110 (
            .O(N__76259),
            .I(\pid_side.error_d_reg_prevZ0Z_5 ));
    Odrv4 I__17109 (
            .O(N__76254),
            .I(\pid_side.error_d_reg_prevZ0Z_5 ));
    InMux I__17108 (
            .O(N__76249),
            .I(N__76246));
    LocalMux I__17107 (
            .O(N__76246),
            .I(N__76243));
    Span4Mux_h I__17106 (
            .O(N__76243),
            .I(N__76240));
    Odrv4 I__17105 (
            .O(N__76240),
            .I(\pid_side.error_p_reg_esr_RNI6FM11_0Z0Z_6 ));
    InMux I__17104 (
            .O(N__76237),
            .I(N__76234));
    LocalMux I__17103 (
            .O(N__76234),
            .I(\pid_side.error_d_reg_esr_RNI2OIO_3Z0Z_13 ));
    CascadeMux I__17102 (
            .O(N__76231),
            .I(\pid_side.error_d_reg_fast_esr_RNIC6BTZ0Z_12_cascade_ ));
    InMux I__17101 (
            .O(N__76228),
            .I(N__76223));
    InMux I__17100 (
            .O(N__76227),
            .I(N__76220));
    CascadeMux I__17099 (
            .O(N__76226),
            .I(N__76217));
    LocalMux I__17098 (
            .O(N__76223),
            .I(N__76213));
    LocalMux I__17097 (
            .O(N__76220),
            .I(N__76210));
    InMux I__17096 (
            .O(N__76217),
            .I(N__76205));
    InMux I__17095 (
            .O(N__76216),
            .I(N__76205));
    Span4Mux_h I__17094 (
            .O(N__76213),
            .I(N__76202));
    Span4Mux_v I__17093 (
            .O(N__76210),
            .I(N__76197));
    LocalMux I__17092 (
            .O(N__76205),
            .I(N__76197));
    Odrv4 I__17091 (
            .O(N__76202),
            .I(\pid_side.error_d_reg_prev_fastZ0Z_12 ));
    Odrv4 I__17090 (
            .O(N__76197),
            .I(\pid_side.error_d_reg_prev_fastZ0Z_12 ));
    InMux I__17089 (
            .O(N__76192),
            .I(N__76189));
    LocalMux I__17088 (
            .O(N__76189),
            .I(N__76185));
    InMux I__17087 (
            .O(N__76188),
            .I(N__76182));
    Span4Mux_v I__17086 (
            .O(N__76185),
            .I(N__76179));
    LocalMux I__17085 (
            .O(N__76182),
            .I(N__76176));
    Span4Mux_h I__17084 (
            .O(N__76179),
            .I(N__76171));
    Span4Mux_v I__17083 (
            .O(N__76176),
            .I(N__76171));
    Span4Mux_v I__17082 (
            .O(N__76171),
            .I(N__76168));
    Odrv4 I__17081 (
            .O(N__76168),
            .I(\pid_front.error_p_regZ0Z_18 ));
    InMux I__17080 (
            .O(N__76165),
            .I(N__76162));
    LocalMux I__17079 (
            .O(N__76162),
            .I(N__76159));
    Span4Mux_h I__17078 (
            .O(N__76159),
            .I(N__76155));
    InMux I__17077 (
            .O(N__76158),
            .I(N__76152));
    Odrv4 I__17076 (
            .O(N__76155),
            .I(\pid_front.error_d_reg_prevZ0Z_18 ));
    LocalMux I__17075 (
            .O(N__76152),
            .I(\pid_front.error_d_reg_prevZ0Z_18 ));
    InMux I__17074 (
            .O(N__76147),
            .I(N__76144));
    LocalMux I__17073 (
            .O(N__76144),
            .I(N__76141));
    Span12Mux_s6_v I__17072 (
            .O(N__76141),
            .I(N__76137));
    InMux I__17071 (
            .O(N__76140),
            .I(N__76134));
    Odrv12 I__17070 (
            .O(N__76137),
            .I(\pid_front.error_p_reg_esr_RNITCC61Z0Z_18 ));
    LocalMux I__17069 (
            .O(N__76134),
            .I(\pid_front.error_p_reg_esr_RNITCC61Z0Z_18 ));
    InMux I__17068 (
            .O(N__76129),
            .I(N__76126));
    LocalMux I__17067 (
            .O(N__76126),
            .I(N__76123));
    Odrv4 I__17066 (
            .O(N__76123),
            .I(\pid_side.error_p_reg_esr_RNI6FM11Z0Z_6 ));
    InMux I__17065 (
            .O(N__76120),
            .I(N__76114));
    InMux I__17064 (
            .O(N__76119),
            .I(N__76114));
    LocalMux I__17063 (
            .O(N__76114),
            .I(N__76111));
    Span4Mux_h I__17062 (
            .O(N__76111),
            .I(N__76108));
    Odrv4 I__17061 (
            .O(N__76108),
            .I(\pid_side.error_p_reg_esr_RNI76TK1Z0Z_5 ));
    InMux I__17060 (
            .O(N__76105),
            .I(N__76102));
    LocalMux I__17059 (
            .O(N__76102),
            .I(\pid_side.error_p_reg_esr_RNIIHEQZ0Z_4 ));
    CascadeMux I__17058 (
            .O(N__76099),
            .I(\pid_side.error_p_reg_esr_RNIIHEQZ0Z_4_cascade_ ));
    CascadeMux I__17057 (
            .O(N__76096),
            .I(\pid_side.error_p_reg_esr_RNI76TK1_0Z0Z_5_cascade_ ));
    CascadeMux I__17056 (
            .O(N__76093),
            .I(N__76090));
    InMux I__17055 (
            .O(N__76090),
            .I(N__76087));
    LocalMux I__17054 (
            .O(N__76087),
            .I(N__76084));
    Span4Mux_h I__17053 (
            .O(N__76084),
            .I(N__76081));
    Odrv4 I__17052 (
            .O(N__76081),
            .I(\pid_side.error_p_reg_esr_RNIG7MC2Z0Z_5 ));
    InMux I__17051 (
            .O(N__76078),
            .I(N__76075));
    LocalMux I__17050 (
            .O(N__76075),
            .I(N__76072));
    Span4Mux_h I__17049 (
            .O(N__76072),
            .I(N__76068));
    InMux I__17048 (
            .O(N__76071),
            .I(N__76065));
    Odrv4 I__17047 (
            .O(N__76068),
            .I(\pid_side.error_p_reg_esr_RNI76TK1_0Z0Z_5 ));
    LocalMux I__17046 (
            .O(N__76065),
            .I(\pid_side.error_p_reg_esr_RNI76TK1_0Z0Z_5 ));
    InMux I__17045 (
            .O(N__76060),
            .I(N__76056));
    InMux I__17044 (
            .O(N__76059),
            .I(N__76053));
    LocalMux I__17043 (
            .O(N__76056),
            .I(N__76048));
    LocalMux I__17042 (
            .O(N__76053),
            .I(N__76045));
    InMux I__17041 (
            .O(N__76052),
            .I(N__76040));
    InMux I__17040 (
            .O(N__76051),
            .I(N__76040));
    Span4Mux_v I__17039 (
            .O(N__76048),
            .I(N__76035));
    Span4Mux_v I__17038 (
            .O(N__76045),
            .I(N__76035));
    LocalMux I__17037 (
            .O(N__76040),
            .I(N__76032));
    Odrv4 I__17036 (
            .O(N__76035),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_4_c_RNI91PN ));
    Odrv12 I__17035 (
            .O(N__76032),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_4_c_RNI91PN ));
    InMux I__17034 (
            .O(N__76027),
            .I(N__76024));
    LocalMux I__17033 (
            .O(N__76024),
            .I(N__76021));
    Span4Mux_v I__17032 (
            .O(N__76021),
            .I(N__76018));
    Span4Mux_h I__17031 (
            .O(N__76018),
            .I(N__76015));
    Odrv4 I__17030 (
            .O(N__76015),
            .I(\pid_side.error_p_reg_esr_RNIG7MC2_0Z0Z_5 ));
    InMux I__17029 (
            .O(N__76012),
            .I(N__76004));
    InMux I__17028 (
            .O(N__76011),
            .I(N__76004));
    InMux I__17027 (
            .O(N__76010),
            .I(N__76001));
    InMux I__17026 (
            .O(N__76009),
            .I(N__75995));
    LocalMux I__17025 (
            .O(N__76004),
            .I(N__75990));
    LocalMux I__17024 (
            .O(N__76001),
            .I(N__75990));
    InMux I__17023 (
            .O(N__76000),
            .I(N__75983));
    InMux I__17022 (
            .O(N__75999),
            .I(N__75983));
    InMux I__17021 (
            .O(N__75998),
            .I(N__75983));
    LocalMux I__17020 (
            .O(N__75995),
            .I(N__75980));
    Span4Mux_v I__17019 (
            .O(N__75990),
            .I(N__75977));
    LocalMux I__17018 (
            .O(N__75983),
            .I(N__75972));
    Span4Mux_h I__17017 (
            .O(N__75980),
            .I(N__75972));
    Odrv4 I__17016 (
            .O(N__75977),
            .I(\pid_front.N_227 ));
    Odrv4 I__17015 (
            .O(N__75972),
            .I(\pid_front.N_227 ));
    CascadeMux I__17014 (
            .O(N__75967),
            .I(N__75959));
    InMux I__17013 (
            .O(N__75966),
            .I(N__75953));
    InMux I__17012 (
            .O(N__75965),
            .I(N__75946));
    InMux I__17011 (
            .O(N__75964),
            .I(N__75946));
    InMux I__17010 (
            .O(N__75963),
            .I(N__75946));
    CascadeMux I__17009 (
            .O(N__75962),
            .I(N__75943));
    InMux I__17008 (
            .O(N__75959),
            .I(N__75934));
    InMux I__17007 (
            .O(N__75958),
            .I(N__75934));
    CascadeMux I__17006 (
            .O(N__75957),
            .I(N__75930));
    CascadeMux I__17005 (
            .O(N__75956),
            .I(N__75927));
    LocalMux I__17004 (
            .O(N__75953),
            .I(N__75922));
    LocalMux I__17003 (
            .O(N__75946),
            .I(N__75922));
    InMux I__17002 (
            .O(N__75943),
            .I(N__75913));
    InMux I__17001 (
            .O(N__75942),
            .I(N__75913));
    InMux I__17000 (
            .O(N__75941),
            .I(N__75913));
    InMux I__16999 (
            .O(N__75940),
            .I(N__75913));
    CascadeMux I__16998 (
            .O(N__75939),
            .I(N__75910));
    LocalMux I__16997 (
            .O(N__75934),
            .I(N__75906));
    InMux I__16996 (
            .O(N__75933),
            .I(N__75903));
    InMux I__16995 (
            .O(N__75930),
            .I(N__75898));
    InMux I__16994 (
            .O(N__75927),
            .I(N__75898));
    Span4Mux_v I__16993 (
            .O(N__75922),
            .I(N__75895));
    LocalMux I__16992 (
            .O(N__75913),
            .I(N__75892));
    InMux I__16991 (
            .O(N__75910),
            .I(N__75887));
    InMux I__16990 (
            .O(N__75909),
            .I(N__75887));
    Span4Mux_h I__16989 (
            .O(N__75906),
            .I(N__75884));
    LocalMux I__16988 (
            .O(N__75903),
            .I(N__75877));
    LocalMux I__16987 (
            .O(N__75898),
            .I(N__75877));
    Sp12to4 I__16986 (
            .O(N__75895),
            .I(N__75877));
    Odrv4 I__16985 (
            .O(N__75892),
            .I(\pid_front.error_i_acumm_preregZ0Z_28 ));
    LocalMux I__16984 (
            .O(N__75887),
            .I(\pid_front.error_i_acumm_preregZ0Z_28 ));
    Odrv4 I__16983 (
            .O(N__75884),
            .I(\pid_front.error_i_acumm_preregZ0Z_28 ));
    Odrv12 I__16982 (
            .O(N__75877),
            .I(\pid_front.error_i_acumm_preregZ0Z_28 ));
    InMux I__16981 (
            .O(N__75868),
            .I(N__75862));
    InMux I__16980 (
            .O(N__75867),
            .I(N__75854));
    InMux I__16979 (
            .O(N__75866),
            .I(N__75854));
    InMux I__16978 (
            .O(N__75865),
            .I(N__75854));
    LocalMux I__16977 (
            .O(N__75862),
            .I(N__75851));
    CascadeMux I__16976 (
            .O(N__75861),
            .I(N__75846));
    LocalMux I__16975 (
            .O(N__75854),
            .I(N__75843));
    Span4Mux_h I__16974 (
            .O(N__75851),
            .I(N__75840));
    InMux I__16973 (
            .O(N__75850),
            .I(N__75837));
    InMux I__16972 (
            .O(N__75849),
            .I(N__75832));
    InMux I__16971 (
            .O(N__75846),
            .I(N__75832));
    Span4Mux_v I__16970 (
            .O(N__75843),
            .I(N__75829));
    Span4Mux_v I__16969 (
            .O(N__75840),
            .I(N__75826));
    LocalMux I__16968 (
            .O(N__75837),
            .I(N__75821));
    LocalMux I__16967 (
            .O(N__75832),
            .I(N__75821));
    Span4Mux_h I__16966 (
            .O(N__75829),
            .I(N__75818));
    Span4Mux_h I__16965 (
            .O(N__75826),
            .I(N__75813));
    Span4Mux_v I__16964 (
            .O(N__75821),
            .I(N__75813));
    Span4Mux_v I__16963 (
            .O(N__75818),
            .I(N__75810));
    Span4Mux_v I__16962 (
            .O(N__75813),
            .I(N__75807));
    Span4Mux_v I__16961 (
            .O(N__75810),
            .I(N__75804));
    Span4Mux_h I__16960 (
            .O(N__75807),
            .I(N__75801));
    Odrv4 I__16959 (
            .O(N__75804),
            .I(\pid_front.N_205 ));
    Odrv4 I__16958 (
            .O(N__75801),
            .I(\pid_front.N_205 ));
    CascadeMux I__16957 (
            .O(N__75796),
            .I(\pid_front.N_242_cascade_ ));
    InMux I__16956 (
            .O(N__75793),
            .I(N__75784));
    InMux I__16955 (
            .O(N__75792),
            .I(N__75784));
    InMux I__16954 (
            .O(N__75791),
            .I(N__75784));
    LocalMux I__16953 (
            .O(N__75784),
            .I(\pid_front.N_285 ));
    InMux I__16952 (
            .O(N__75781),
            .I(N__75778));
    LocalMux I__16951 (
            .O(N__75778),
            .I(N__75775));
    Span4Mux_h I__16950 (
            .O(N__75775),
            .I(N__75772));
    Odrv4 I__16949 (
            .O(N__75772),
            .I(\pid_front.error_i_acummZ0Z_12 ));
    CEMux I__16948 (
            .O(N__75769),
            .I(N__75761));
    CEMux I__16947 (
            .O(N__75768),
            .I(N__75758));
    CEMux I__16946 (
            .O(N__75767),
            .I(N__75755));
    CEMux I__16945 (
            .O(N__75766),
            .I(N__75752));
    CEMux I__16944 (
            .O(N__75765),
            .I(N__75749));
    CEMux I__16943 (
            .O(N__75764),
            .I(N__75746));
    LocalMux I__16942 (
            .O(N__75761),
            .I(N__75743));
    LocalMux I__16941 (
            .O(N__75758),
            .I(N__75738));
    LocalMux I__16940 (
            .O(N__75755),
            .I(N__75738));
    LocalMux I__16939 (
            .O(N__75752),
            .I(N__75735));
    LocalMux I__16938 (
            .O(N__75749),
            .I(N__75732));
    LocalMux I__16937 (
            .O(N__75746),
            .I(N__75729));
    Span4Mux_h I__16936 (
            .O(N__75743),
            .I(N__75726));
    Span4Mux_v I__16935 (
            .O(N__75738),
            .I(N__75723));
    Span4Mux_v I__16934 (
            .O(N__75735),
            .I(N__75720));
    Span4Mux_v I__16933 (
            .O(N__75732),
            .I(N__75717));
    Span4Mux_v I__16932 (
            .O(N__75729),
            .I(N__75710));
    Span4Mux_h I__16931 (
            .O(N__75726),
            .I(N__75710));
    Span4Mux_h I__16930 (
            .O(N__75723),
            .I(N__75710));
    Span4Mux_h I__16929 (
            .O(N__75720),
            .I(N__75707));
    Odrv4 I__16928 (
            .O(N__75717),
            .I(\pid_front.N_64 ));
    Odrv4 I__16927 (
            .O(N__75710),
            .I(\pid_front.N_64 ));
    Odrv4 I__16926 (
            .O(N__75707),
            .I(\pid_front.N_64 ));
    InMux I__16925 (
            .O(N__75700),
            .I(N__75697));
    LocalMux I__16924 (
            .O(N__75697),
            .I(N__75692));
    InMux I__16923 (
            .O(N__75696),
            .I(N__75687));
    InMux I__16922 (
            .O(N__75695),
            .I(N__75687));
    Span4Mux_h I__16921 (
            .O(N__75692),
            .I(N__75684));
    LocalMux I__16920 (
            .O(N__75687),
            .I(N__75681));
    Odrv4 I__16919 (
            .O(N__75684),
            .I(\pid_front.error_i_reg_esr_RNIV4AUZ0Z_12 ));
    Odrv12 I__16918 (
            .O(N__75681),
            .I(\pid_front.error_i_reg_esr_RNIV4AUZ0Z_12 ));
    CascadeMux I__16917 (
            .O(N__75676),
            .I(N__75672));
    InMux I__16916 (
            .O(N__75675),
            .I(N__75666));
    InMux I__16915 (
            .O(N__75672),
            .I(N__75661));
    InMux I__16914 (
            .O(N__75671),
            .I(N__75661));
    InMux I__16913 (
            .O(N__75670),
            .I(N__75658));
    InMux I__16912 (
            .O(N__75669),
            .I(N__75655));
    LocalMux I__16911 (
            .O(N__75666),
            .I(N__75646));
    LocalMux I__16910 (
            .O(N__75661),
            .I(N__75646));
    LocalMux I__16909 (
            .O(N__75658),
            .I(N__75641));
    LocalMux I__16908 (
            .O(N__75655),
            .I(N__75641));
    InMux I__16907 (
            .O(N__75654),
            .I(N__75636));
    InMux I__16906 (
            .O(N__75653),
            .I(N__75636));
    InMux I__16905 (
            .O(N__75652),
            .I(N__75631));
    InMux I__16904 (
            .O(N__75651),
            .I(N__75631));
    Span4Mux_v I__16903 (
            .O(N__75646),
            .I(N__75628));
    Span4Mux_h I__16902 (
            .O(N__75641),
            .I(N__75625));
    LocalMux I__16901 (
            .O(N__75636),
            .I(\pid_front.un10lto12 ));
    LocalMux I__16900 (
            .O(N__75631),
            .I(\pid_front.un10lto12 ));
    Odrv4 I__16899 (
            .O(N__75628),
            .I(\pid_front.un10lto12 ));
    Odrv4 I__16898 (
            .O(N__75625),
            .I(\pid_front.un10lto12 ));
    InMux I__16897 (
            .O(N__75616),
            .I(N__75611));
    InMux I__16896 (
            .O(N__75615),
            .I(N__75608));
    InMux I__16895 (
            .O(N__75614),
            .I(N__75605));
    LocalMux I__16894 (
            .O(N__75611),
            .I(N__75602));
    LocalMux I__16893 (
            .O(N__75608),
            .I(N__75599));
    LocalMux I__16892 (
            .O(N__75605),
            .I(N__75596));
    Span12Mux_h I__16891 (
            .O(N__75602),
            .I(N__75593));
    Span4Mux_v I__16890 (
            .O(N__75599),
            .I(N__75590));
    Span4Mux_v I__16889 (
            .O(N__75596),
            .I(N__75587));
    Odrv12 I__16888 (
            .O(N__75593),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_0_c_RNI9AGE ));
    Odrv4 I__16887 (
            .O(N__75590),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_0_c_RNI9AGE ));
    Odrv4 I__16886 (
            .O(N__75587),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_0_c_RNI9AGE ));
    InMux I__16885 (
            .O(N__75580),
            .I(N__75577));
    LocalMux I__16884 (
            .O(N__75577),
            .I(N__75574));
    Span4Mux_h I__16883 (
            .O(N__75574),
            .I(N__75571));
    Odrv4 I__16882 (
            .O(N__75571),
            .I(\pid_front.error_i_acumm_preregZ0Z_1 ));
    InMux I__16881 (
            .O(N__75568),
            .I(N__75565));
    LocalMux I__16880 (
            .O(N__75565),
            .I(N__75561));
    CascadeMux I__16879 (
            .O(N__75564),
            .I(N__75558));
    Span4Mux_h I__16878 (
            .O(N__75561),
            .I(N__75554));
    InMux I__16877 (
            .O(N__75558),
            .I(N__75551));
    InMux I__16876 (
            .O(N__75557),
            .I(N__75548));
    Span4Mux_v I__16875 (
            .O(N__75554),
            .I(N__75543));
    LocalMux I__16874 (
            .O(N__75551),
            .I(N__75543));
    LocalMux I__16873 (
            .O(N__75548),
            .I(N__75540));
    Span4Mux_h I__16872 (
            .O(N__75543),
            .I(N__75537));
    Span4Mux_v I__16871 (
            .O(N__75540),
            .I(N__75532));
    Span4Mux_v I__16870 (
            .O(N__75537),
            .I(N__75532));
    Odrv4 I__16869 (
            .O(N__75532),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_1_c_RNICEHE ));
    CascadeMux I__16868 (
            .O(N__75529),
            .I(N__75526));
    InMux I__16867 (
            .O(N__75526),
            .I(N__75523));
    LocalMux I__16866 (
            .O(N__75523),
            .I(N__75520));
    Span4Mux_h I__16865 (
            .O(N__75520),
            .I(N__75517));
    Span4Mux_h I__16864 (
            .O(N__75517),
            .I(N__75514));
    Odrv4 I__16863 (
            .O(N__75514),
            .I(\pid_front.error_i_acumm_preregZ0Z_2 ));
    InMux I__16862 (
            .O(N__75511),
            .I(N__75506));
    InMux I__16861 (
            .O(N__75510),
            .I(N__75501));
    InMux I__16860 (
            .O(N__75509),
            .I(N__75501));
    LocalMux I__16859 (
            .O(N__75506),
            .I(N__75498));
    LocalMux I__16858 (
            .O(N__75501),
            .I(N__75495));
    Span4Mux_v I__16857 (
            .O(N__75498),
            .I(N__75492));
    Span4Mux_h I__16856 (
            .O(N__75495),
            .I(N__75489));
    Odrv4 I__16855 (
            .O(N__75492),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_3_c_RNI9CPM ));
    Odrv4 I__16854 (
            .O(N__75489),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_3_c_RNI9CPM ));
    InMux I__16853 (
            .O(N__75484),
            .I(N__75480));
    InMux I__16852 (
            .O(N__75483),
            .I(N__75477));
    LocalMux I__16851 (
            .O(N__75480),
            .I(N__75472));
    LocalMux I__16850 (
            .O(N__75477),
            .I(N__75472));
    Span4Mux_v I__16849 (
            .O(N__75472),
            .I(N__75467));
    InMux I__16848 (
            .O(N__75471),
            .I(N__75462));
    InMux I__16847 (
            .O(N__75470),
            .I(N__75462));
    Span4Mux_h I__16846 (
            .O(N__75467),
            .I(N__75459));
    LocalMux I__16845 (
            .O(N__75462),
            .I(N__75456));
    Odrv4 I__16844 (
            .O(N__75459),
            .I(\pid_front.error_i_acumm_preregZ0Z_4 ));
    Odrv4 I__16843 (
            .O(N__75456),
            .I(\pid_front.error_i_acumm_preregZ0Z_4 ));
    InMux I__16842 (
            .O(N__75451),
            .I(N__75446));
    InMux I__16841 (
            .O(N__75450),
            .I(N__75443));
    InMux I__16840 (
            .O(N__75449),
            .I(N__75440));
    LocalMux I__16839 (
            .O(N__75446),
            .I(N__75437));
    LocalMux I__16838 (
            .O(N__75443),
            .I(N__75434));
    LocalMux I__16837 (
            .O(N__75440),
            .I(N__75431));
    Span4Mux_v I__16836 (
            .O(N__75437),
            .I(N__75428));
    Span4Mux_v I__16835 (
            .O(N__75434),
            .I(N__75425));
    Span4Mux_v I__16834 (
            .O(N__75431),
            .I(N__75420));
    Span4Mux_v I__16833 (
            .O(N__75428),
            .I(N__75420));
    Span4Mux_h I__16832 (
            .O(N__75425),
            .I(N__75417));
    Odrv4 I__16831 (
            .O(N__75420),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_6_c_RNIIOSM ));
    Odrv4 I__16830 (
            .O(N__75417),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_6_c_RNIIOSM ));
    CascadeMux I__16829 (
            .O(N__75412),
            .I(N__75409));
    InMux I__16828 (
            .O(N__75409),
            .I(N__75404));
    InMux I__16827 (
            .O(N__75408),
            .I(N__75399));
    InMux I__16826 (
            .O(N__75407),
            .I(N__75399));
    LocalMux I__16825 (
            .O(N__75404),
            .I(N__75396));
    LocalMux I__16824 (
            .O(N__75399),
            .I(N__75393));
    Span4Mux_v I__16823 (
            .O(N__75396),
            .I(N__75390));
    Span4Mux_h I__16822 (
            .O(N__75393),
            .I(N__75387));
    Odrv4 I__16821 (
            .O(N__75390),
            .I(\pid_front.error_i_acumm_preregZ0Z_7 ));
    Odrv4 I__16820 (
            .O(N__75387),
            .I(\pid_front.error_i_acumm_preregZ0Z_7 ));
    InMux I__16819 (
            .O(N__75382),
            .I(N__75377));
    InMux I__16818 (
            .O(N__75381),
            .I(N__75372));
    InMux I__16817 (
            .O(N__75380),
            .I(N__75372));
    LocalMux I__16816 (
            .O(N__75377),
            .I(N__75369));
    LocalMux I__16815 (
            .O(N__75372),
            .I(N__75366));
    Span4Mux_v I__16814 (
            .O(N__75369),
            .I(N__75363));
    Span4Mux_v I__16813 (
            .O(N__75366),
            .I(N__75360));
    Odrv4 I__16812 (
            .O(N__75363),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_7_c_RNIU6OE ));
    Odrv4 I__16811 (
            .O(N__75360),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_7_c_RNIU6OE ));
    InMux I__16810 (
            .O(N__75355),
            .I(N__75350));
    InMux I__16809 (
            .O(N__75354),
            .I(N__75345));
    InMux I__16808 (
            .O(N__75353),
            .I(N__75345));
    LocalMux I__16807 (
            .O(N__75350),
            .I(N__75342));
    LocalMux I__16806 (
            .O(N__75345),
            .I(N__75339));
    Span4Mux_v I__16805 (
            .O(N__75342),
            .I(N__75336));
    Span4Mux_h I__16804 (
            .O(N__75339),
            .I(N__75333));
    Odrv4 I__16803 (
            .O(N__75336),
            .I(\pid_front.error_i_acumm_preregZ0Z_8 ));
    Odrv4 I__16802 (
            .O(N__75333),
            .I(\pid_front.error_i_acumm_preregZ0Z_8 ));
    CEMux I__16801 (
            .O(N__75328),
            .I(N__75289));
    CEMux I__16800 (
            .O(N__75327),
            .I(N__75289));
    CEMux I__16799 (
            .O(N__75326),
            .I(N__75289));
    CEMux I__16798 (
            .O(N__75325),
            .I(N__75289));
    CEMux I__16797 (
            .O(N__75324),
            .I(N__75289));
    CEMux I__16796 (
            .O(N__75323),
            .I(N__75289));
    CEMux I__16795 (
            .O(N__75322),
            .I(N__75289));
    CEMux I__16794 (
            .O(N__75321),
            .I(N__75289));
    CEMux I__16793 (
            .O(N__75320),
            .I(N__75289));
    CEMux I__16792 (
            .O(N__75319),
            .I(N__75289));
    CEMux I__16791 (
            .O(N__75318),
            .I(N__75289));
    CEMux I__16790 (
            .O(N__75317),
            .I(N__75289));
    CEMux I__16789 (
            .O(N__75316),
            .I(N__75289));
    GlobalMux I__16788 (
            .O(N__75289),
            .I(N__75286));
    gio2CtrlBuf I__16787 (
            .O(N__75286),
            .I(\pid_front.state_0_g_0 ));
    InMux I__16786 (
            .O(N__75283),
            .I(N__75277));
    InMux I__16785 (
            .O(N__75282),
            .I(N__75274));
    InMux I__16784 (
            .O(N__75281),
            .I(N__75269));
    InMux I__16783 (
            .O(N__75280),
            .I(N__75269));
    LocalMux I__16782 (
            .O(N__75277),
            .I(N__75266));
    LocalMux I__16781 (
            .O(N__75274),
            .I(N__75261));
    LocalMux I__16780 (
            .O(N__75269),
            .I(N__75261));
    Span4Mux_h I__16779 (
            .O(N__75266),
            .I(N__75258));
    Span4Mux_v I__16778 (
            .O(N__75261),
            .I(N__75255));
    Odrv4 I__16777 (
            .O(N__75258),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_4_c_RNICGQM ));
    Odrv4 I__16776 (
            .O(N__75255),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_4_c_RNICGQM ));
    InMux I__16775 (
            .O(N__75250),
            .I(N__75247));
    LocalMux I__16774 (
            .O(N__75247),
            .I(N__75244));
    Span4Mux_h I__16773 (
            .O(N__75244),
            .I(N__75239));
    InMux I__16772 (
            .O(N__75243),
            .I(N__75236));
    InMux I__16771 (
            .O(N__75242),
            .I(N__75233));
    Odrv4 I__16770 (
            .O(N__75239),
            .I(\pid_front.error_i_acumm_preregZ0Z_5 ));
    LocalMux I__16769 (
            .O(N__75236),
            .I(\pid_front.error_i_acumm_preregZ0Z_5 ));
    LocalMux I__16768 (
            .O(N__75233),
            .I(\pid_front.error_i_acumm_preregZ0Z_5 ));
    InMux I__16767 (
            .O(N__75226),
            .I(N__75219));
    InMux I__16766 (
            .O(N__75225),
            .I(N__75219));
    InMux I__16765 (
            .O(N__75224),
            .I(N__75216));
    LocalMux I__16764 (
            .O(N__75219),
            .I(N__75213));
    LocalMux I__16763 (
            .O(N__75216),
            .I(N__75210));
    Span4Mux_h I__16762 (
            .O(N__75213),
            .I(N__75207));
    Span4Mux_h I__16761 (
            .O(N__75210),
            .I(N__75204));
    Span4Mux_v I__16760 (
            .O(N__75207),
            .I(N__75201));
    Odrv4 I__16759 (
            .O(N__75204),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_5_c_RNIOULE ));
    Odrv4 I__16758 (
            .O(N__75201),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_5_c_RNIOULE ));
    InMux I__16757 (
            .O(N__75196),
            .I(N__75193));
    LocalMux I__16756 (
            .O(N__75193),
            .I(N__75189));
    CascadeMux I__16755 (
            .O(N__75192),
            .I(N__75185));
    Span4Mux_v I__16754 (
            .O(N__75189),
            .I(N__75182));
    InMux I__16753 (
            .O(N__75188),
            .I(N__75177));
    InMux I__16752 (
            .O(N__75185),
            .I(N__75177));
    Odrv4 I__16751 (
            .O(N__75182),
            .I(\pid_front.error_i_acumm_preregZ0Z_6 ));
    LocalMux I__16750 (
            .O(N__75177),
            .I(\pid_front.error_i_acumm_preregZ0Z_6 ));
    InMux I__16749 (
            .O(N__75172),
            .I(N__75167));
    InMux I__16748 (
            .O(N__75171),
            .I(N__75162));
    InMux I__16747 (
            .O(N__75170),
            .I(N__75162));
    LocalMux I__16746 (
            .O(N__75167),
            .I(N__75157));
    LocalMux I__16745 (
            .O(N__75162),
            .I(N__75157));
    Span4Mux_v I__16744 (
            .O(N__75157),
            .I(N__75154));
    Odrv4 I__16743 (
            .O(N__75154),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_9_c_RNIIPQK ));
    CascadeMux I__16742 (
            .O(N__75151),
            .I(N__75148));
    InMux I__16741 (
            .O(N__75148),
            .I(N__75145));
    LocalMux I__16740 (
            .O(N__75145),
            .I(N__75141));
    InMux I__16739 (
            .O(N__75144),
            .I(N__75138));
    Span4Mux_v I__16738 (
            .O(N__75141),
            .I(N__75131));
    LocalMux I__16737 (
            .O(N__75138),
            .I(N__75131));
    InMux I__16736 (
            .O(N__75137),
            .I(N__75126));
    InMux I__16735 (
            .O(N__75136),
            .I(N__75126));
    Span4Mux_h I__16734 (
            .O(N__75131),
            .I(N__75123));
    LocalMux I__16733 (
            .O(N__75126),
            .I(N__75120));
    Odrv4 I__16732 (
            .O(N__75123),
            .I(\pid_front.error_i_reg_esr_RNIS09UZ0Z_11 ));
    Odrv4 I__16731 (
            .O(N__75120),
            .I(\pid_front.error_i_reg_esr_RNIS09UZ0Z_11 ));
    InMux I__16730 (
            .O(N__75115),
            .I(N__75112));
    LocalMux I__16729 (
            .O(N__75112),
            .I(N__75105));
    InMux I__16728 (
            .O(N__75111),
            .I(N__75102));
    InMux I__16727 (
            .O(N__75110),
            .I(N__75095));
    InMux I__16726 (
            .O(N__75109),
            .I(N__75095));
    InMux I__16725 (
            .O(N__75108),
            .I(N__75092));
    Span4Mux_v I__16724 (
            .O(N__75105),
            .I(N__75087));
    LocalMux I__16723 (
            .O(N__75102),
            .I(N__75087));
    InMux I__16722 (
            .O(N__75101),
            .I(N__75082));
    InMux I__16721 (
            .O(N__75100),
            .I(N__75082));
    LocalMux I__16720 (
            .O(N__75095),
            .I(\pid_front.error_i_acumm_preregZ0Z_10 ));
    LocalMux I__16719 (
            .O(N__75092),
            .I(\pid_front.error_i_acumm_preregZ0Z_10 ));
    Odrv4 I__16718 (
            .O(N__75087),
            .I(\pid_front.error_i_acumm_preregZ0Z_10 ));
    LocalMux I__16717 (
            .O(N__75082),
            .I(\pid_front.error_i_acumm_preregZ0Z_10 ));
    CascadeMux I__16716 (
            .O(N__75073),
            .I(\pid_front.N_355_cascade_ ));
    InMux I__16715 (
            .O(N__75070),
            .I(N__75067));
    LocalMux I__16714 (
            .O(N__75067),
            .I(N__75064));
    Span4Mux_h I__16713 (
            .O(N__75064),
            .I(N__75061));
    Odrv4 I__16712 (
            .O(N__75061),
            .I(\pid_front.error_i_acummZ0Z_10 ));
    InMux I__16711 (
            .O(N__75058),
            .I(N__75052));
    InMux I__16710 (
            .O(N__75057),
            .I(N__75047));
    InMux I__16709 (
            .O(N__75056),
            .I(N__75047));
    InMux I__16708 (
            .O(N__75055),
            .I(N__75044));
    LocalMux I__16707 (
            .O(N__75052),
            .I(N__75041));
    LocalMux I__16706 (
            .O(N__75047),
            .I(N__75036));
    LocalMux I__16705 (
            .O(N__75044),
            .I(N__75036));
    Odrv4 I__16704 (
            .O(N__75041),
            .I(\pid_front.N_203 ));
    Odrv4 I__16703 (
            .O(N__75036),
            .I(\pid_front.N_203 ));
    InMux I__16702 (
            .O(N__75031),
            .I(N__75028));
    LocalMux I__16701 (
            .O(N__75028),
            .I(N__75021));
    InMux I__16700 (
            .O(N__75027),
            .I(N__75017));
    CascadeMux I__16699 (
            .O(N__75026),
            .I(N__75014));
    InMux I__16698 (
            .O(N__75025),
            .I(N__75008));
    InMux I__16697 (
            .O(N__75024),
            .I(N__75008));
    Span4Mux_h I__16696 (
            .O(N__75021),
            .I(N__75005));
    InMux I__16695 (
            .O(N__75020),
            .I(N__75002));
    LocalMux I__16694 (
            .O(N__75017),
            .I(N__74999));
    InMux I__16693 (
            .O(N__75014),
            .I(N__74994));
    InMux I__16692 (
            .O(N__75013),
            .I(N__74994));
    LocalMux I__16691 (
            .O(N__75008),
            .I(\pid_front.error_i_acumm_preregZ0Z_11 ));
    Odrv4 I__16690 (
            .O(N__75005),
            .I(\pid_front.error_i_acumm_preregZ0Z_11 ));
    LocalMux I__16689 (
            .O(N__75002),
            .I(\pid_front.error_i_acumm_preregZ0Z_11 ));
    Odrv4 I__16688 (
            .O(N__74999),
            .I(\pid_front.error_i_acumm_preregZ0Z_11 ));
    LocalMux I__16687 (
            .O(N__74994),
            .I(\pid_front.error_i_acumm_preregZ0Z_11 ));
    CascadeMux I__16686 (
            .O(N__74983),
            .I(\pid_front.N_353_cascade_ ));
    InMux I__16685 (
            .O(N__74980),
            .I(N__74977));
    LocalMux I__16684 (
            .O(N__74977),
            .I(N__74974));
    Span4Mux_h I__16683 (
            .O(N__74974),
            .I(N__74971));
    Odrv4 I__16682 (
            .O(N__74971),
            .I(\pid_front.error_i_acummZ0Z_11 ));
    InMux I__16681 (
            .O(N__74968),
            .I(N__74959));
    CascadeMux I__16680 (
            .O(N__74967),
            .I(N__74955));
    InMux I__16679 (
            .O(N__74966),
            .I(N__74952));
    InMux I__16678 (
            .O(N__74965),
            .I(N__74949));
    InMux I__16677 (
            .O(N__74964),
            .I(N__74946));
    InMux I__16676 (
            .O(N__74963),
            .I(N__74943));
    InMux I__16675 (
            .O(N__74962),
            .I(N__74939));
    LocalMux I__16674 (
            .O(N__74959),
            .I(N__74936));
    InMux I__16673 (
            .O(N__74958),
            .I(N__74932));
    InMux I__16672 (
            .O(N__74955),
            .I(N__74929));
    LocalMux I__16671 (
            .O(N__74952),
            .I(N__74920));
    LocalMux I__16670 (
            .O(N__74949),
            .I(N__74920));
    LocalMux I__16669 (
            .O(N__74946),
            .I(N__74920));
    LocalMux I__16668 (
            .O(N__74943),
            .I(N__74920));
    InMux I__16667 (
            .O(N__74942),
            .I(N__74917));
    LocalMux I__16666 (
            .O(N__74939),
            .I(N__74914));
    Span4Mux_h I__16665 (
            .O(N__74936),
            .I(N__74911));
    InMux I__16664 (
            .O(N__74935),
            .I(N__74908));
    LocalMux I__16663 (
            .O(N__74932),
            .I(N__74905));
    LocalMux I__16662 (
            .O(N__74929),
            .I(N__74902));
    Span4Mux_v I__16661 (
            .O(N__74920),
            .I(N__74897));
    LocalMux I__16660 (
            .O(N__74917),
            .I(N__74897));
    Span4Mux_h I__16659 (
            .O(N__74914),
            .I(N__74890));
    Span4Mux_v I__16658 (
            .O(N__74911),
            .I(N__74890));
    LocalMux I__16657 (
            .O(N__74908),
            .I(N__74890));
    Span4Mux_v I__16656 (
            .O(N__74905),
            .I(N__74885));
    Span4Mux_v I__16655 (
            .O(N__74902),
            .I(N__74885));
    Span4Mux_h I__16654 (
            .O(N__74897),
            .I(N__74882));
    Odrv4 I__16653 (
            .O(N__74890),
            .I(pid_side_N_495));
    Odrv4 I__16652 (
            .O(N__74885),
            .I(pid_side_N_495));
    Odrv4 I__16651 (
            .O(N__74882),
            .I(pid_side_N_495));
    CascadeMux I__16650 (
            .O(N__74875),
            .I(\pid_front.N_569_cascade_ ));
    CascadeMux I__16649 (
            .O(N__74872),
            .I(N__74868));
    InMux I__16648 (
            .O(N__74871),
            .I(N__74865));
    InMux I__16647 (
            .O(N__74868),
            .I(N__74862));
    LocalMux I__16646 (
            .O(N__74865),
            .I(N__74859));
    LocalMux I__16645 (
            .O(N__74862),
            .I(N__74853));
    Span4Mux_s1_h I__16644 (
            .O(N__74859),
            .I(N__74850));
    InMux I__16643 (
            .O(N__74858),
            .I(N__74846));
    InMux I__16642 (
            .O(N__74857),
            .I(N__74843));
    InMux I__16641 (
            .O(N__74856),
            .I(N__74840));
    Span4Mux_h I__16640 (
            .O(N__74853),
            .I(N__74836));
    Span4Mux_h I__16639 (
            .O(N__74850),
            .I(N__74833));
    InMux I__16638 (
            .O(N__74849),
            .I(N__74830));
    LocalMux I__16637 (
            .O(N__74846),
            .I(N__74827));
    LocalMux I__16636 (
            .O(N__74843),
            .I(N__74824));
    LocalMux I__16635 (
            .O(N__74840),
            .I(N__74821));
    InMux I__16634 (
            .O(N__74839),
            .I(N__74818));
    Span4Mux_v I__16633 (
            .O(N__74836),
            .I(N__74815));
    Span4Mux_h I__16632 (
            .O(N__74833),
            .I(N__74811));
    LocalMux I__16631 (
            .O(N__74830),
            .I(N__74806));
    Span4Mux_h I__16630 (
            .O(N__74827),
            .I(N__74806));
    Span4Mux_h I__16629 (
            .O(N__74824),
            .I(N__74803));
    Span4Mux_v I__16628 (
            .O(N__74821),
            .I(N__74800));
    LocalMux I__16627 (
            .O(N__74818),
            .I(N__74795));
    Span4Mux_v I__16626 (
            .O(N__74815),
            .I(N__74795));
    InMux I__16625 (
            .O(N__74814),
            .I(N__74792));
    Span4Mux_h I__16624 (
            .O(N__74811),
            .I(N__74788));
    Span4Mux_h I__16623 (
            .O(N__74806),
            .I(N__74783));
    Span4Mux_h I__16622 (
            .O(N__74803),
            .I(N__74783));
    Sp12to4 I__16621 (
            .O(N__74800),
            .I(N__74776));
    Sp12to4 I__16620 (
            .O(N__74795),
            .I(N__74776));
    LocalMux I__16619 (
            .O(N__74792),
            .I(N__74776));
    InMux I__16618 (
            .O(N__74791),
            .I(N__74773));
    Span4Mux_v I__16617 (
            .O(N__74788),
            .I(N__74768));
    Span4Mux_h I__16616 (
            .O(N__74783),
            .I(N__74768));
    Odrv12 I__16615 (
            .O(N__74776),
            .I(\pid_front.error_8 ));
    LocalMux I__16614 (
            .O(N__74773),
            .I(\pid_front.error_8 ));
    Odrv4 I__16613 (
            .O(N__74768),
            .I(\pid_front.error_8 ));
    InMux I__16612 (
            .O(N__74761),
            .I(N__74758));
    LocalMux I__16611 (
            .O(N__74758),
            .I(\pid_front.error_i_reg_9_sn_13 ));
    InMux I__16610 (
            .O(N__74755),
            .I(N__74752));
    LocalMux I__16609 (
            .O(N__74752),
            .I(N__74749));
    Span4Mux_v I__16608 (
            .O(N__74749),
            .I(N__74746));
    Span4Mux_v I__16607 (
            .O(N__74746),
            .I(N__74743));
    Odrv4 I__16606 (
            .O(N__74743),
            .I(\pid_front.error_i_reg_9_rn_2_13 ));
    CascadeMux I__16605 (
            .O(N__74740),
            .I(\pid_front.N_436_cascade_ ));
    CascadeMux I__16604 (
            .O(N__74737),
            .I(N__74734));
    InMux I__16603 (
            .O(N__74734),
            .I(N__74731));
    LocalMux I__16602 (
            .O(N__74731),
            .I(N__74728));
    Span4Mux_h I__16601 (
            .O(N__74728),
            .I(N__74725));
    Odrv4 I__16600 (
            .O(N__74725),
            .I(\pid_front.error_i_regZ0Z_13 ));
    InMux I__16599 (
            .O(N__74722),
            .I(N__74718));
    InMux I__16598 (
            .O(N__74721),
            .I(N__74713));
    LocalMux I__16597 (
            .O(N__74718),
            .I(N__74710));
    InMux I__16596 (
            .O(N__74717),
            .I(N__74707));
    InMux I__16595 (
            .O(N__74716),
            .I(N__74704));
    LocalMux I__16594 (
            .O(N__74713),
            .I(N__74699));
    Span4Mux_v I__16593 (
            .O(N__74710),
            .I(N__74699));
    LocalMux I__16592 (
            .O(N__74707),
            .I(\pid_front.N_184 ));
    LocalMux I__16591 (
            .O(N__74704),
            .I(\pid_front.N_184 ));
    Odrv4 I__16590 (
            .O(N__74699),
            .I(\pid_front.N_184 ));
    CascadeMux I__16589 (
            .O(N__74692),
            .I(N__74687));
    InMux I__16588 (
            .O(N__74691),
            .I(N__74684));
    InMux I__16587 (
            .O(N__74690),
            .I(N__74681));
    InMux I__16586 (
            .O(N__74687),
            .I(N__74678));
    LocalMux I__16585 (
            .O(N__74684),
            .I(N__74674));
    LocalMux I__16584 (
            .O(N__74681),
            .I(N__74671));
    LocalMux I__16583 (
            .O(N__74678),
            .I(N__74668));
    InMux I__16582 (
            .O(N__74677),
            .I(N__74665));
    Span4Mux_v I__16581 (
            .O(N__74674),
            .I(N__74662));
    Span4Mux_h I__16580 (
            .O(N__74671),
            .I(N__74655));
    Span4Mux_v I__16579 (
            .O(N__74668),
            .I(N__74655));
    LocalMux I__16578 (
            .O(N__74665),
            .I(N__74655));
    Span4Mux_h I__16577 (
            .O(N__74662),
            .I(N__74652));
    Span4Mux_h I__16576 (
            .O(N__74655),
            .I(N__74649));
    Odrv4 I__16575 (
            .O(N__74652),
            .I(\pid_front.N_231 ));
    Odrv4 I__16574 (
            .O(N__74649),
            .I(\pid_front.N_231 ));
    InMux I__16573 (
            .O(N__74644),
            .I(N__74641));
    LocalMux I__16572 (
            .O(N__74641),
            .I(\pid_front.N_437 ));
    InMux I__16571 (
            .O(N__74638),
            .I(N__74635));
    LocalMux I__16570 (
            .O(N__74635),
            .I(N__74632));
    Span4Mux_h I__16569 (
            .O(N__74632),
            .I(N__74629));
    Span4Mux_h I__16568 (
            .O(N__74629),
            .I(N__74626));
    Odrv4 I__16567 (
            .O(N__74626),
            .I(\pid_front.m10_2_03_3_i_0_a2_0 ));
    InMux I__16566 (
            .O(N__74623),
            .I(N__74620));
    LocalMux I__16565 (
            .O(N__74620),
            .I(\pid_front.error_i_acumm_13_0_a2_2_2_2 ));
    InMux I__16564 (
            .O(N__74617),
            .I(N__74614));
    LocalMux I__16563 (
            .O(N__74614),
            .I(N__74611));
    Odrv12 I__16562 (
            .O(N__74611),
            .I(\pid_front.N_603 ));
    CascadeMux I__16561 (
            .O(N__74608),
            .I(\pid_front.N_603_cascade_ ));
    InMux I__16560 (
            .O(N__74605),
            .I(N__74602));
    LocalMux I__16559 (
            .O(N__74602),
            .I(N__74599));
    Span4Mux_v I__16558 (
            .O(N__74599),
            .I(N__74596));
    Odrv4 I__16557 (
            .O(N__74596),
            .I(\pid_front.error_i_acumm_13_0_a2_3_1_2 ));
    InMux I__16556 (
            .O(N__74593),
            .I(N__74590));
    LocalMux I__16555 (
            .O(N__74590),
            .I(N__74585));
    InMux I__16554 (
            .O(N__74589),
            .I(N__74580));
    InMux I__16553 (
            .O(N__74588),
            .I(N__74580));
    Span4Mux_v I__16552 (
            .O(N__74585),
            .I(N__74577));
    LocalMux I__16551 (
            .O(N__74580),
            .I(N__74574));
    Odrv4 I__16550 (
            .O(N__74577),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_2_c_RNI68OM ));
    Odrv4 I__16549 (
            .O(N__74574),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_2_c_RNI68OM ));
    InMux I__16548 (
            .O(N__74569),
            .I(N__74565));
    CascadeMux I__16547 (
            .O(N__74568),
            .I(N__74561));
    LocalMux I__16546 (
            .O(N__74565),
            .I(N__74558));
    InMux I__16545 (
            .O(N__74564),
            .I(N__74555));
    InMux I__16544 (
            .O(N__74561),
            .I(N__74552));
    Odrv12 I__16543 (
            .O(N__74558),
            .I(\pid_front.error_i_acumm16lto3 ));
    LocalMux I__16542 (
            .O(N__74555),
            .I(\pid_front.error_i_acumm16lto3 ));
    LocalMux I__16541 (
            .O(N__74552),
            .I(\pid_front.error_i_acumm16lto3 ));
    CascadeMux I__16540 (
            .O(N__74545),
            .I(\pid_front.N_226_cascade_ ));
    InMux I__16539 (
            .O(N__74542),
            .I(N__74539));
    LocalMux I__16538 (
            .O(N__74539),
            .I(N__74536));
    Span4Mux_h I__16537 (
            .O(N__74536),
            .I(N__74533));
    Odrv4 I__16536 (
            .O(N__74533),
            .I(\pid_front.m21_2_03_0_0 ));
    InMux I__16535 (
            .O(N__74530),
            .I(N__74527));
    LocalMux I__16534 (
            .O(N__74527),
            .I(N__74524));
    Span4Mux_h I__16533 (
            .O(N__74524),
            .I(N__74521));
    Odrv4 I__16532 (
            .O(N__74521),
            .I(\pid_front.m22_2_03_0_0 ));
    InMux I__16531 (
            .O(N__74518),
            .I(N__74515));
    LocalMux I__16530 (
            .O(N__74515),
            .I(N__74511));
    InMux I__16529 (
            .O(N__74514),
            .I(N__74508));
    Span4Mux_v I__16528 (
            .O(N__74511),
            .I(N__74500));
    LocalMux I__16527 (
            .O(N__74508),
            .I(N__74497));
    InMux I__16526 (
            .O(N__74507),
            .I(N__74491));
    InMux I__16525 (
            .O(N__74506),
            .I(N__74488));
    InMux I__16524 (
            .O(N__74505),
            .I(N__74485));
    InMux I__16523 (
            .O(N__74504),
            .I(N__74480));
    InMux I__16522 (
            .O(N__74503),
            .I(N__74480));
    Span4Mux_h I__16521 (
            .O(N__74500),
            .I(N__74477));
    Span4Mux_v I__16520 (
            .O(N__74497),
            .I(N__74474));
    InMux I__16519 (
            .O(N__74496),
            .I(N__74470));
    InMux I__16518 (
            .O(N__74495),
            .I(N__74465));
    InMux I__16517 (
            .O(N__74494),
            .I(N__74465));
    LocalMux I__16516 (
            .O(N__74491),
            .I(N__74460));
    LocalMux I__16515 (
            .O(N__74488),
            .I(N__74460));
    LocalMux I__16514 (
            .O(N__74485),
            .I(N__74457));
    LocalMux I__16513 (
            .O(N__74480),
            .I(N__74454));
    Span4Mux_h I__16512 (
            .O(N__74477),
            .I(N__74451));
    Span4Mux_h I__16511 (
            .O(N__74474),
            .I(N__74448));
    InMux I__16510 (
            .O(N__74473),
            .I(N__74445));
    LocalMux I__16509 (
            .O(N__74470),
            .I(N__74442));
    LocalMux I__16508 (
            .O(N__74465),
            .I(N__74439));
    Span4Mux_v I__16507 (
            .O(N__74460),
            .I(N__74432));
    Span4Mux_v I__16506 (
            .O(N__74457),
            .I(N__74432));
    Span4Mux_v I__16505 (
            .O(N__74454),
            .I(N__74432));
    Span4Mux_h I__16504 (
            .O(N__74451),
            .I(N__74429));
    Span4Mux_h I__16503 (
            .O(N__74448),
            .I(N__74426));
    LocalMux I__16502 (
            .O(N__74445),
            .I(N__74421));
    Span4Mux_h I__16501 (
            .O(N__74442),
            .I(N__74421));
    Span4Mux_v I__16500 (
            .O(N__74439),
            .I(N__74418));
    Span4Mux_h I__16499 (
            .O(N__74432),
            .I(N__74415));
    Odrv4 I__16498 (
            .O(N__74429),
            .I(\pid_front.error_11 ));
    Odrv4 I__16497 (
            .O(N__74426),
            .I(\pid_front.error_11 ));
    Odrv4 I__16496 (
            .O(N__74421),
            .I(\pid_front.error_11 ));
    Odrv4 I__16495 (
            .O(N__74418),
            .I(\pid_front.error_11 ));
    Odrv4 I__16494 (
            .O(N__74415),
            .I(\pid_front.error_11 ));
    InMux I__16493 (
            .O(N__74404),
            .I(N__74401));
    LocalMux I__16492 (
            .O(N__74401),
            .I(\pid_front.N_254 ));
    CascadeMux I__16491 (
            .O(N__74398),
            .I(\pid_front.N_254_cascade_ ));
    CascadeMux I__16490 (
            .O(N__74395),
            .I(\pid_front.error_i_reg_9_N_2L1_1_cascade_ ));
    InMux I__16489 (
            .O(N__74392),
            .I(N__74383));
    InMux I__16488 (
            .O(N__74391),
            .I(N__74383));
    InMux I__16487 (
            .O(N__74390),
            .I(N__74383));
    LocalMux I__16486 (
            .O(N__74383),
            .I(\pid_front.N_226 ));
    InMux I__16485 (
            .O(N__74380),
            .I(N__74377));
    LocalMux I__16484 (
            .O(N__74377),
            .I(\pid_front.error_i_reg_esr_RNO_0Z0Z_16 ));
    InMux I__16483 (
            .O(N__74374),
            .I(N__74368));
    InMux I__16482 (
            .O(N__74373),
            .I(N__74363));
    InMux I__16481 (
            .O(N__74372),
            .I(N__74363));
    InMux I__16480 (
            .O(N__74371),
            .I(N__74360));
    LocalMux I__16479 (
            .O(N__74368),
            .I(N__74357));
    LocalMux I__16478 (
            .O(N__74363),
            .I(N__74353));
    LocalMux I__16477 (
            .O(N__74360),
            .I(N__74350));
    Span4Mux_h I__16476 (
            .O(N__74357),
            .I(N__74347));
    InMux I__16475 (
            .O(N__74356),
            .I(N__74344));
    Sp12to4 I__16474 (
            .O(N__74353),
            .I(N__74339));
    Span12Mux_v I__16473 (
            .O(N__74350),
            .I(N__74339));
    Odrv4 I__16472 (
            .O(N__74347),
            .I(\pid_front.N_594 ));
    LocalMux I__16471 (
            .O(N__74344),
            .I(\pid_front.N_594 ));
    Odrv12 I__16470 (
            .O(N__74339),
            .I(\pid_front.N_594 ));
    InMux I__16469 (
            .O(N__74332),
            .I(N__74329));
    LocalMux I__16468 (
            .O(N__74329),
            .I(N__74326));
    Span4Mux_h I__16467 (
            .O(N__74326),
            .I(N__74323));
    Odrv4 I__16466 (
            .O(N__74323),
            .I(\pid_front.N_611 ));
    InMux I__16465 (
            .O(N__74320),
            .I(N__74314));
    InMux I__16464 (
            .O(N__74319),
            .I(N__74308));
    InMux I__16463 (
            .O(N__74318),
            .I(N__74305));
    CascadeMux I__16462 (
            .O(N__74317),
            .I(N__74301));
    LocalMux I__16461 (
            .O(N__74314),
            .I(N__74297));
    InMux I__16460 (
            .O(N__74313),
            .I(N__74294));
    InMux I__16459 (
            .O(N__74312),
            .I(N__74289));
    InMux I__16458 (
            .O(N__74311),
            .I(N__74289));
    LocalMux I__16457 (
            .O(N__74308),
            .I(N__74284));
    LocalMux I__16456 (
            .O(N__74305),
            .I(N__74284));
    InMux I__16455 (
            .O(N__74304),
            .I(N__74277));
    InMux I__16454 (
            .O(N__74301),
            .I(N__74277));
    InMux I__16453 (
            .O(N__74300),
            .I(N__74277));
    Span4Mux_v I__16452 (
            .O(N__74297),
            .I(N__74274));
    LocalMux I__16451 (
            .O(N__74294),
            .I(N__74271));
    LocalMux I__16450 (
            .O(N__74289),
            .I(N__74267));
    Span4Mux_v I__16449 (
            .O(N__74284),
            .I(N__74261));
    LocalMux I__16448 (
            .O(N__74277),
            .I(N__74261));
    Span4Mux_v I__16447 (
            .O(N__74274),
            .I(N__74258));
    Span12Mux_v I__16446 (
            .O(N__74271),
            .I(N__74255));
    InMux I__16445 (
            .O(N__74270),
            .I(N__74252));
    Span4Mux_v I__16444 (
            .O(N__74267),
            .I(N__74249));
    InMux I__16443 (
            .O(N__74266),
            .I(N__74246));
    Span4Mux_h I__16442 (
            .O(N__74261),
            .I(N__74243));
    Sp12to4 I__16441 (
            .O(N__74258),
            .I(N__74232));
    Span12Mux_h I__16440 (
            .O(N__74255),
            .I(N__74232));
    LocalMux I__16439 (
            .O(N__74252),
            .I(N__74232));
    Sp12to4 I__16438 (
            .O(N__74249),
            .I(N__74232));
    LocalMux I__16437 (
            .O(N__74246),
            .I(N__74232));
    Span4Mux_v I__16436 (
            .O(N__74243),
            .I(N__74229));
    Odrv12 I__16435 (
            .O(N__74232),
            .I(\pid_front.error_12 ));
    Odrv4 I__16434 (
            .O(N__74229),
            .I(\pid_front.error_12 ));
    CascadeMux I__16433 (
            .O(N__74224),
            .I(\pid_front.error_cry_1_0_c_RNI590GZ0Z1_cascade_ ));
    InMux I__16432 (
            .O(N__74221),
            .I(N__74218));
    LocalMux I__16431 (
            .O(N__74218),
            .I(N__74215));
    Span4Mux_h I__16430 (
            .O(N__74215),
            .I(N__74211));
    InMux I__16429 (
            .O(N__74214),
            .I(N__74208));
    Sp12to4 I__16428 (
            .O(N__74211),
            .I(N__74202));
    LocalMux I__16427 (
            .O(N__74208),
            .I(N__74202));
    InMux I__16426 (
            .O(N__74207),
            .I(N__74199));
    Odrv12 I__16425 (
            .O(N__74202),
            .I(\pid_front.N_183 ));
    LocalMux I__16424 (
            .O(N__74199),
            .I(\pid_front.N_183 ));
    InMux I__16423 (
            .O(N__74194),
            .I(N__74191));
    LocalMux I__16422 (
            .O(N__74191),
            .I(\pid_front.error_cry_1_0_c_RNINTZ0Z963 ));
    InMux I__16421 (
            .O(N__74188),
            .I(N__74185));
    LocalMux I__16420 (
            .O(N__74185),
            .I(N__74180));
    InMux I__16419 (
            .O(N__74184),
            .I(N__74177));
    CascadeMux I__16418 (
            .O(N__74183),
            .I(N__74172));
    Span4Mux_v I__16417 (
            .O(N__74180),
            .I(N__74168));
    LocalMux I__16416 (
            .O(N__74177),
            .I(N__74165));
    InMux I__16415 (
            .O(N__74176),
            .I(N__74161));
    InMux I__16414 (
            .O(N__74175),
            .I(N__74158));
    InMux I__16413 (
            .O(N__74172),
            .I(N__74153));
    InMux I__16412 (
            .O(N__74171),
            .I(N__74153));
    Span4Mux_h I__16411 (
            .O(N__74168),
            .I(N__74150));
    Span4Mux_v I__16410 (
            .O(N__74165),
            .I(N__74147));
    InMux I__16409 (
            .O(N__74164),
            .I(N__74143));
    LocalMux I__16408 (
            .O(N__74161),
            .I(N__74138));
    LocalMux I__16407 (
            .O(N__74158),
            .I(N__74138));
    LocalMux I__16406 (
            .O(N__74153),
            .I(N__74135));
    Span4Mux_v I__16405 (
            .O(N__74150),
            .I(N__74129));
    Sp12to4 I__16404 (
            .O(N__74147),
            .I(N__74126));
    InMux I__16403 (
            .O(N__74146),
            .I(N__74123));
    LocalMux I__16402 (
            .O(N__74143),
            .I(N__74116));
    Span4Mux_v I__16401 (
            .O(N__74138),
            .I(N__74116));
    Span4Mux_v I__16400 (
            .O(N__74135),
            .I(N__74116));
    InMux I__16399 (
            .O(N__74134),
            .I(N__74113));
    InMux I__16398 (
            .O(N__74133),
            .I(N__74108));
    InMux I__16397 (
            .O(N__74132),
            .I(N__74108));
    Sp12to4 I__16396 (
            .O(N__74129),
            .I(N__74097));
    Span12Mux_s7_h I__16395 (
            .O(N__74126),
            .I(N__74097));
    LocalMux I__16394 (
            .O(N__74123),
            .I(N__74097));
    Sp12to4 I__16393 (
            .O(N__74116),
            .I(N__74097));
    LocalMux I__16392 (
            .O(N__74113),
            .I(N__74097));
    LocalMux I__16391 (
            .O(N__74108),
            .I(N__74094));
    Odrv12 I__16390 (
            .O(N__74097),
            .I(\pid_front.error_1 ));
    Odrv4 I__16389 (
            .O(N__74094),
            .I(\pid_front.error_1 ));
    CascadeMux I__16388 (
            .O(N__74089),
            .I(\pid_front.N_40_0_i_i_o2_0_cascade_ ));
    InMux I__16387 (
            .O(N__74086),
            .I(N__74083));
    LocalMux I__16386 (
            .O(N__74083),
            .I(N__74078));
    InMux I__16385 (
            .O(N__74082),
            .I(N__74073));
    InMux I__16384 (
            .O(N__74081),
            .I(N__74070));
    Span4Mux_v I__16383 (
            .O(N__74078),
            .I(N__74067));
    InMux I__16382 (
            .O(N__74077),
            .I(N__74063));
    InMux I__16381 (
            .O(N__74076),
            .I(N__74059));
    LocalMux I__16380 (
            .O(N__74073),
            .I(N__74056));
    LocalMux I__16379 (
            .O(N__74070),
            .I(N__74053));
    Span4Mux_h I__16378 (
            .O(N__74067),
            .I(N__74048));
    InMux I__16377 (
            .O(N__74066),
            .I(N__74045));
    LocalMux I__16376 (
            .O(N__74063),
            .I(N__74042));
    InMux I__16375 (
            .O(N__74062),
            .I(N__74039));
    LocalMux I__16374 (
            .O(N__74059),
            .I(N__74034));
    Span4Mux_h I__16373 (
            .O(N__74056),
            .I(N__74034));
    Span4Mux_v I__16372 (
            .O(N__74053),
            .I(N__74031));
    InMux I__16371 (
            .O(N__74052),
            .I(N__74026));
    InMux I__16370 (
            .O(N__74051),
            .I(N__74026));
    Span4Mux_h I__16369 (
            .O(N__74048),
            .I(N__74023));
    LocalMux I__16368 (
            .O(N__74045),
            .I(N__74020));
    Span4Mux_h I__16367 (
            .O(N__74042),
            .I(N__74017));
    LocalMux I__16366 (
            .O(N__74039),
            .I(N__74012));
    Span4Mux_h I__16365 (
            .O(N__74034),
            .I(N__74012));
    Span4Mux_h I__16364 (
            .O(N__74031),
            .I(N__74005));
    LocalMux I__16363 (
            .O(N__74026),
            .I(N__74005));
    Span4Mux_h I__16362 (
            .O(N__74023),
            .I(N__74005));
    Span12Mux_h I__16361 (
            .O(N__74020),
            .I(N__74002));
    Odrv4 I__16360 (
            .O(N__74017),
            .I(\pid_front.error_3 ));
    Odrv4 I__16359 (
            .O(N__74012),
            .I(\pid_front.error_3 ));
    Odrv4 I__16358 (
            .O(N__74005),
            .I(\pid_front.error_3 ));
    Odrv12 I__16357 (
            .O(N__74002),
            .I(\pid_front.error_3 ));
    CascadeMux I__16356 (
            .O(N__73993),
            .I(\pid_front.error_cry_2_c_RNIKGVOZ0Z2_cascade_ ));
    InMux I__16355 (
            .O(N__73990),
            .I(N__73987));
    LocalMux I__16354 (
            .O(N__73987),
            .I(N__73984));
    Span4Mux_v I__16353 (
            .O(N__73984),
            .I(N__73980));
    InMux I__16352 (
            .O(N__73983),
            .I(N__73977));
    Odrv4 I__16351 (
            .O(N__73980),
            .I(\pid_front.N_245 ));
    LocalMux I__16350 (
            .O(N__73977),
            .I(\pid_front.N_245 ));
    CascadeMux I__16349 (
            .O(N__73972),
            .I(\pid_front.error_i_reg_9_sn_rn_0_15_cascade_ ));
    InMux I__16348 (
            .O(N__73969),
            .I(N__73966));
    LocalMux I__16347 (
            .O(N__73966),
            .I(N__73963));
    Odrv12 I__16346 (
            .O(N__73963),
            .I(\pid_front.m19_2_03_0_0 ));
    InMux I__16345 (
            .O(N__73960),
            .I(N__73957));
    LocalMux I__16344 (
            .O(N__73957),
            .I(N__73954));
    Odrv4 I__16343 (
            .O(N__73954),
            .I(\pid_front.error_i_reg_9_rn_1_15 ));
    CascadeMux I__16342 (
            .O(N__73951),
            .I(\pid_front.error_i_reg_9_sn_15_cascade_ ));
    InMux I__16341 (
            .O(N__73948),
            .I(N__73945));
    LocalMux I__16340 (
            .O(N__73945),
            .I(\pid_front.m19_2_03_0_1 ));
    CascadeMux I__16339 (
            .O(N__73942),
            .I(N__73939));
    InMux I__16338 (
            .O(N__73939),
            .I(N__73936));
    LocalMux I__16337 (
            .O(N__73936),
            .I(N__73933));
    Span4Mux_h I__16336 (
            .O(N__73933),
            .I(N__73930));
    Odrv4 I__16335 (
            .O(N__73930),
            .I(\pid_front.error_i_regZ0Z_15 ));
    CascadeMux I__16334 (
            .O(N__73927),
            .I(\pid_side.N_185_cascade_ ));
    InMux I__16333 (
            .O(N__73924),
            .I(N__73921));
    LocalMux I__16332 (
            .O(N__73921),
            .I(N__73918));
    Odrv12 I__16331 (
            .O(N__73918),
            .I(\pid_side.m11_2_03_3_i_0_o2_1 ));
    InMux I__16330 (
            .O(N__73915),
            .I(N__73912));
    LocalMux I__16329 (
            .O(N__73912),
            .I(N__73909));
    Span4Mux_s1_h I__16328 (
            .O(N__73909),
            .I(N__73903));
    InMux I__16327 (
            .O(N__73908),
            .I(N__73900));
    InMux I__16326 (
            .O(N__73907),
            .I(N__73888));
    InMux I__16325 (
            .O(N__73906),
            .I(N__73888));
    Span4Mux_h I__16324 (
            .O(N__73903),
            .I(N__73884));
    LocalMux I__16323 (
            .O(N__73900),
            .I(N__73881));
    InMux I__16322 (
            .O(N__73899),
            .I(N__73876));
    InMux I__16321 (
            .O(N__73898),
            .I(N__73876));
    InMux I__16320 (
            .O(N__73897),
            .I(N__73873));
    InMux I__16319 (
            .O(N__73896),
            .I(N__73864));
    InMux I__16318 (
            .O(N__73895),
            .I(N__73864));
    InMux I__16317 (
            .O(N__73894),
            .I(N__73864));
    InMux I__16316 (
            .O(N__73893),
            .I(N__73864));
    LocalMux I__16315 (
            .O(N__73888),
            .I(N__73861));
    InMux I__16314 (
            .O(N__73887),
            .I(N__73857));
    Span4Mux_h I__16313 (
            .O(N__73884),
            .I(N__73854));
    Span4Mux_h I__16312 (
            .O(N__73881),
            .I(N__73851));
    LocalMux I__16311 (
            .O(N__73876),
            .I(N__73848));
    LocalMux I__16310 (
            .O(N__73873),
            .I(N__73845));
    LocalMux I__16309 (
            .O(N__73864),
            .I(N__73840));
    Span4Mux_v I__16308 (
            .O(N__73861),
            .I(N__73840));
    InMux I__16307 (
            .O(N__73860),
            .I(N__73837));
    LocalMux I__16306 (
            .O(N__73857),
            .I(N__73834));
    Span4Mux_h I__16305 (
            .O(N__73854),
            .I(N__73831));
    Span4Mux_h I__16304 (
            .O(N__73851),
            .I(N__73828));
    Span4Mux_v I__16303 (
            .O(N__73848),
            .I(N__73825));
    Span4Mux_v I__16302 (
            .O(N__73845),
            .I(N__73820));
    Span4Mux_h I__16301 (
            .O(N__73840),
            .I(N__73820));
    LocalMux I__16300 (
            .O(N__73837),
            .I(N__73815));
    Span4Mux_v I__16299 (
            .O(N__73834),
            .I(N__73815));
    Span4Mux_v I__16298 (
            .O(N__73831),
            .I(N__73810));
    Span4Mux_h I__16297 (
            .O(N__73828),
            .I(N__73810));
    Odrv4 I__16296 (
            .O(N__73825),
            .I(\pid_front.error_13 ));
    Odrv4 I__16295 (
            .O(N__73820),
            .I(\pid_front.error_13 ));
    Odrv4 I__16294 (
            .O(N__73815),
            .I(\pid_front.error_13 ));
    Odrv4 I__16293 (
            .O(N__73810),
            .I(\pid_front.error_13 ));
    InMux I__16292 (
            .O(N__73801),
            .I(N__73798));
    LocalMux I__16291 (
            .O(N__73798),
            .I(N__73790));
    InMux I__16290 (
            .O(N__73797),
            .I(N__73787));
    InMux I__16289 (
            .O(N__73796),
            .I(N__73782));
    InMux I__16288 (
            .O(N__73795),
            .I(N__73782));
    InMux I__16287 (
            .O(N__73794),
            .I(N__73779));
    CascadeMux I__16286 (
            .O(N__73793),
            .I(N__73776));
    Span4Mux_v I__16285 (
            .O(N__73790),
            .I(N__73773));
    LocalMux I__16284 (
            .O(N__73787),
            .I(N__73770));
    LocalMux I__16283 (
            .O(N__73782),
            .I(N__73766));
    LocalMux I__16282 (
            .O(N__73779),
            .I(N__73763));
    InMux I__16281 (
            .O(N__73776),
            .I(N__73760));
    Span4Mux_h I__16280 (
            .O(N__73773),
            .I(N__73757));
    Span4Mux_h I__16279 (
            .O(N__73770),
            .I(N__73754));
    InMux I__16278 (
            .O(N__73769),
            .I(N__73751));
    Span4Mux_h I__16277 (
            .O(N__73766),
            .I(N__73744));
    Span4Mux_v I__16276 (
            .O(N__73763),
            .I(N__73744));
    LocalMux I__16275 (
            .O(N__73760),
            .I(N__73744));
    Span4Mux_h I__16274 (
            .O(N__73757),
            .I(N__73741));
    Span4Mux_h I__16273 (
            .O(N__73754),
            .I(N__73738));
    LocalMux I__16272 (
            .O(N__73751),
            .I(N__73735));
    Span4Mux_h I__16271 (
            .O(N__73744),
            .I(N__73732));
    Span4Mux_h I__16270 (
            .O(N__73741),
            .I(N__73729));
    Span4Mux_h I__16269 (
            .O(N__73738),
            .I(N__73726));
    Odrv12 I__16268 (
            .O(N__73735),
            .I(\pid_front.error_9 ));
    Odrv4 I__16267 (
            .O(N__73732),
            .I(\pid_front.error_9 ));
    Odrv4 I__16266 (
            .O(N__73729),
            .I(\pid_front.error_9 ));
    Odrv4 I__16265 (
            .O(N__73726),
            .I(\pid_front.error_9 ));
    InMux I__16264 (
            .O(N__73717),
            .I(N__73714));
    LocalMux I__16263 (
            .O(N__73714),
            .I(N__73710));
    InMux I__16262 (
            .O(N__73713),
            .I(N__73707));
    Odrv4 I__16261 (
            .O(N__73710),
            .I(\pid_side.N_185 ));
    LocalMux I__16260 (
            .O(N__73707),
            .I(\pid_side.N_185 ));
    InMux I__16259 (
            .O(N__73702),
            .I(N__73699));
    LocalMux I__16258 (
            .O(N__73699),
            .I(N__73695));
    InMux I__16257 (
            .O(N__73698),
            .I(N__73692));
    Odrv4 I__16256 (
            .O(N__73695),
            .I(\pid_side.N_207 ));
    LocalMux I__16255 (
            .O(N__73692),
            .I(\pid_side.N_207 ));
    InMux I__16254 (
            .O(N__73687),
            .I(N__73681));
    InMux I__16253 (
            .O(N__73686),
            .I(N__73681));
    LocalMux I__16252 (
            .O(N__73681),
            .I(N__73678));
    Odrv4 I__16251 (
            .O(N__73678),
            .I(\pid_side.m10_2_03_3_i_0_o2_1 ));
    CascadeMux I__16250 (
            .O(N__73675),
            .I(N__73672));
    InMux I__16249 (
            .O(N__73672),
            .I(N__73669));
    LocalMux I__16248 (
            .O(N__73669),
            .I(N__73666));
    Span4Mux_v I__16247 (
            .O(N__73666),
            .I(N__73663));
    Span4Mux_v I__16246 (
            .O(N__73663),
            .I(N__73660));
    Odrv4 I__16245 (
            .O(N__73660),
            .I(\pid_front.m78_0_a2_sx ));
    InMux I__16244 (
            .O(N__73657),
            .I(N__73654));
    LocalMux I__16243 (
            .O(N__73654),
            .I(N__73650));
    InMux I__16242 (
            .O(N__73653),
            .I(N__73647));
    Span4Mux_h I__16241 (
            .O(N__73650),
            .I(N__73642));
    LocalMux I__16240 (
            .O(N__73647),
            .I(N__73642));
    Span4Mux_v I__16239 (
            .O(N__73642),
            .I(N__73639));
    Odrv4 I__16238 (
            .O(N__73639),
            .I(\pid_front.N_524 ));
    CascadeMux I__16237 (
            .O(N__73636),
            .I(\pid_front.error_cry_1_c_RNIJE4MZ0Z2_cascade_ ));
    CascadeMux I__16236 (
            .O(N__73633),
            .I(N__73628));
    InMux I__16235 (
            .O(N__73632),
            .I(N__73625));
    InMux I__16234 (
            .O(N__73631),
            .I(N__73622));
    InMux I__16233 (
            .O(N__73628),
            .I(N__73619));
    LocalMux I__16232 (
            .O(N__73625),
            .I(N__73616));
    LocalMux I__16231 (
            .O(N__73622),
            .I(\pid_front.N_182 ));
    LocalMux I__16230 (
            .O(N__73619),
            .I(\pid_front.N_182 ));
    Odrv12 I__16229 (
            .O(N__73616),
            .I(\pid_front.N_182 ));
    InMux I__16228 (
            .O(N__73609),
            .I(N__73606));
    LocalMux I__16227 (
            .O(N__73606),
            .I(N__73603));
    Odrv4 I__16226 (
            .O(N__73603),
            .I(\pid_front.m8_2_03_3_i_0 ));
    CascadeMux I__16225 (
            .O(N__73600),
            .I(\pid_front.m8_2_03_3_i_0_cascade_ ));
    InMux I__16224 (
            .O(N__73597),
            .I(N__73594));
    LocalMux I__16223 (
            .O(N__73594),
            .I(N__73590));
    InMux I__16222 (
            .O(N__73593),
            .I(N__73587));
    Span4Mux_v I__16221 (
            .O(N__73590),
            .I(N__73584));
    LocalMux I__16220 (
            .O(N__73587),
            .I(\pid_front.error_i_regZ0Z_4 ));
    Odrv4 I__16219 (
            .O(N__73584),
            .I(\pid_front.error_i_regZ0Z_4 ));
    InMux I__16218 (
            .O(N__73579),
            .I(N__73576));
    LocalMux I__16217 (
            .O(N__73576),
            .I(N__73573));
    Odrv4 I__16216 (
            .O(N__73573),
            .I(\pid_front.m58_0_o2_N_2LZ0Z1 ));
    CascadeMux I__16215 (
            .O(N__73570),
            .I(\pid_side.error_i_reg_9_1_26_cascade_ ));
    CascadeMux I__16214 (
            .O(N__73567),
            .I(N__73564));
    InMux I__16213 (
            .O(N__73564),
            .I(N__73561));
    LocalMux I__16212 (
            .O(N__73561),
            .I(N__73558));
    Span4Mux_h I__16211 (
            .O(N__73558),
            .I(N__73555));
    Span4Mux_h I__16210 (
            .O(N__73555),
            .I(N__73552));
    Odrv4 I__16209 (
            .O(N__73552),
            .I(\pid_side.error_i_regZ0Z_26 ));
    CascadeMux I__16208 (
            .O(N__73549),
            .I(\pid_side.m10_2_03_3_i_0_o2_1_1_cascade_ ));
    CascadeMux I__16207 (
            .O(N__73546),
            .I(N__73543));
    InMux I__16206 (
            .O(N__73543),
            .I(N__73537));
    InMux I__16205 (
            .O(N__73542),
            .I(N__73537));
    LocalMux I__16204 (
            .O(N__73537),
            .I(\pid_side.m51_0_o2_0 ));
    InMux I__16203 (
            .O(N__73534),
            .I(N__73531));
    LocalMux I__16202 (
            .O(N__73531),
            .I(\pid_side.N_228 ));
    CascadeMux I__16201 (
            .O(N__73528),
            .I(N__73525));
    InMux I__16200 (
            .O(N__73525),
            .I(N__73522));
    LocalMux I__16199 (
            .O(N__73522),
            .I(N__73519));
    Span4Mux_h I__16198 (
            .O(N__73519),
            .I(N__73516));
    Span4Mux_v I__16197 (
            .O(N__73516),
            .I(N__73513));
    Odrv4 I__16196 (
            .O(N__73513),
            .I(\pid_side.error_i_regZ0Z_10 ));
    CascadeMux I__16195 (
            .O(N__73510),
            .I(N__73507));
    InMux I__16194 (
            .O(N__73507),
            .I(N__73504));
    LocalMux I__16193 (
            .O(N__73504),
            .I(\pid_side.m10_2_03_3_i_3 ));
    CascadeMux I__16192 (
            .O(N__73501),
            .I(N__73498));
    InMux I__16191 (
            .O(N__73498),
            .I(N__73495));
    LocalMux I__16190 (
            .O(N__73495),
            .I(N__73492));
    Span4Mux_h I__16189 (
            .O(N__73492),
            .I(N__73489));
    Span4Mux_v I__16188 (
            .O(N__73489),
            .I(N__73486));
    Odrv4 I__16187 (
            .O(N__73486),
            .I(\pid_side.error_i_regZ0Z_22 ));
    InMux I__16186 (
            .O(N__73483),
            .I(N__73480));
    LocalMux I__16185 (
            .O(N__73480),
            .I(\pid_front.N_186_0 ));
    InMux I__16184 (
            .O(N__73477),
            .I(N__73474));
    LocalMux I__16183 (
            .O(N__73474),
            .I(\pid_front.error_i_reg_esr_RNO_5_0_12 ));
    CascadeMux I__16182 (
            .O(N__73471),
            .I(\pid_side.m10_2_03_3_i_0_o2_0_1_cascade_ ));
    CascadeMux I__16181 (
            .O(N__73468),
            .I(\pid_side.error_cry_2_0_c_RNI7C2SZ0_cascade_ ));
    InMux I__16180 (
            .O(N__73465),
            .I(N__73462));
    LocalMux I__16179 (
            .O(N__73462),
            .I(\pid_side.N_155 ));
    CascadeMux I__16178 (
            .O(N__73459),
            .I(\pid_side.error_cry_2_0_c_RNI7A6PZ0Z2_cascade_ ));
    InMux I__16177 (
            .O(N__73456),
            .I(N__73453));
    LocalMux I__16176 (
            .O(N__73453),
            .I(N__73450));
    Span12Mux_s6_v I__16175 (
            .O(N__73450),
            .I(N__73446));
    InMux I__16174 (
            .O(N__73449),
            .I(N__73443));
    Odrv12 I__16173 (
            .O(N__73446),
            .I(\pid_side.N_204 ));
    LocalMux I__16172 (
            .O(N__73443),
            .I(\pid_side.N_204 ));
    CascadeMux I__16171 (
            .O(N__73438),
            .I(\pid_side.N_204_cascade_ ));
    InMux I__16170 (
            .O(N__73435),
            .I(N__73432));
    LocalMux I__16169 (
            .O(N__73432),
            .I(N__73429));
    Span4Mux_h I__16168 (
            .O(N__73429),
            .I(N__73425));
    InMux I__16167 (
            .O(N__73428),
            .I(N__73422));
    Odrv4 I__16166 (
            .O(N__73425),
            .I(\pid_side.N_186 ));
    LocalMux I__16165 (
            .O(N__73422),
            .I(\pid_side.N_186 ));
    CascadeMux I__16164 (
            .O(N__73417),
            .I(\pid_side.g0_16_1_cascade_ ));
    CascadeMux I__16163 (
            .O(N__73414),
            .I(\pid_side.N_228_cascade_ ));
    InMux I__16162 (
            .O(N__73411),
            .I(N__73408));
    LocalMux I__16161 (
            .O(N__73408),
            .I(\pid_side.error_i_reg_esr_RNO_5Z0Z_17 ));
    InMux I__16160 (
            .O(N__73405),
            .I(N__73401));
    InMux I__16159 (
            .O(N__73404),
            .I(N__73398));
    LocalMux I__16158 (
            .O(N__73401),
            .I(N__73395));
    LocalMux I__16157 (
            .O(N__73398),
            .I(N__73390));
    Span4Mux_h I__16156 (
            .O(N__73395),
            .I(N__73390));
    Odrv4 I__16155 (
            .O(N__73390),
            .I(xy_ki_fast_fast_3));
    CascadeMux I__16154 (
            .O(N__73387),
            .I(N__73384));
    InMux I__16153 (
            .O(N__73384),
            .I(N__73380));
    CascadeMux I__16152 (
            .O(N__73383),
            .I(N__73376));
    LocalMux I__16151 (
            .O(N__73380),
            .I(N__73373));
    InMux I__16150 (
            .O(N__73379),
            .I(N__73368));
    InMux I__16149 (
            .O(N__73376),
            .I(N__73368));
    Span4Mux_v I__16148 (
            .O(N__73373),
            .I(N__73364));
    LocalMux I__16147 (
            .O(N__73368),
            .I(N__73361));
    InMux I__16146 (
            .O(N__73367),
            .I(N__73358));
    Span4Mux_h I__16145 (
            .O(N__73364),
            .I(N__73355));
    Span12Mux_v I__16144 (
            .O(N__73361),
            .I(N__73350));
    LocalMux I__16143 (
            .O(N__73358),
            .I(N__73350));
    Odrv4 I__16142 (
            .O(N__73355),
            .I(pid_side_N_235));
    Odrv12 I__16141 (
            .O(N__73350),
            .I(pid_side_N_235));
    CascadeMux I__16140 (
            .O(N__73345),
            .I(pid_side_N_235_cascade_));
    CascadeMux I__16139 (
            .O(N__73342),
            .I(\pid_side.m28_2_03_0_0_cascade_ ));
    CascadeMux I__16138 (
            .O(N__73339),
            .I(\pid_side.m28_2_03_0_cascade_ ));
    CascadeMux I__16137 (
            .O(N__73336),
            .I(\pid_side.error_i_reg_9_rn_0_24_cascade_ ));
    CascadeMux I__16136 (
            .O(N__73333),
            .I(N__73330));
    InMux I__16135 (
            .O(N__73330),
            .I(N__73327));
    LocalMux I__16134 (
            .O(N__73327),
            .I(N__73324));
    Span4Mux_h I__16133 (
            .O(N__73324),
            .I(N__73321));
    Odrv4 I__16132 (
            .O(N__73321),
            .I(\pid_side.error_i_regZ0Z_24 ));
    InMux I__16131 (
            .O(N__73318),
            .I(N__73315));
    LocalMux I__16130 (
            .O(N__73315),
            .I(N__73312));
    Span12Mux_s6_v I__16129 (
            .O(N__73312),
            .I(N__73308));
    InMux I__16128 (
            .O(N__73311),
            .I(N__73305));
    Odrv12 I__16127 (
            .O(N__73308),
            .I(\pid_side.m56_0_o2_0 ));
    LocalMux I__16126 (
            .O(N__73305),
            .I(\pid_side.m56_0_o2_0 ));
    CascadeMux I__16125 (
            .O(N__73300),
            .I(\pid_side.m56_0_o2_0_cascade_ ));
    InMux I__16124 (
            .O(N__73297),
            .I(N__73294));
    LocalMux I__16123 (
            .O(N__73294),
            .I(\pid_side.error_i_reg_9_sn_24 ));
    InMux I__16122 (
            .O(N__73291),
            .I(N__73288));
    LocalMux I__16121 (
            .O(N__73288),
            .I(N__73285));
    Span4Mux_v I__16120 (
            .O(N__73285),
            .I(N__73282));
    Odrv4 I__16119 (
            .O(N__73282),
            .I(\pid_front.m78_0_m2_1_ns_1 ));
    InMux I__16118 (
            .O(N__73279),
            .I(N__73276));
    LocalMux I__16117 (
            .O(N__73276),
            .I(N__73272));
    InMux I__16116 (
            .O(N__73275),
            .I(N__73269));
    Span4Mux_v I__16115 (
            .O(N__73272),
            .I(N__73266));
    LocalMux I__16114 (
            .O(N__73269),
            .I(N__73261));
    Span4Mux_h I__16113 (
            .O(N__73266),
            .I(N__73261));
    Odrv4 I__16112 (
            .O(N__73261),
            .I(pid_side_m27_2_03_0_a2_0_0));
    CascadeMux I__16111 (
            .O(N__73258),
            .I(\pid_side.N_253_cascade_ ));
    CascadeMux I__16110 (
            .O(N__73255),
            .I(\pid_side.m27_2_03_0_cascade_ ));
    InMux I__16109 (
            .O(N__73252),
            .I(N__73249));
    LocalMux I__16108 (
            .O(N__73249),
            .I(N__73246));
    Span4Mux_h I__16107 (
            .O(N__73246),
            .I(N__73243));
    Odrv4 I__16106 (
            .O(N__73243),
            .I(\pid_side.error_i_regZ0Z_23 ));
    InMux I__16105 (
            .O(N__73240),
            .I(N__73237));
    LocalMux I__16104 (
            .O(N__73237),
            .I(\pid_side.N_576 ));
    InMux I__16103 (
            .O(N__73234),
            .I(N__73231));
    LocalMux I__16102 (
            .O(N__73231),
            .I(N__73227));
    InMux I__16101 (
            .O(N__73230),
            .I(N__73224));
    Odrv4 I__16100 (
            .O(N__73227),
            .I(\pid_side.m11_2_03_3_i_3 ));
    LocalMux I__16099 (
            .O(N__73224),
            .I(\pid_side.m11_2_03_3_i_3 ));
    InMux I__16098 (
            .O(N__73219),
            .I(N__73216));
    LocalMux I__16097 (
            .O(N__73216),
            .I(N__73213));
    Span4Mux_h I__16096 (
            .O(N__73213),
            .I(N__73210));
    Odrv4 I__16095 (
            .O(N__73210),
            .I(\pid_side.error_i_reg_esr_RNO_3Z0Z_14 ));
    CascadeMux I__16094 (
            .O(N__73207),
            .I(pid_side_N_216_cascade_));
    CascadeMux I__16093 (
            .O(N__73204),
            .I(\pid_side.error_i_reg_esr_RNO_6Z0Z_17_cascade_ ));
    InMux I__16092 (
            .O(N__73201),
            .I(N__73198));
    LocalMux I__16091 (
            .O(N__73198),
            .I(\pid_side.m21_2_03_0_0 ));
    CascadeMux I__16090 (
            .O(N__73195),
            .I(\pid_side.m21_2_03_0_1_cascade_ ));
    InMux I__16089 (
            .O(N__73192),
            .I(N__73189));
    LocalMux I__16088 (
            .O(N__73189),
            .I(\pid_side.error_i_reg_esr_RNO_0_0_17 ));
    InMux I__16087 (
            .O(N__73186),
            .I(N__73183));
    LocalMux I__16086 (
            .O(N__73183),
            .I(\pid_side.error_p_reg_esr_RNI1VTC1Z0Z_9 ));
    InMux I__16085 (
            .O(N__73180),
            .I(N__73177));
    LocalMux I__16084 (
            .O(N__73177),
            .I(N__73172));
    InMux I__16083 (
            .O(N__73176),
            .I(N__73167));
    InMux I__16082 (
            .O(N__73175),
            .I(N__73167));
    Span4Mux_v I__16081 (
            .O(N__73172),
            .I(N__73164));
    LocalMux I__16080 (
            .O(N__73167),
            .I(N__73161));
    Odrv4 I__16079 (
            .O(N__73164),
            .I(\pid_side.error_i_reg_esr_RNI6OOIZ0Z_10 ));
    Odrv4 I__16078 (
            .O(N__73161),
            .I(\pid_side.error_i_reg_esr_RNI6OOIZ0Z_10 ));
    CascadeMux I__16077 (
            .O(N__73156),
            .I(N__73153));
    InMux I__16076 (
            .O(N__73153),
            .I(N__73149));
    InMux I__16075 (
            .O(N__73152),
            .I(N__73146));
    LocalMux I__16074 (
            .O(N__73149),
            .I(N__73143));
    LocalMux I__16073 (
            .O(N__73146),
            .I(N__73140));
    Span4Mux_v I__16072 (
            .O(N__73143),
            .I(N__73137));
    Span4Mux_v I__16071 (
            .O(N__73140),
            .I(N__73134));
    Span4Mux_h I__16070 (
            .O(N__73137),
            .I(N__73131));
    Span4Mux_v I__16069 (
            .O(N__73134),
            .I(N__73128));
    Odrv4 I__16068 (
            .O(N__73131),
            .I(\pid_side.error_d_reg_prev_esr_RNITU3P4_0Z0Z_10 ));
    Odrv4 I__16067 (
            .O(N__73128),
            .I(\pid_side.error_d_reg_prev_esr_RNITU3P4_0Z0Z_10 ));
    InMux I__16066 (
            .O(N__73123),
            .I(N__73117));
    InMux I__16065 (
            .O(N__73122),
            .I(N__73117));
    LocalMux I__16064 (
            .O(N__73117),
            .I(\pid_side.error_p_reg_esr_RNIRE1B1Z0Z_10 ));
    CascadeMux I__16063 (
            .O(N__73114),
            .I(N__73111));
    InMux I__16062 (
            .O(N__73111),
            .I(N__73108));
    LocalMux I__16061 (
            .O(N__73108),
            .I(N__73105));
    Span4Mux_h I__16060 (
            .O(N__73105),
            .I(N__73102));
    Odrv4 I__16059 (
            .O(N__73102),
            .I(\pid_side.error_p_reg_esr_RNIV4S38Z0Z_10 ));
    InMux I__16058 (
            .O(N__73099),
            .I(N__73093));
    InMux I__16057 (
            .O(N__73098),
            .I(N__73090));
    InMux I__16056 (
            .O(N__73097),
            .I(N__73085));
    InMux I__16055 (
            .O(N__73096),
            .I(N__73085));
    LocalMux I__16054 (
            .O(N__73093),
            .I(\pid_side.error_d_reg_prevZ0Z_9 ));
    LocalMux I__16053 (
            .O(N__73090),
            .I(\pid_side.error_d_reg_prevZ0Z_9 ));
    LocalMux I__16052 (
            .O(N__73085),
            .I(\pid_side.error_d_reg_prevZ0Z_9 ));
    CascadeMux I__16051 (
            .O(N__73078),
            .I(N__73074));
    InMux I__16050 (
            .O(N__73077),
            .I(N__73070));
    InMux I__16049 (
            .O(N__73074),
            .I(N__73065));
    InMux I__16048 (
            .O(N__73073),
            .I(N__73065));
    LocalMux I__16047 (
            .O(N__73070),
            .I(N__73059));
    LocalMux I__16046 (
            .O(N__73065),
            .I(N__73059));
    InMux I__16045 (
            .O(N__73064),
            .I(N__73056));
    Odrv4 I__16044 (
            .O(N__73059),
            .I(\pid_side.error_d_reg_prevZ0Z_10 ));
    LocalMux I__16043 (
            .O(N__73056),
            .I(\pid_side.error_d_reg_prevZ0Z_10 ));
    InMux I__16042 (
            .O(N__73051),
            .I(N__73048));
    LocalMux I__16041 (
            .O(N__73048),
            .I(N__73045));
    Span4Mux_h I__16040 (
            .O(N__73045),
            .I(N__73042));
    Span4Mux_v I__16039 (
            .O(N__73042),
            .I(N__73039));
    Span4Mux_h I__16038 (
            .O(N__73039),
            .I(N__73036));
    Odrv4 I__16037 (
            .O(N__73036),
            .I(\pid_side.O_1_13 ));
    CascadeMux I__16036 (
            .O(N__73033),
            .I(N__73026));
    InMux I__16035 (
            .O(N__73032),
            .I(N__73020));
    InMux I__16034 (
            .O(N__73031),
            .I(N__73020));
    InMux I__16033 (
            .O(N__73030),
            .I(N__73011));
    InMux I__16032 (
            .O(N__73029),
            .I(N__73011));
    InMux I__16031 (
            .O(N__73026),
            .I(N__73011));
    InMux I__16030 (
            .O(N__73025),
            .I(N__73011));
    LocalMux I__16029 (
            .O(N__73020),
            .I(\pid_side.error_d_regZ0Z_10 ));
    LocalMux I__16028 (
            .O(N__73011),
            .I(\pid_side.error_d_regZ0Z_10 ));
    InMux I__16027 (
            .O(N__73006),
            .I(N__73003));
    LocalMux I__16026 (
            .O(N__73003),
            .I(N__73000));
    Span4Mux_h I__16025 (
            .O(N__73000),
            .I(N__72997));
    Span4Mux_h I__16024 (
            .O(N__72997),
            .I(N__72994));
    Odrv4 I__16023 (
            .O(N__72994),
            .I(\pid_side.O_2_14 ));
    CascadeMux I__16022 (
            .O(N__72991),
            .I(N__72986));
    InMux I__16021 (
            .O(N__72990),
            .I(N__72983));
    InMux I__16020 (
            .O(N__72989),
            .I(N__72978));
    InMux I__16019 (
            .O(N__72986),
            .I(N__72978));
    LocalMux I__16018 (
            .O(N__72983),
            .I(\pid_side.error_p_regZ0Z_10 ));
    LocalMux I__16017 (
            .O(N__72978),
            .I(\pid_side.error_p_regZ0Z_10 ));
    CascadeMux I__16016 (
            .O(N__72973),
            .I(\pid_front.m19_2_03_0_0_1_cascade_ ));
    InMux I__16015 (
            .O(N__72970),
            .I(N__72967));
    LocalMux I__16014 (
            .O(N__72967),
            .I(N__72964));
    Span4Mux_h I__16013 (
            .O(N__72964),
            .I(N__72960));
    InMux I__16012 (
            .O(N__72963),
            .I(N__72957));
    Odrv4 I__16011 (
            .O(N__72960),
            .I(\pid_front.N_161 ));
    LocalMux I__16010 (
            .O(N__72957),
            .I(\pid_front.N_161 ));
    CascadeMux I__16009 (
            .O(N__72952),
            .I(N__72944));
    CascadeMux I__16008 (
            .O(N__72951),
            .I(N__72941));
    CascadeMux I__16007 (
            .O(N__72950),
            .I(N__72937));
    CascadeMux I__16006 (
            .O(N__72949),
            .I(N__72934));
    CascadeMux I__16005 (
            .O(N__72948),
            .I(N__72931));
    CascadeMux I__16004 (
            .O(N__72947),
            .I(N__72920));
    InMux I__16003 (
            .O(N__72944),
            .I(N__72917));
    InMux I__16002 (
            .O(N__72941),
            .I(N__72914));
    InMux I__16001 (
            .O(N__72940),
            .I(N__72909));
    InMux I__16000 (
            .O(N__72937),
            .I(N__72909));
    InMux I__15999 (
            .O(N__72934),
            .I(N__72904));
    InMux I__15998 (
            .O(N__72931),
            .I(N__72904));
    CascadeMux I__15997 (
            .O(N__72930),
            .I(N__72901));
    InMux I__15996 (
            .O(N__72929),
            .I(N__72896));
    InMux I__15995 (
            .O(N__72928),
            .I(N__72896));
    CascadeMux I__15994 (
            .O(N__72927),
            .I(N__72893));
    CascadeMux I__15993 (
            .O(N__72926),
            .I(N__72890));
    CascadeMux I__15992 (
            .O(N__72925),
            .I(N__72887));
    InMux I__15991 (
            .O(N__72924),
            .I(N__72880));
    InMux I__15990 (
            .O(N__72923),
            .I(N__72880));
    InMux I__15989 (
            .O(N__72920),
            .I(N__72880));
    LocalMux I__15988 (
            .O(N__72917),
            .I(N__72875));
    LocalMux I__15987 (
            .O(N__72914),
            .I(N__72875));
    LocalMux I__15986 (
            .O(N__72909),
            .I(N__72870));
    LocalMux I__15985 (
            .O(N__72904),
            .I(N__72870));
    InMux I__15984 (
            .O(N__72901),
            .I(N__72867));
    LocalMux I__15983 (
            .O(N__72896),
            .I(N__72864));
    InMux I__15982 (
            .O(N__72893),
            .I(N__72857));
    InMux I__15981 (
            .O(N__72890),
            .I(N__72857));
    InMux I__15980 (
            .O(N__72887),
            .I(N__72857));
    LocalMux I__15979 (
            .O(N__72880),
            .I(N__72854));
    Span4Mux_h I__15978 (
            .O(N__72875),
            .I(N__72849));
    Span4Mux_h I__15977 (
            .O(N__72870),
            .I(N__72849));
    LocalMux I__15976 (
            .O(N__72867),
            .I(N__72844));
    Span4Mux_v I__15975 (
            .O(N__72864),
            .I(N__72844));
    LocalMux I__15974 (
            .O(N__72857),
            .I(\pid_side.error_d_reg_prevZ0Z_21 ));
    Odrv4 I__15973 (
            .O(N__72854),
            .I(\pid_side.error_d_reg_prevZ0Z_21 ));
    Odrv4 I__15972 (
            .O(N__72849),
            .I(\pid_side.error_d_reg_prevZ0Z_21 ));
    Odrv4 I__15971 (
            .O(N__72844),
            .I(\pid_side.error_d_reg_prevZ0Z_21 ));
    CascadeMux I__15970 (
            .O(N__72835),
            .I(N__72832));
    InMux I__15969 (
            .O(N__72832),
            .I(N__72825));
    InMux I__15968 (
            .O(N__72831),
            .I(N__72825));
    InMux I__15967 (
            .O(N__72830),
            .I(N__72822));
    LocalMux I__15966 (
            .O(N__72825),
            .I(N__72819));
    LocalMux I__15965 (
            .O(N__72822),
            .I(\pid_side.error_d_reg_prevZ0Z_8 ));
    Odrv4 I__15964 (
            .O(N__72819),
            .I(\pid_side.error_d_reg_prevZ0Z_8 ));
    CascadeMux I__15963 (
            .O(N__72814),
            .I(N__72811));
    InMux I__15962 (
            .O(N__72811),
            .I(N__72807));
    InMux I__15961 (
            .O(N__72810),
            .I(N__72804));
    LocalMux I__15960 (
            .O(N__72807),
            .I(N__72801));
    LocalMux I__15959 (
            .O(N__72804),
            .I(N__72798));
    Span4Mux_h I__15958 (
            .O(N__72801),
            .I(N__72795));
    Odrv12 I__15957 (
            .O(N__72798),
            .I(\pid_side.error_p_reg_esr_RNI9GJD3Z0Z_8 ));
    Odrv4 I__15956 (
            .O(N__72795),
            .I(\pid_side.error_p_reg_esr_RNI9GJD3Z0Z_8 ));
    CascadeMux I__15955 (
            .O(N__72790),
            .I(\pid_side.error_p_reg_esr_RNI1VTC1Z0Z_9_cascade_ ));
    InMux I__15954 (
            .O(N__72787),
            .I(N__72784));
    LocalMux I__15953 (
            .O(N__72784),
            .I(N__72781));
    Span4Mux_h I__15952 (
            .O(N__72781),
            .I(N__72778));
    Odrv4 I__15951 (
            .O(N__72778),
            .I(\pid_side.error_p_reg_esr_RNIBMBO6Z0Z_10 ));
    CascadeMux I__15950 (
            .O(N__72775),
            .I(\pid_side.N_2589_i_cascade_ ));
    InMux I__15949 (
            .O(N__72772),
            .I(N__72768));
    InMux I__15948 (
            .O(N__72771),
            .I(N__72765));
    LocalMux I__15947 (
            .O(N__72768),
            .I(N__72762));
    LocalMux I__15946 (
            .O(N__72765),
            .I(\pid_side.N_2583_i ));
    Odrv4 I__15945 (
            .O(N__72762),
            .I(\pid_side.N_2583_i ));
    InMux I__15944 (
            .O(N__72757),
            .I(N__72751));
    InMux I__15943 (
            .O(N__72756),
            .I(N__72751));
    LocalMux I__15942 (
            .O(N__72751),
            .I(N__72745));
    InMux I__15941 (
            .O(N__72750),
            .I(N__72738));
    InMux I__15940 (
            .O(N__72749),
            .I(N__72738));
    InMux I__15939 (
            .O(N__72748),
            .I(N__72738));
    Odrv4 I__15938 (
            .O(N__72745),
            .I(\pid_side.un1_pid_prereg_0_25 ));
    LocalMux I__15937 (
            .O(N__72738),
            .I(\pid_side.un1_pid_prereg_0_25 ));
    CascadeMux I__15936 (
            .O(N__72733),
            .I(\pid_side.un1_pid_prereg_0_25_cascade_ ));
    CascadeMux I__15935 (
            .O(N__72730),
            .I(N__72727));
    InMux I__15934 (
            .O(N__72727),
            .I(N__72723));
    InMux I__15933 (
            .O(N__72726),
            .I(N__72720));
    LocalMux I__15932 (
            .O(N__72723),
            .I(\pid_side.un1_pid_prereg_0_24 ));
    LocalMux I__15931 (
            .O(N__72720),
            .I(\pid_side.un1_pid_prereg_0_24 ));
    CascadeMux I__15930 (
            .O(N__72715),
            .I(N__72712));
    InMux I__15929 (
            .O(N__72712),
            .I(N__72709));
    LocalMux I__15928 (
            .O(N__72709),
            .I(N__72706));
    Odrv4 I__15927 (
            .O(N__72706),
            .I(\pid_side.error_d_reg_prev_esr_RNITP9B3Z0Z_21 ));
    InMux I__15926 (
            .O(N__72703),
            .I(N__72699));
    CascadeMux I__15925 (
            .O(N__72702),
            .I(N__72696));
    LocalMux I__15924 (
            .O(N__72699),
            .I(N__72693));
    InMux I__15923 (
            .O(N__72696),
            .I(N__72690));
    Span4Mux_v I__15922 (
            .O(N__72693),
            .I(N__72685));
    LocalMux I__15921 (
            .O(N__72690),
            .I(N__72685));
    Span4Mux_h I__15920 (
            .O(N__72685),
            .I(N__72682));
    Odrv4 I__15919 (
            .O(N__72682),
            .I(\pid_side.un1_pid_prereg_0 ));
    InMux I__15918 (
            .O(N__72679),
            .I(N__72676));
    LocalMux I__15917 (
            .O(N__72676),
            .I(N__72673));
    Sp12to4 I__15916 (
            .O(N__72673),
            .I(N__72670));
    Span12Mux_s6_v I__15915 (
            .O(N__72670),
            .I(N__72667));
    Odrv12 I__15914 (
            .O(N__72667),
            .I(\pid_side.error_d_reg_prev_esr_RNIHEJ01Z0Z_0 ));
    InMux I__15913 (
            .O(N__72664),
            .I(N__72661));
    LocalMux I__15912 (
            .O(N__72661),
            .I(N__72656));
    InMux I__15911 (
            .O(N__72660),
            .I(N__72653));
    InMux I__15910 (
            .O(N__72659),
            .I(N__72650));
    Span4Mux_h I__15909 (
            .O(N__72656),
            .I(N__72647));
    LocalMux I__15908 (
            .O(N__72653),
            .I(\pid_side.error_i_reg_esr_RNISESSZ0Z_25 ));
    LocalMux I__15907 (
            .O(N__72650),
            .I(\pid_side.error_i_reg_esr_RNISESSZ0Z_25 ));
    Odrv4 I__15906 (
            .O(N__72647),
            .I(\pid_side.error_i_reg_esr_RNISESSZ0Z_25 ));
    InMux I__15905 (
            .O(N__72640),
            .I(N__72637));
    LocalMux I__15904 (
            .O(N__72637),
            .I(N__72634));
    Span4Mux_h I__15903 (
            .O(N__72634),
            .I(N__72631));
    Span4Mux_v I__15902 (
            .O(N__72631),
            .I(N__72626));
    InMux I__15901 (
            .O(N__72630),
            .I(N__72621));
    InMux I__15900 (
            .O(N__72629),
            .I(N__72621));
    Odrv4 I__15899 (
            .O(N__72626),
            .I(\pid_side.un1_pid_prereg_0_19 ));
    LocalMux I__15898 (
            .O(N__72621),
            .I(\pid_side.un1_pid_prereg_0_19 ));
    CascadeMux I__15897 (
            .O(N__72616),
            .I(N__72612));
    CascadeMux I__15896 (
            .O(N__72615),
            .I(N__72609));
    InMux I__15895 (
            .O(N__72612),
            .I(N__72604));
    InMux I__15894 (
            .O(N__72609),
            .I(N__72604));
    LocalMux I__15893 (
            .O(N__72604),
            .I(N__72600));
    InMux I__15892 (
            .O(N__72603),
            .I(N__72597));
    Span4Mux_h I__15891 (
            .O(N__72600),
            .I(N__72594));
    LocalMux I__15890 (
            .O(N__72597),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_27_c_RNI1NVS ));
    Odrv4 I__15889 (
            .O(N__72594),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_27_c_RNI1NVS ));
    CascadeMux I__15888 (
            .O(N__72589),
            .I(N__72586));
    InMux I__15887 (
            .O(N__72586),
            .I(N__72580));
    InMux I__15886 (
            .O(N__72585),
            .I(N__72580));
    LocalMux I__15885 (
            .O(N__72580),
            .I(N__72576));
    InMux I__15884 (
            .O(N__72579),
            .I(N__72573));
    Odrv4 I__15883 (
            .O(N__72576),
            .I(\pid_side.un1_pid_prereg_0_26 ));
    LocalMux I__15882 (
            .O(N__72573),
            .I(\pid_side.un1_pid_prereg_0_26 ));
    InMux I__15881 (
            .O(N__72568),
            .I(N__72562));
    InMux I__15880 (
            .O(N__72567),
            .I(N__72559));
    InMux I__15879 (
            .O(N__72566),
            .I(N__72556));
    InMux I__15878 (
            .O(N__72565),
            .I(N__72553));
    LocalMux I__15877 (
            .O(N__72562),
            .I(N__72550));
    LocalMux I__15876 (
            .O(N__72559),
            .I(N__72547));
    LocalMux I__15875 (
            .O(N__72556),
            .I(N__72544));
    LocalMux I__15874 (
            .O(N__72553),
            .I(N__72541));
    Span4Mux_h I__15873 (
            .O(N__72550),
            .I(N__72536));
    Span4Mux_v I__15872 (
            .O(N__72547),
            .I(N__72536));
    Span4Mux_v I__15871 (
            .O(N__72544),
            .I(N__72529));
    Span4Mux_v I__15870 (
            .O(N__72541),
            .I(N__72529));
    Span4Mux_v I__15869 (
            .O(N__72536),
            .I(N__72529));
    Odrv4 I__15868 (
            .O(N__72529),
            .I(\pid_side.error_i_reg_esr_RNIGRJRZ0Z_11 ));
    InMux I__15867 (
            .O(N__72526),
            .I(N__72521));
    InMux I__15866 (
            .O(N__72525),
            .I(N__72518));
    InMux I__15865 (
            .O(N__72524),
            .I(N__72515));
    LocalMux I__15864 (
            .O(N__72521),
            .I(N__72512));
    LocalMux I__15863 (
            .O(N__72518),
            .I(\pid_side.error_d_reg_prev_esr_RNID3GT3_0Z0Z_10 ));
    LocalMux I__15862 (
            .O(N__72515),
            .I(\pid_side.error_d_reg_prev_esr_RNID3GT3_0Z0Z_10 ));
    Odrv12 I__15861 (
            .O(N__72512),
            .I(\pid_side.error_d_reg_prev_esr_RNID3GT3_0Z0Z_10 ));
    CascadeMux I__15860 (
            .O(N__72505),
            .I(N__72502));
    InMux I__15859 (
            .O(N__72502),
            .I(N__72499));
    LocalMux I__15858 (
            .O(N__72499),
            .I(N__72496));
    Span4Mux_h I__15857 (
            .O(N__72496),
            .I(N__72493));
    Odrv4 I__15856 (
            .O(N__72493),
            .I(\pid_side.error_d_reg_prev_esr_RNITU3P4Z0Z_10 ));
    InMux I__15855 (
            .O(N__72490),
            .I(N__72484));
    InMux I__15854 (
            .O(N__72489),
            .I(N__72484));
    LocalMux I__15853 (
            .O(N__72484),
            .I(N__72481));
    Odrv4 I__15852 (
            .O(N__72481),
            .I(\pid_side.N_2571_i ));
    CascadeMux I__15851 (
            .O(N__72478),
            .I(N__72475));
    InMux I__15850 (
            .O(N__72475),
            .I(N__72469));
    InMux I__15849 (
            .O(N__72474),
            .I(N__72469));
    LocalMux I__15848 (
            .O(N__72469),
            .I(N__72465));
    InMux I__15847 (
            .O(N__72468),
            .I(N__72462));
    Odrv4 I__15846 (
            .O(N__72465),
            .I(\pid_side.error_d_reg_prevZ0Z_7 ));
    LocalMux I__15845 (
            .O(N__72462),
            .I(\pid_side.error_d_reg_prevZ0Z_7 ));
    InMux I__15844 (
            .O(N__72457),
            .I(N__72454));
    LocalMux I__15843 (
            .O(N__72454),
            .I(N__72451));
    Span4Mux_v I__15842 (
            .O(N__72451),
            .I(N__72448));
    Span4Mux_h I__15841 (
            .O(N__72448),
            .I(N__72445));
    Odrv4 I__15840 (
            .O(N__72445),
            .I(\pid_side.state_RNIL5IFZ0Z_0 ));
    InMux I__15839 (
            .O(N__72442),
            .I(N__72438));
    CascadeMux I__15838 (
            .O(N__72441),
            .I(N__72435));
    LocalMux I__15837 (
            .O(N__72438),
            .I(N__72432));
    InMux I__15836 (
            .O(N__72435),
            .I(N__72429));
    Odrv4 I__15835 (
            .O(N__72432),
            .I(\pid_side.error_p_reg_esr_RNI5SNH3Z0Z_7 ));
    LocalMux I__15834 (
            .O(N__72429),
            .I(\pid_side.error_p_reg_esr_RNI5SNH3Z0Z_7 ));
    CascadeMux I__15833 (
            .O(N__72424),
            .I(\pid_side.error_p_reg_esr_RNISPTC1Z0Z_8_cascade_ ));
    InMux I__15832 (
            .O(N__72421),
            .I(N__72418));
    LocalMux I__15831 (
            .O(N__72418),
            .I(N__72415));
    Span4Mux_h I__15830 (
            .O(N__72415),
            .I(N__72412));
    Odrv4 I__15829 (
            .O(N__72412),
            .I(\pid_side.error_p_reg_esr_RNIECBV6Z0Z_8 ));
    InMux I__15828 (
            .O(N__72409),
            .I(N__72402));
    InMux I__15827 (
            .O(N__72408),
            .I(N__72402));
    InMux I__15826 (
            .O(N__72407),
            .I(N__72399));
    LocalMux I__15825 (
            .O(N__72402),
            .I(N__72396));
    LocalMux I__15824 (
            .O(N__72399),
            .I(N__72393));
    Span4Mux_h I__15823 (
            .O(N__72396),
            .I(N__72390));
    Odrv4 I__15822 (
            .O(N__72393),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_8_c_RNICNNJ ));
    Odrv4 I__15821 (
            .O(N__72390),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_8_c_RNICNNJ ));
    CascadeMux I__15820 (
            .O(N__72385),
            .I(N__72382));
    InMux I__15819 (
            .O(N__72382),
            .I(N__72379));
    LocalMux I__15818 (
            .O(N__72379),
            .I(\pid_side.error_p_reg_esr_RNISPTC1Z0Z_8 ));
    InMux I__15817 (
            .O(N__72376),
            .I(N__72370));
    InMux I__15816 (
            .O(N__72375),
            .I(N__72370));
    LocalMux I__15815 (
            .O(N__72370),
            .I(\pid_side.error_p_reg_esr_RNI1VTC1_0Z0Z_9 ));
    InMux I__15814 (
            .O(N__72367),
            .I(N__72364));
    LocalMux I__15813 (
            .O(N__72364),
            .I(\pid_side.N_2577_i ));
    CascadeMux I__15812 (
            .O(N__72361),
            .I(\pid_side.N_2577_i_cascade_ ));
    InMux I__15811 (
            .O(N__72358),
            .I(N__72355));
    LocalMux I__15810 (
            .O(N__72355),
            .I(N__72352));
    Span4Mux_h I__15809 (
            .O(N__72352),
            .I(N__72348));
    InMux I__15808 (
            .O(N__72351),
            .I(N__72345));
    Odrv4 I__15807 (
            .O(N__72348),
            .I(\pid_side.error_p_reg_esr_RNISPTC1_0Z0Z_8 ));
    LocalMux I__15806 (
            .O(N__72345),
            .I(\pid_side.error_p_reg_esr_RNISPTC1_0Z0Z_8 ));
    CascadeMux I__15805 (
            .O(N__72340),
            .I(\pid_side.un1_pid_prereg_9_0_cascade_ ));
    InMux I__15804 (
            .O(N__72337),
            .I(N__72333));
    CascadeMux I__15803 (
            .O(N__72336),
            .I(N__72330));
    LocalMux I__15802 (
            .O(N__72333),
            .I(N__72326));
    InMux I__15801 (
            .O(N__72330),
            .I(N__72323));
    InMux I__15800 (
            .O(N__72329),
            .I(N__72320));
    Span4Mux_v I__15799 (
            .O(N__72326),
            .I(N__72315));
    LocalMux I__15798 (
            .O(N__72323),
            .I(N__72315));
    LocalMux I__15797 (
            .O(N__72320),
            .I(N__72310));
    Span4Mux_h I__15796 (
            .O(N__72315),
            .I(N__72310));
    Odrv4 I__15795 (
            .O(N__72310),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_0_c_RNITGKN ));
    InMux I__15794 (
            .O(N__72307),
            .I(N__72304));
    LocalMux I__15793 (
            .O(N__72304),
            .I(N__72301));
    Span4Mux_v I__15792 (
            .O(N__72301),
            .I(N__72298));
    Odrv4 I__15791 (
            .O(N__72298),
            .I(\pid_side.error_d_reg_prev_esr_RNIM6H42Z0Z_0 ));
    CascadeMux I__15790 (
            .O(N__72295),
            .I(\pid_side.N_2565_i_cascade_ ));
    InMux I__15789 (
            .O(N__72292),
            .I(N__72289));
    LocalMux I__15788 (
            .O(N__72289),
            .I(\pid_side.error_p_reg_esr_RNINKTC1_0Z0Z_7 ));
    InMux I__15787 (
            .O(N__72286),
            .I(N__72280));
    InMux I__15786 (
            .O(N__72285),
            .I(N__72280));
    LocalMux I__15785 (
            .O(N__72280),
            .I(\pid_side.error_p_reg_esr_RNIIFTC1Z0Z_6 ));
    CascadeMux I__15784 (
            .O(N__72277),
            .I(\pid_side.error_p_reg_esr_RNINKTC1_0Z0Z_7_cascade_ ));
    InMux I__15783 (
            .O(N__72274),
            .I(N__72267));
    InMux I__15782 (
            .O(N__72273),
            .I(N__72267));
    InMux I__15781 (
            .O(N__72272),
            .I(N__72264));
    LocalMux I__15780 (
            .O(N__72267),
            .I(N__72261));
    LocalMux I__15779 (
            .O(N__72264),
            .I(N__72256));
    Span4Mux_h I__15778 (
            .O(N__72261),
            .I(N__72256));
    Odrv4 I__15777 (
            .O(N__72256),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_6_c_RNI6FLJ ));
    InMux I__15776 (
            .O(N__72253),
            .I(N__72250));
    LocalMux I__15775 (
            .O(N__72250),
            .I(N__72247));
    Odrv12 I__15774 (
            .O(N__72247),
            .I(\pid_side.error_p_reg_esr_RNIFJGD3_0Z0Z_6 ));
    CascadeMux I__15773 (
            .O(N__72244),
            .I(N__72241));
    InMux I__15772 (
            .O(N__72241),
            .I(N__72231));
    InMux I__15771 (
            .O(N__72240),
            .I(N__72231));
    InMux I__15770 (
            .O(N__72239),
            .I(N__72231));
    InMux I__15769 (
            .O(N__72238),
            .I(N__72228));
    LocalMux I__15768 (
            .O(N__72231),
            .I(\pid_side.error_d_reg_prevZ0Z_6 ));
    LocalMux I__15767 (
            .O(N__72228),
            .I(\pid_side.error_d_reg_prevZ0Z_6 ));
    InMux I__15766 (
            .O(N__72223),
            .I(N__72220));
    LocalMux I__15765 (
            .O(N__72220),
            .I(\pid_side.error_p_reg_esr_RNINKTC1Z0Z_7 ));
    InMux I__15764 (
            .O(N__72217),
            .I(N__72213));
    InMux I__15763 (
            .O(N__72216),
            .I(N__72210));
    LocalMux I__15762 (
            .O(N__72213),
            .I(N__72207));
    LocalMux I__15761 (
            .O(N__72210),
            .I(\pid_side.error_p_reg_esr_RNIFJGD3Z0Z_6 ));
    Odrv4 I__15760 (
            .O(N__72207),
            .I(\pid_side.error_p_reg_esr_RNIFJGD3Z0Z_6 ));
    CascadeMux I__15759 (
            .O(N__72202),
            .I(\pid_side.error_p_reg_esr_RNINKTC1Z0Z_7_cascade_ ));
    InMux I__15758 (
            .O(N__72199),
            .I(N__72195));
    InMux I__15757 (
            .O(N__72198),
            .I(N__72192));
    LocalMux I__15756 (
            .O(N__72195),
            .I(N__72188));
    LocalMux I__15755 (
            .O(N__72192),
            .I(N__72185));
    InMux I__15754 (
            .O(N__72191),
            .I(N__72182));
    Span4Mux_v I__15753 (
            .O(N__72188),
            .I(N__72179));
    Span4Mux_v I__15752 (
            .O(N__72185),
            .I(N__72174));
    LocalMux I__15751 (
            .O(N__72182),
            .I(N__72174));
    Span4Mux_v I__15750 (
            .O(N__72179),
            .I(N__72171));
    Span4Mux_h I__15749 (
            .O(N__72174),
            .I(N__72168));
    Odrv4 I__15748 (
            .O(N__72171),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_7_c_RNIIDSN ));
    Odrv4 I__15747 (
            .O(N__72168),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_7_c_RNIIDSN ));
    CascadeMux I__15746 (
            .O(N__72163),
            .I(N__72160));
    InMux I__15745 (
            .O(N__72160),
            .I(N__72157));
    LocalMux I__15744 (
            .O(N__72157),
            .I(N__72154));
    Odrv4 I__15743 (
            .O(N__72154),
            .I(\pid_side.error_p_reg_esr_RNIKF8V6Z0Z_7 ));
    CascadeMux I__15742 (
            .O(N__72151),
            .I(N__72148));
    InMux I__15741 (
            .O(N__72148),
            .I(N__72145));
    LocalMux I__15740 (
            .O(N__72145),
            .I(N__72142));
    Span4Mux_v I__15739 (
            .O(N__72142),
            .I(N__72139));
    Odrv4 I__15738 (
            .O(N__72139),
            .I(\pid_side.error_i_regZ0Z_8 ));
    InMux I__15737 (
            .O(N__72136),
            .I(N__72133));
    LocalMux I__15736 (
            .O(N__72133),
            .I(N__72128));
    InMux I__15735 (
            .O(N__72132),
            .I(N__72125));
    CascadeMux I__15734 (
            .O(N__72131),
            .I(N__72122));
    Span4Mux_v I__15733 (
            .O(N__72128),
            .I(N__72119));
    LocalMux I__15732 (
            .O(N__72125),
            .I(N__72116));
    InMux I__15731 (
            .O(N__72122),
            .I(N__72113));
    Odrv4 I__15730 (
            .O(N__72119),
            .I(\pid_front.error_i_reg_esr_RNI4EFVZ0Z_23 ));
    Odrv4 I__15729 (
            .O(N__72116),
            .I(\pid_front.error_i_reg_esr_RNI4EFVZ0Z_23 ));
    LocalMux I__15728 (
            .O(N__72113),
            .I(\pid_front.error_i_reg_esr_RNI4EFVZ0Z_23 ));
    CascadeMux I__15727 (
            .O(N__72106),
            .I(N__72102));
    CascadeMux I__15726 (
            .O(N__72105),
            .I(N__72099));
    InMux I__15725 (
            .O(N__72102),
            .I(N__72094));
    InMux I__15724 (
            .O(N__72099),
            .I(N__72094));
    LocalMux I__15723 (
            .O(N__72094),
            .I(\pid_front.error_i_acumm_preregZ0Z_23 ));
    InMux I__15722 (
            .O(N__72091),
            .I(N__72088));
    LocalMux I__15721 (
            .O(N__72088),
            .I(N__72085));
    Span4Mux_h I__15720 (
            .O(N__72085),
            .I(N__72081));
    CascadeMux I__15719 (
            .O(N__72084),
            .I(N__72078));
    Span4Mux_h I__15718 (
            .O(N__72081),
            .I(N__72075));
    InMux I__15717 (
            .O(N__72078),
            .I(N__72072));
    Span4Mux_v I__15716 (
            .O(N__72075),
            .I(N__72069));
    LocalMux I__15715 (
            .O(N__72072),
            .I(N__72066));
    Odrv4 I__15714 (
            .O(N__72069),
            .I(\pid_front.error_p_reg_esr_RNI0GC61_0Z0Z_19 ));
    Odrv12 I__15713 (
            .O(N__72066),
            .I(\pid_front.error_p_reg_esr_RNI0GC61_0Z0Z_19 ));
    InMux I__15712 (
            .O(N__72061),
            .I(N__72058));
    LocalMux I__15711 (
            .O(N__72058),
            .I(N__72053));
    InMux I__15710 (
            .O(N__72057),
            .I(N__72048));
    InMux I__15709 (
            .O(N__72056),
            .I(N__72048));
    Span4Mux_h I__15708 (
            .O(N__72053),
            .I(N__72045));
    LocalMux I__15707 (
            .O(N__72048),
            .I(N__72042));
    Span4Mux_v I__15706 (
            .O(N__72045),
            .I(N__72037));
    Span4Mux_v I__15705 (
            .O(N__72042),
            .I(N__72037));
    Odrv4 I__15704 (
            .O(N__72037),
            .I(\pid_front.error_i_reg_esr_RNIERHUZ0Z_19 ));
    InMux I__15703 (
            .O(N__72034),
            .I(N__72030));
    InMux I__15702 (
            .O(N__72033),
            .I(N__72027));
    LocalMux I__15701 (
            .O(N__72030),
            .I(N__72024));
    LocalMux I__15700 (
            .O(N__72027),
            .I(N__72021));
    Odrv12 I__15699 (
            .O(N__72024),
            .I(\pid_front.un1_pid_prereg_0_7 ));
    Odrv4 I__15698 (
            .O(N__72021),
            .I(\pid_front.un1_pid_prereg_0_7 ));
    CascadeMux I__15697 (
            .O(N__72016),
            .I(\pid_front.un1_pid_prereg_0_7_cascade_ ));
    InMux I__15696 (
            .O(N__72013),
            .I(N__72009));
    InMux I__15695 (
            .O(N__72012),
            .I(N__72006));
    LocalMux I__15694 (
            .O(N__72009),
            .I(N__72003));
    LocalMux I__15693 (
            .O(N__72006),
            .I(N__72000));
    Odrv4 I__15692 (
            .O(N__72003),
            .I(\pid_front.un1_pid_prereg_0_6 ));
    Odrv4 I__15691 (
            .O(N__72000),
            .I(\pid_front.un1_pid_prereg_0_6 ));
    CascadeMux I__15690 (
            .O(N__71995),
            .I(N__71992));
    InMux I__15689 (
            .O(N__71992),
            .I(N__71989));
    LocalMux I__15688 (
            .O(N__71989),
            .I(N__71986));
    Span4Mux_h I__15687 (
            .O(N__71986),
            .I(N__71983));
    Odrv4 I__15686 (
            .O(N__71983),
            .I(\pid_front.error_p_reg_esr_RNIE7KM6Z0Z_17 ));
    CascadeMux I__15685 (
            .O(N__71980),
            .I(N__71977));
    InMux I__15684 (
            .O(N__71977),
            .I(N__71974));
    LocalMux I__15683 (
            .O(N__71974),
            .I(N__71971));
    Span4Mux_h I__15682 (
            .O(N__71971),
            .I(N__71965));
    InMux I__15681 (
            .O(N__71970),
            .I(N__71960));
    InMux I__15680 (
            .O(N__71969),
            .I(N__71960));
    InMux I__15679 (
            .O(N__71968),
            .I(N__71957));
    Odrv4 I__15678 (
            .O(N__71965),
            .I(\pid_front.error_d_reg_fastZ0Z_12 ));
    LocalMux I__15677 (
            .O(N__71960),
            .I(\pid_front.error_d_reg_fastZ0Z_12 ));
    LocalMux I__15676 (
            .O(N__71957),
            .I(\pid_front.error_d_reg_fastZ0Z_12 ));
    CascadeMux I__15675 (
            .O(N__71950),
            .I(N__71947));
    InMux I__15674 (
            .O(N__71947),
            .I(N__71940));
    InMux I__15673 (
            .O(N__71946),
            .I(N__71940));
    CascadeMux I__15672 (
            .O(N__71945),
            .I(N__71936));
    LocalMux I__15671 (
            .O(N__71940),
            .I(N__71932));
    InMux I__15670 (
            .O(N__71939),
            .I(N__71929));
    InMux I__15669 (
            .O(N__71936),
            .I(N__71924));
    InMux I__15668 (
            .O(N__71935),
            .I(N__71924));
    Odrv4 I__15667 (
            .O(N__71932),
            .I(\pid_front.error_p_regZ0Z_11 ));
    LocalMux I__15666 (
            .O(N__71929),
            .I(\pid_front.error_p_regZ0Z_11 ));
    LocalMux I__15665 (
            .O(N__71924),
            .I(\pid_front.error_p_regZ0Z_11 ));
    CascadeMux I__15664 (
            .O(N__71917),
            .I(\pid_front.g0_1_0_1_cascade_ ));
    CascadeMux I__15663 (
            .O(N__71914),
            .I(N__71909));
    CascadeMux I__15662 (
            .O(N__71913),
            .I(N__71906));
    CascadeMux I__15661 (
            .O(N__71912),
            .I(N__71899));
    InMux I__15660 (
            .O(N__71909),
            .I(N__71892));
    InMux I__15659 (
            .O(N__71906),
            .I(N__71892));
    InMux I__15658 (
            .O(N__71905),
            .I(N__71892));
    InMux I__15657 (
            .O(N__71904),
            .I(N__71889));
    InMux I__15656 (
            .O(N__71903),
            .I(N__71886));
    InMux I__15655 (
            .O(N__71902),
            .I(N__71881));
    InMux I__15654 (
            .O(N__71899),
            .I(N__71881));
    LocalMux I__15653 (
            .O(N__71892),
            .I(N__71878));
    LocalMux I__15652 (
            .O(N__71889),
            .I(\pid_front.error_p_regZ0Z_12 ));
    LocalMux I__15651 (
            .O(N__71886),
            .I(\pid_front.error_p_regZ0Z_12 ));
    LocalMux I__15650 (
            .O(N__71881),
            .I(\pid_front.error_p_regZ0Z_12 ));
    Odrv4 I__15649 (
            .O(N__71878),
            .I(\pid_front.error_p_regZ0Z_12 ));
    InMux I__15648 (
            .O(N__71869),
            .I(N__71866));
    LocalMux I__15647 (
            .O(N__71866),
            .I(\pid_front.g0_1 ));
    InMux I__15646 (
            .O(N__71863),
            .I(N__71860));
    LocalMux I__15645 (
            .O(N__71860),
            .I(N__71857));
    Odrv4 I__15644 (
            .O(N__71857),
            .I(\pid_front.N_5 ));
    InMux I__15643 (
            .O(N__71854),
            .I(N__71848));
    InMux I__15642 (
            .O(N__71853),
            .I(N__71848));
    LocalMux I__15641 (
            .O(N__71848),
            .I(N__71845));
    Span4Mux_h I__15640 (
            .O(N__71845),
            .I(N__71839));
    InMux I__15639 (
            .O(N__71844),
            .I(N__71836));
    InMux I__15638 (
            .O(N__71843),
            .I(N__71831));
    InMux I__15637 (
            .O(N__71842),
            .I(N__71831));
    Odrv4 I__15636 (
            .O(N__71839),
            .I(\pid_front.error_d_reg_prevZ0Z_11 ));
    LocalMux I__15635 (
            .O(N__71836),
            .I(\pid_front.error_d_reg_prevZ0Z_11 ));
    LocalMux I__15634 (
            .O(N__71831),
            .I(\pid_front.error_d_reg_prevZ0Z_11 ));
    CEMux I__15633 (
            .O(N__71824),
            .I(N__71821));
    LocalMux I__15632 (
            .O(N__71821),
            .I(N__71818));
    Span4Mux_v I__15631 (
            .O(N__71818),
            .I(N__71813));
    CEMux I__15630 (
            .O(N__71817),
            .I(N__71810));
    CEMux I__15629 (
            .O(N__71816),
            .I(N__71806));
    Span4Mux_h I__15628 (
            .O(N__71813),
            .I(N__71799));
    LocalMux I__15627 (
            .O(N__71810),
            .I(N__71799));
    CEMux I__15626 (
            .O(N__71809),
            .I(N__71796));
    LocalMux I__15625 (
            .O(N__71806),
            .I(N__71791));
    CEMux I__15624 (
            .O(N__71805),
            .I(N__71788));
    CEMux I__15623 (
            .O(N__71804),
            .I(N__71782));
    Span4Mux_h I__15622 (
            .O(N__71799),
            .I(N__71777));
    LocalMux I__15621 (
            .O(N__71796),
            .I(N__71777));
    CEMux I__15620 (
            .O(N__71795),
            .I(N__71774));
    CEMux I__15619 (
            .O(N__71794),
            .I(N__71771));
    Span4Mux_h I__15618 (
            .O(N__71791),
            .I(N__71766));
    LocalMux I__15617 (
            .O(N__71788),
            .I(N__71766));
    CEMux I__15616 (
            .O(N__71787),
            .I(N__71763));
    CEMux I__15615 (
            .O(N__71786),
            .I(N__71760));
    CEMux I__15614 (
            .O(N__71785),
            .I(N__71757));
    LocalMux I__15613 (
            .O(N__71782),
            .I(N__71748));
    Span4Mux_h I__15612 (
            .O(N__71777),
            .I(N__71748));
    LocalMux I__15611 (
            .O(N__71774),
            .I(N__71748));
    LocalMux I__15610 (
            .O(N__71771),
            .I(N__71748));
    Span4Mux_h I__15609 (
            .O(N__71766),
            .I(N__71742));
    LocalMux I__15608 (
            .O(N__71763),
            .I(N__71742));
    LocalMux I__15607 (
            .O(N__71760),
            .I(N__71739));
    LocalMux I__15606 (
            .O(N__71757),
            .I(N__71734));
    Span4Mux_v I__15605 (
            .O(N__71748),
            .I(N__71734));
    CEMux I__15604 (
            .O(N__71747),
            .I(N__71731));
    Span4Mux_v I__15603 (
            .O(N__71742),
            .I(N__71726));
    Span4Mux_h I__15602 (
            .O(N__71739),
            .I(N__71726));
    Span4Mux_h I__15601 (
            .O(N__71734),
            .I(N__71721));
    LocalMux I__15600 (
            .O(N__71731),
            .I(N__71721));
    Odrv4 I__15599 (
            .O(N__71726),
            .I(\pid_front.N_763_0 ));
    Odrv4 I__15598 (
            .O(N__71721),
            .I(\pid_front.N_763_0 ));
    SRMux I__15597 (
            .O(N__71716),
            .I(N__71711));
    SRMux I__15596 (
            .O(N__71715),
            .I(N__71708));
    SRMux I__15595 (
            .O(N__71714),
            .I(N__71701));
    LocalMux I__15594 (
            .O(N__71711),
            .I(N__71696));
    LocalMux I__15593 (
            .O(N__71708),
            .I(N__71693));
    SRMux I__15592 (
            .O(N__71707),
            .I(N__71690));
    SRMux I__15591 (
            .O(N__71706),
            .I(N__71687));
    SRMux I__15590 (
            .O(N__71705),
            .I(N__71684));
    SRMux I__15589 (
            .O(N__71704),
            .I(N__71680));
    LocalMux I__15588 (
            .O(N__71701),
            .I(N__71677));
    SRMux I__15587 (
            .O(N__71700),
            .I(N__71674));
    SRMux I__15586 (
            .O(N__71699),
            .I(N__71671));
    Span4Mux_v I__15585 (
            .O(N__71696),
            .I(N__71668));
    Span4Mux_h I__15584 (
            .O(N__71693),
            .I(N__71661));
    LocalMux I__15583 (
            .O(N__71690),
            .I(N__71661));
    LocalMux I__15582 (
            .O(N__71687),
            .I(N__71661));
    LocalMux I__15581 (
            .O(N__71684),
            .I(N__71658));
    SRMux I__15580 (
            .O(N__71683),
            .I(N__71655));
    LocalMux I__15579 (
            .O(N__71680),
            .I(N__71652));
    Span4Mux_v I__15578 (
            .O(N__71677),
            .I(N__71645));
    LocalMux I__15577 (
            .O(N__71674),
            .I(N__71645));
    LocalMux I__15576 (
            .O(N__71671),
            .I(N__71645));
    Span4Mux_h I__15575 (
            .O(N__71668),
            .I(N__71640));
    Span4Mux_v I__15574 (
            .O(N__71661),
            .I(N__71640));
    Span4Mux_v I__15573 (
            .O(N__71658),
            .I(N__71635));
    LocalMux I__15572 (
            .O(N__71655),
            .I(N__71635));
    Span4Mux_v I__15571 (
            .O(N__71652),
            .I(N__71630));
    Span4Mux_v I__15570 (
            .O(N__71645),
            .I(N__71630));
    Span4Mux_v I__15569 (
            .O(N__71640),
            .I(N__71624));
    Span4Mux_h I__15568 (
            .O(N__71635),
            .I(N__71621));
    Sp12to4 I__15567 (
            .O(N__71630),
            .I(N__71618));
    SRMux I__15566 (
            .O(N__71629),
            .I(N__71615));
    SRMux I__15565 (
            .O(N__71628),
            .I(N__71612));
    InMux I__15564 (
            .O(N__71627),
            .I(N__71609));
    Odrv4 I__15563 (
            .O(N__71624),
            .I(\pid_front.state_RNIM14NZ0Z_0 ));
    Odrv4 I__15562 (
            .O(N__71621),
            .I(\pid_front.state_RNIM14NZ0Z_0 ));
    Odrv12 I__15561 (
            .O(N__71618),
            .I(\pid_front.state_RNIM14NZ0Z_0 ));
    LocalMux I__15560 (
            .O(N__71615),
            .I(\pid_front.state_RNIM14NZ0Z_0 ));
    LocalMux I__15559 (
            .O(N__71612),
            .I(\pid_front.state_RNIM14NZ0Z_0 ));
    LocalMux I__15558 (
            .O(N__71609),
            .I(\pid_front.state_RNIM14NZ0Z_0 ));
    InMux I__15557 (
            .O(N__71596),
            .I(N__71592));
    CascadeMux I__15556 (
            .O(N__71595),
            .I(N__71589));
    LocalMux I__15555 (
            .O(N__71592),
            .I(N__71586));
    InMux I__15554 (
            .O(N__71589),
            .I(N__71583));
    Span4Mux_v I__15553 (
            .O(N__71586),
            .I(N__71580));
    LocalMux I__15552 (
            .O(N__71583),
            .I(N__71577));
    Span4Mux_v I__15551 (
            .O(N__71580),
            .I(N__71574));
    Span4Mux_h I__15550 (
            .O(N__71577),
            .I(N__71571));
    Odrv4 I__15549 (
            .O(N__71574),
            .I(\pid_front.error_p_reg_esr_RNIOH2JDZ0Z_12 ));
    Odrv4 I__15548 (
            .O(N__71571),
            .I(\pid_front.error_p_reg_esr_RNIOH2JDZ0Z_12 ));
    CascadeMux I__15547 (
            .O(N__71566),
            .I(\pid_front.error_p_reg_esr_RNIBJ5B3_0Z0Z_14_cascade_ ));
    InMux I__15546 (
            .O(N__71563),
            .I(N__71559));
    InMux I__15545 (
            .O(N__71562),
            .I(N__71556));
    LocalMux I__15544 (
            .O(N__71559),
            .I(N__71553));
    LocalMux I__15543 (
            .O(N__71556),
            .I(N__71549));
    Span4Mux_v I__15542 (
            .O(N__71553),
            .I(N__71546));
    InMux I__15541 (
            .O(N__71552),
            .I(N__71543));
    Span4Mux_h I__15540 (
            .O(N__71549),
            .I(N__71540));
    Span4Mux_v I__15539 (
            .O(N__71546),
            .I(N__71535));
    LocalMux I__15538 (
            .O(N__71543),
            .I(N__71535));
    Odrv4 I__15537 (
            .O(N__71540),
            .I(\pid_front.error_d_reg_prev_esr_RNI13Q1DZ0Z_12 ));
    Odrv4 I__15536 (
            .O(N__71535),
            .I(\pid_front.error_d_reg_prev_esr_RNI13Q1DZ0Z_12 ));
    InMux I__15535 (
            .O(N__71530),
            .I(N__71527));
    LocalMux I__15534 (
            .O(N__71527),
            .I(N__71524));
    Span4Mux_h I__15533 (
            .O(N__71524),
            .I(N__71521));
    Odrv4 I__15532 (
            .O(N__71521),
            .I(\pid_front.error_p_reg_esr_RNI4820UZ0Z_12 ));
    InMux I__15531 (
            .O(N__71518),
            .I(N__71515));
    LocalMux I__15530 (
            .O(N__71515),
            .I(\pid_front.error_i_acumm_13_i_o2_0_9_3 ));
    CascadeMux I__15529 (
            .O(N__71512),
            .I(N__71509));
    InMux I__15528 (
            .O(N__71509),
            .I(N__71506));
    LocalMux I__15527 (
            .O(N__71506),
            .I(N__71503));
    Span4Mux_v I__15526 (
            .O(N__71503),
            .I(N__71500));
    Odrv4 I__15525 (
            .O(N__71500),
            .I(\pid_front.error_i_acumm_13_i_o2_0_10_3 ));
    InMux I__15524 (
            .O(N__71497),
            .I(N__71494));
    LocalMux I__15523 (
            .O(N__71494),
            .I(N__71491));
    Span4Mux_v I__15522 (
            .O(N__71491),
            .I(N__71488));
    Odrv4 I__15521 (
            .O(N__71488),
            .I(\pid_front.error_i_acumm_13_i_o2_0_7_3 ));
    InMux I__15520 (
            .O(N__71485),
            .I(N__71482));
    LocalMux I__15519 (
            .O(N__71482),
            .I(\pid_front.error_i_acumm_13_i_o2_0_9_12 ));
    CascadeMux I__15518 (
            .O(N__71479),
            .I(N__71476));
    InMux I__15517 (
            .O(N__71476),
            .I(N__71473));
    LocalMux I__15516 (
            .O(N__71473),
            .I(N__71470));
    Span4Mux_h I__15515 (
            .O(N__71470),
            .I(N__71467));
    Odrv4 I__15514 (
            .O(N__71467),
            .I(\pid_front.error_i_acumm_13_i_o2_0_10_12 ));
    InMux I__15513 (
            .O(N__71464),
            .I(N__71461));
    LocalMux I__15512 (
            .O(N__71461),
            .I(N__71458));
    Odrv12 I__15511 (
            .O(N__71458),
            .I(\pid_front.error_i_acumm_13_i_o2_0_7_12 ));
    InMux I__15510 (
            .O(N__71455),
            .I(N__71452));
    LocalMux I__15509 (
            .O(N__71452),
            .I(\pid_front.error_i_acumm_13_i_o2_0_8_12 ));
    InMux I__15508 (
            .O(N__71449),
            .I(N__71443));
    InMux I__15507 (
            .O(N__71448),
            .I(N__71443));
    LocalMux I__15506 (
            .O(N__71443),
            .I(\pid_front.error_i_acumm_preregZ0Z_19 ));
    InMux I__15505 (
            .O(N__71440),
            .I(N__71437));
    LocalMux I__15504 (
            .O(N__71437),
            .I(\pid_front.error_i_acumm_13_i_o2_0_8_3 ));
    InMux I__15503 (
            .O(N__71434),
            .I(N__71429));
    InMux I__15502 (
            .O(N__71433),
            .I(N__71424));
    InMux I__15501 (
            .O(N__71432),
            .I(N__71424));
    LocalMux I__15500 (
            .O(N__71429),
            .I(N__71421));
    LocalMux I__15499 (
            .O(N__71424),
            .I(N__71418));
    Span4Mux_v I__15498 (
            .O(N__71421),
            .I(N__71415));
    Span4Mux_v I__15497 (
            .O(N__71418),
            .I(N__71412));
    Odrv4 I__15496 (
            .O(N__71415),
            .I(\pid_front.error_i_reg_esr_RNI7MJUZ0Z_20 ));
    Odrv4 I__15495 (
            .O(N__71412),
            .I(\pid_front.error_i_reg_esr_RNI7MJUZ0Z_20 ));
    InMux I__15494 (
            .O(N__71407),
            .I(N__71401));
    InMux I__15493 (
            .O(N__71406),
            .I(N__71401));
    LocalMux I__15492 (
            .O(N__71401),
            .I(\pid_front.error_i_acumm_preregZ0Z_20 ));
    InMux I__15491 (
            .O(N__71398),
            .I(N__71394));
    InMux I__15490 (
            .O(N__71397),
            .I(N__71391));
    LocalMux I__15489 (
            .O(N__71394),
            .I(N__71387));
    LocalMux I__15488 (
            .O(N__71391),
            .I(N__71384));
    InMux I__15487 (
            .O(N__71390),
            .I(N__71381));
    Span4Mux_v I__15486 (
            .O(N__71387),
            .I(N__71376));
    Span4Mux_v I__15485 (
            .O(N__71384),
            .I(N__71376));
    LocalMux I__15484 (
            .O(N__71381),
            .I(\pid_front.error_i_reg_esr_RNI08DVZ0Z_21 ));
    Odrv4 I__15483 (
            .O(N__71376),
            .I(\pid_front.error_i_reg_esr_RNI08DVZ0Z_21 ));
    InMux I__15482 (
            .O(N__71371),
            .I(N__71365));
    InMux I__15481 (
            .O(N__71370),
            .I(N__71365));
    LocalMux I__15480 (
            .O(N__71365),
            .I(\pid_front.error_i_acumm_preregZ0Z_21 ));
    InMux I__15479 (
            .O(N__71362),
            .I(N__71354));
    InMux I__15478 (
            .O(N__71361),
            .I(N__71354));
    InMux I__15477 (
            .O(N__71360),
            .I(N__71349));
    InMux I__15476 (
            .O(N__71359),
            .I(N__71349));
    LocalMux I__15475 (
            .O(N__71354),
            .I(\pid_front.error_d_reg_prevZ0Z_9 ));
    LocalMux I__15474 (
            .O(N__71349),
            .I(\pid_front.error_d_reg_prevZ0Z_9 ));
    InMux I__15473 (
            .O(N__71344),
            .I(N__71341));
    LocalMux I__15472 (
            .O(N__71341),
            .I(\pid_front.N_2376_i ));
    InMux I__15471 (
            .O(N__71338),
            .I(N__71333));
    InMux I__15470 (
            .O(N__71337),
            .I(N__71328));
    InMux I__15469 (
            .O(N__71336),
            .I(N__71328));
    LocalMux I__15468 (
            .O(N__71333),
            .I(N__71325));
    LocalMux I__15467 (
            .O(N__71328),
            .I(\pid_front.error_d_reg_prevZ0Z_8 ));
    Odrv4 I__15466 (
            .O(N__71325),
            .I(\pid_front.error_d_reg_prevZ0Z_8 ));
    CascadeMux I__15465 (
            .O(N__71320),
            .I(N__71317));
    InMux I__15464 (
            .O(N__71317),
            .I(N__71311));
    InMux I__15463 (
            .O(N__71316),
            .I(N__71311));
    LocalMux I__15462 (
            .O(N__71311),
            .I(N__71308));
    Span4Mux_v I__15461 (
            .O(N__71308),
            .I(N__71305));
    Span4Mux_h I__15460 (
            .O(N__71305),
            .I(N__71302));
    Span4Mux_h I__15459 (
            .O(N__71302),
            .I(N__71299));
    Span4Mux_v I__15458 (
            .O(N__71299),
            .I(N__71296));
    Odrv4 I__15457 (
            .O(N__71296),
            .I(\pid_front.error_p_regZ0Z_9 ));
    CascadeMux I__15456 (
            .O(N__71293),
            .I(\pid_front.N_2376_i_cascade_ ));
    InMux I__15455 (
            .O(N__71290),
            .I(N__71287));
    LocalMux I__15454 (
            .O(N__71287),
            .I(N__71283));
    InMux I__15453 (
            .O(N__71286),
            .I(N__71280));
    Span4Mux_h I__15452 (
            .O(N__71283),
            .I(N__71277));
    LocalMux I__15451 (
            .O(N__71280),
            .I(N__71274));
    Span4Mux_h I__15450 (
            .O(N__71277),
            .I(N__71271));
    Odrv4 I__15449 (
            .O(N__71274),
            .I(\pid_front.error_p_reg_esr_RNILQ6F_0Z0Z_9 ));
    Odrv4 I__15448 (
            .O(N__71271),
            .I(\pid_front.error_p_reg_esr_RNILQ6F_0Z0Z_9 ));
    InMux I__15447 (
            .O(N__71266),
            .I(N__71260));
    InMux I__15446 (
            .O(N__71265),
            .I(N__71260));
    LocalMux I__15445 (
            .O(N__71260),
            .I(\pid_front.error_i_acumm_preregZ0Z_15 ));
    InMux I__15444 (
            .O(N__71257),
            .I(N__71252));
    InMux I__15443 (
            .O(N__71256),
            .I(N__71247));
    InMux I__15442 (
            .O(N__71255),
            .I(N__71247));
    LocalMux I__15441 (
            .O(N__71252),
            .I(N__71244));
    LocalMux I__15440 (
            .O(N__71247),
            .I(N__71241));
    Span4Mux_h I__15439 (
            .O(N__71244),
            .I(N__71236));
    Span4Mux_v I__15438 (
            .O(N__71241),
            .I(N__71236));
    Odrv4 I__15437 (
            .O(N__71236),
            .I(\pid_front.error_i_reg_esr_RNI8IEUZ0Z_16 ));
    InMux I__15436 (
            .O(N__71233),
            .I(N__71227));
    InMux I__15435 (
            .O(N__71232),
            .I(N__71227));
    LocalMux I__15434 (
            .O(N__71227),
            .I(\pid_front.error_i_acumm_preregZ0Z_16 ));
    InMux I__15433 (
            .O(N__71224),
            .I(N__71220));
    InMux I__15432 (
            .O(N__71223),
            .I(N__71216));
    LocalMux I__15431 (
            .O(N__71220),
            .I(N__71213));
    InMux I__15430 (
            .O(N__71219),
            .I(N__71210));
    LocalMux I__15429 (
            .O(N__71216),
            .I(N__71207));
    Span4Mux_h I__15428 (
            .O(N__71213),
            .I(N__71202));
    LocalMux I__15427 (
            .O(N__71210),
            .I(N__71202));
    Span4Mux_v I__15426 (
            .O(N__71207),
            .I(N__71197));
    Span4Mux_v I__15425 (
            .O(N__71202),
            .I(N__71197));
    Odrv4 I__15424 (
            .O(N__71197),
            .I(\pid_front.error_i_reg_esr_RNIALFUZ0Z_17 ));
    InMux I__15423 (
            .O(N__71194),
            .I(N__71188));
    InMux I__15422 (
            .O(N__71193),
            .I(N__71188));
    LocalMux I__15421 (
            .O(N__71188),
            .I(\pid_front.error_i_acumm_preregZ0Z_17 ));
    InMux I__15420 (
            .O(N__71185),
            .I(N__71180));
    InMux I__15419 (
            .O(N__71184),
            .I(N__71175));
    InMux I__15418 (
            .O(N__71183),
            .I(N__71175));
    LocalMux I__15417 (
            .O(N__71180),
            .I(N__71172));
    LocalMux I__15416 (
            .O(N__71175),
            .I(N__71169));
    Span4Mux_v I__15415 (
            .O(N__71172),
            .I(N__71164));
    Span4Mux_v I__15414 (
            .O(N__71169),
            .I(N__71164));
    Odrv4 I__15413 (
            .O(N__71164),
            .I(\pid_front.error_i_reg_esr_RNI6HGVZ0Z_24 ));
    CascadeMux I__15412 (
            .O(N__71161),
            .I(N__71157));
    CascadeMux I__15411 (
            .O(N__71160),
            .I(N__71154));
    InMux I__15410 (
            .O(N__71157),
            .I(N__71149));
    InMux I__15409 (
            .O(N__71154),
            .I(N__71149));
    LocalMux I__15408 (
            .O(N__71149),
            .I(\pid_front.error_i_acumm_preregZ0Z_24 ));
    InMux I__15407 (
            .O(N__71146),
            .I(N__71143));
    LocalMux I__15406 (
            .O(N__71143),
            .I(N__71139));
    InMux I__15405 (
            .O(N__71142),
            .I(N__71136));
    Odrv12 I__15404 (
            .O(N__71139),
            .I(\pid_front.error_p_reg_esr_RNIK3C61_0Z0Z_15 ));
    LocalMux I__15403 (
            .O(N__71136),
            .I(\pid_front.error_p_reg_esr_RNIK3C61_0Z0Z_15 ));
    InMux I__15402 (
            .O(N__71131),
            .I(N__71128));
    LocalMux I__15401 (
            .O(N__71128),
            .I(N__71124));
    InMux I__15400 (
            .O(N__71127),
            .I(N__71121));
    Odrv4 I__15399 (
            .O(N__71124),
            .I(\pid_front.error_p_reg_esr_RNIH0C61Z0Z_14 ));
    LocalMux I__15398 (
            .O(N__71121),
            .I(\pid_front.error_p_reg_esr_RNIH0C61Z0Z_14 ));
    InMux I__15397 (
            .O(N__71116),
            .I(N__71111));
    InMux I__15396 (
            .O(N__71115),
            .I(N__71106));
    InMux I__15395 (
            .O(N__71114),
            .I(N__71106));
    LocalMux I__15394 (
            .O(N__71111),
            .I(N__71103));
    LocalMux I__15393 (
            .O(N__71106),
            .I(N__71100));
    Span4Mux_v I__15392 (
            .O(N__71103),
            .I(N__71095));
    Span4Mux_h I__15391 (
            .O(N__71100),
            .I(N__71095));
    Odrv4 I__15390 (
            .O(N__71095),
            .I(\pid_front.error_i_reg_esr_RNI6FDUZ0Z_15 ));
    InMux I__15389 (
            .O(N__71092),
            .I(N__71088));
    InMux I__15388 (
            .O(N__71091),
            .I(N__71085));
    LocalMux I__15387 (
            .O(N__71088),
            .I(N__71082));
    LocalMux I__15386 (
            .O(N__71085),
            .I(N__71079));
    Span4Mux_v I__15385 (
            .O(N__71082),
            .I(N__71076));
    Span12Mux_v I__15384 (
            .O(N__71079),
            .I(N__71073));
    Odrv4 I__15383 (
            .O(N__71076),
            .I(\pid_front.error_p_reg_esr_RNIBJ5B3_0Z0Z_14 ));
    Odrv12 I__15382 (
            .O(N__71073),
            .I(\pid_front.error_p_reg_esr_RNIBJ5B3_0Z0Z_14 ));
    CascadeMux I__15381 (
            .O(N__71068),
            .I(N__71065));
    InMux I__15380 (
            .O(N__71065),
            .I(N__71058));
    InMux I__15379 (
            .O(N__71064),
            .I(N__71052));
    InMux I__15378 (
            .O(N__71063),
            .I(N__71052));
    CascadeMux I__15377 (
            .O(N__71062),
            .I(N__71048));
    CascadeMux I__15376 (
            .O(N__71061),
            .I(N__71041));
    LocalMux I__15375 (
            .O(N__71058),
            .I(N__71034));
    InMux I__15374 (
            .O(N__71057),
            .I(N__71031));
    LocalMux I__15373 (
            .O(N__71052),
            .I(N__71019));
    InMux I__15372 (
            .O(N__71051),
            .I(N__71008));
    InMux I__15371 (
            .O(N__71048),
            .I(N__71008));
    InMux I__15370 (
            .O(N__71047),
            .I(N__71008));
    InMux I__15369 (
            .O(N__71046),
            .I(N__71008));
    IoInMux I__15368 (
            .O(N__71045),
            .I(N__71005));
    InMux I__15367 (
            .O(N__71044),
            .I(N__70998));
    InMux I__15366 (
            .O(N__71041),
            .I(N__70998));
    InMux I__15365 (
            .O(N__71040),
            .I(N__70998));
    InMux I__15364 (
            .O(N__71039),
            .I(N__70993));
    InMux I__15363 (
            .O(N__71038),
            .I(N__70993));
    InMux I__15362 (
            .O(N__71037),
            .I(N__70990));
    Span4Mux_h I__15361 (
            .O(N__71034),
            .I(N__70985));
    LocalMux I__15360 (
            .O(N__71031),
            .I(N__70985));
    InMux I__15359 (
            .O(N__71030),
            .I(N__70974));
    InMux I__15358 (
            .O(N__71029),
            .I(N__70967));
    InMux I__15357 (
            .O(N__71028),
            .I(N__70967));
    InMux I__15356 (
            .O(N__71027),
            .I(N__70955));
    InMux I__15355 (
            .O(N__71026),
            .I(N__70955));
    InMux I__15354 (
            .O(N__71025),
            .I(N__70948));
    InMux I__15353 (
            .O(N__71024),
            .I(N__70948));
    InMux I__15352 (
            .O(N__71023),
            .I(N__70948));
    InMux I__15351 (
            .O(N__71022),
            .I(N__70945));
    Span4Mux_v I__15350 (
            .O(N__71019),
            .I(N__70942));
    InMux I__15349 (
            .O(N__71018),
            .I(N__70939));
    InMux I__15348 (
            .O(N__71017),
            .I(N__70935));
    LocalMux I__15347 (
            .O(N__71008),
            .I(N__70930));
    LocalMux I__15346 (
            .O(N__71005),
            .I(N__70930));
    LocalMux I__15345 (
            .O(N__70998),
            .I(N__70926));
    LocalMux I__15344 (
            .O(N__70993),
            .I(N__70919));
    LocalMux I__15343 (
            .O(N__70990),
            .I(N__70919));
    Span4Mux_h I__15342 (
            .O(N__70985),
            .I(N__70919));
    InMux I__15341 (
            .O(N__70984),
            .I(N__70911));
    InMux I__15340 (
            .O(N__70983),
            .I(N__70911));
    InMux I__15339 (
            .O(N__70982),
            .I(N__70911));
    InMux I__15338 (
            .O(N__70981),
            .I(N__70906));
    InMux I__15337 (
            .O(N__70980),
            .I(N__70906));
    InMux I__15336 (
            .O(N__70979),
            .I(N__70899));
    InMux I__15335 (
            .O(N__70978),
            .I(N__70899));
    InMux I__15334 (
            .O(N__70977),
            .I(N__70899));
    LocalMux I__15333 (
            .O(N__70974),
            .I(N__70896));
    InMux I__15332 (
            .O(N__70973),
            .I(N__70893));
    InMux I__15331 (
            .O(N__70972),
            .I(N__70890));
    LocalMux I__15330 (
            .O(N__70967),
            .I(N__70887));
    InMux I__15329 (
            .O(N__70966),
            .I(N__70884));
    InMux I__15328 (
            .O(N__70965),
            .I(N__70881));
    InMux I__15327 (
            .O(N__70964),
            .I(N__70875));
    InMux I__15326 (
            .O(N__70963),
            .I(N__70875));
    InMux I__15325 (
            .O(N__70962),
            .I(N__70870));
    InMux I__15324 (
            .O(N__70961),
            .I(N__70870));
    InMux I__15323 (
            .O(N__70960),
            .I(N__70867));
    LocalMux I__15322 (
            .O(N__70955),
            .I(N__70864));
    LocalMux I__15321 (
            .O(N__70948),
            .I(N__70861));
    LocalMux I__15320 (
            .O(N__70945),
            .I(N__70858));
    Span4Mux_v I__15319 (
            .O(N__70942),
            .I(N__70855));
    LocalMux I__15318 (
            .O(N__70939),
            .I(N__70852));
    InMux I__15317 (
            .O(N__70938),
            .I(N__70847));
    LocalMux I__15316 (
            .O(N__70935),
            .I(N__70844));
    Span4Mux_s3_v I__15315 (
            .O(N__70930),
            .I(N__70840));
    InMux I__15314 (
            .O(N__70929),
            .I(N__70835));
    Span4Mux_h I__15313 (
            .O(N__70926),
            .I(N__70830));
    Span4Mux_v I__15312 (
            .O(N__70919),
            .I(N__70830));
    InMux I__15311 (
            .O(N__70918),
            .I(N__70827));
    LocalMux I__15310 (
            .O(N__70911),
            .I(N__70820));
    LocalMux I__15309 (
            .O(N__70906),
            .I(N__70820));
    LocalMux I__15308 (
            .O(N__70899),
            .I(N__70820));
    Span4Mux_h I__15307 (
            .O(N__70896),
            .I(N__70817));
    LocalMux I__15306 (
            .O(N__70893),
            .I(N__70812));
    LocalMux I__15305 (
            .O(N__70890),
            .I(N__70812));
    Span4Mux_v I__15304 (
            .O(N__70887),
            .I(N__70807));
    LocalMux I__15303 (
            .O(N__70884),
            .I(N__70797));
    LocalMux I__15302 (
            .O(N__70881),
            .I(N__70797));
    InMux I__15301 (
            .O(N__70880),
            .I(N__70791));
    LocalMux I__15300 (
            .O(N__70875),
            .I(N__70788));
    LocalMux I__15299 (
            .O(N__70870),
            .I(N__70781));
    LocalMux I__15298 (
            .O(N__70867),
            .I(N__70781));
    Span4Mux_v I__15297 (
            .O(N__70864),
            .I(N__70781));
    Span4Mux_h I__15296 (
            .O(N__70861),
            .I(N__70776));
    Span4Mux_v I__15295 (
            .O(N__70858),
            .I(N__70776));
    Span4Mux_h I__15294 (
            .O(N__70855),
            .I(N__70771));
    Span4Mux_v I__15293 (
            .O(N__70852),
            .I(N__70771));
    InMux I__15292 (
            .O(N__70851),
            .I(N__70766));
    InMux I__15291 (
            .O(N__70850),
            .I(N__70766));
    LocalMux I__15290 (
            .O(N__70847),
            .I(N__70763));
    Span4Mux_v I__15289 (
            .O(N__70844),
            .I(N__70760));
    InMux I__15288 (
            .O(N__70843),
            .I(N__70757));
    Span4Mux_v I__15287 (
            .O(N__70840),
            .I(N__70754));
    InMux I__15286 (
            .O(N__70839),
            .I(N__70750));
    InMux I__15285 (
            .O(N__70838),
            .I(N__70747));
    LocalMux I__15284 (
            .O(N__70835),
            .I(N__70740));
    Span4Mux_v I__15283 (
            .O(N__70830),
            .I(N__70740));
    LocalMux I__15282 (
            .O(N__70827),
            .I(N__70740));
    Span4Mux_v I__15281 (
            .O(N__70820),
            .I(N__70737));
    Span4Mux_h I__15280 (
            .O(N__70817),
            .I(N__70732));
    Span4Mux_v I__15279 (
            .O(N__70812),
            .I(N__70732));
    InMux I__15278 (
            .O(N__70811),
            .I(N__70724));
    InMux I__15277 (
            .O(N__70810),
            .I(N__70724));
    Span4Mux_h I__15276 (
            .O(N__70807),
            .I(N__70721));
    InMux I__15275 (
            .O(N__70806),
            .I(N__70716));
    InMux I__15274 (
            .O(N__70805),
            .I(N__70716));
    InMux I__15273 (
            .O(N__70804),
            .I(N__70709));
    InMux I__15272 (
            .O(N__70803),
            .I(N__70709));
    InMux I__15271 (
            .O(N__70802),
            .I(N__70709));
    Span4Mux_h I__15270 (
            .O(N__70797),
            .I(N__70706));
    InMux I__15269 (
            .O(N__70796),
            .I(N__70697));
    InMux I__15268 (
            .O(N__70795),
            .I(N__70697));
    InMux I__15267 (
            .O(N__70794),
            .I(N__70697));
    LocalMux I__15266 (
            .O(N__70791),
            .I(N__70688));
    Span4Mux_v I__15265 (
            .O(N__70788),
            .I(N__70688));
    Span4Mux_h I__15264 (
            .O(N__70781),
            .I(N__70688));
    Span4Mux_v I__15263 (
            .O(N__70776),
            .I(N__70688));
    Span4Mux_v I__15262 (
            .O(N__70771),
            .I(N__70683));
    LocalMux I__15261 (
            .O(N__70766),
            .I(N__70683));
    Span4Mux_v I__15260 (
            .O(N__70763),
            .I(N__70674));
    Span4Mux_v I__15259 (
            .O(N__70760),
            .I(N__70674));
    LocalMux I__15258 (
            .O(N__70757),
            .I(N__70674));
    Span4Mux_v I__15257 (
            .O(N__70754),
            .I(N__70674));
    InMux I__15256 (
            .O(N__70753),
            .I(N__70671));
    LocalMux I__15255 (
            .O(N__70750),
            .I(N__70666));
    LocalMux I__15254 (
            .O(N__70747),
            .I(N__70666));
    Span4Mux_h I__15253 (
            .O(N__70740),
            .I(N__70659));
    Span4Mux_h I__15252 (
            .O(N__70737),
            .I(N__70659));
    Span4Mux_v I__15251 (
            .O(N__70732),
            .I(N__70659));
    InMux I__15250 (
            .O(N__70731),
            .I(N__70652));
    InMux I__15249 (
            .O(N__70730),
            .I(N__70652));
    InMux I__15248 (
            .O(N__70729),
            .I(N__70652));
    LocalMux I__15247 (
            .O(N__70724),
            .I(N__70641));
    Span4Mux_h I__15246 (
            .O(N__70721),
            .I(N__70641));
    LocalMux I__15245 (
            .O(N__70716),
            .I(N__70641));
    LocalMux I__15244 (
            .O(N__70709),
            .I(N__70641));
    Span4Mux_v I__15243 (
            .O(N__70706),
            .I(N__70641));
    InMux I__15242 (
            .O(N__70705),
            .I(N__70636));
    InMux I__15241 (
            .O(N__70704),
            .I(N__70636));
    LocalMux I__15240 (
            .O(N__70697),
            .I(N__70627));
    Span4Mux_v I__15239 (
            .O(N__70688),
            .I(N__70627));
    Span4Mux_v I__15238 (
            .O(N__70683),
            .I(N__70627));
    Span4Mux_h I__15237 (
            .O(N__70674),
            .I(N__70627));
    LocalMux I__15236 (
            .O(N__70671),
            .I(reset_system));
    Odrv12 I__15235 (
            .O(N__70666),
            .I(reset_system));
    Odrv4 I__15234 (
            .O(N__70659),
            .I(reset_system));
    LocalMux I__15233 (
            .O(N__70652),
            .I(reset_system));
    Odrv4 I__15232 (
            .O(N__70641),
            .I(reset_system));
    LocalMux I__15231 (
            .O(N__70636),
            .I(reset_system));
    Odrv4 I__15230 (
            .O(N__70627),
            .I(reset_system));
    CascadeMux I__15229 (
            .O(N__70612),
            .I(N__70607));
    CascadeMux I__15228 (
            .O(N__70611),
            .I(N__70601));
    InMux I__15227 (
            .O(N__70610),
            .I(N__70596));
    InMux I__15226 (
            .O(N__70607),
            .I(N__70596));
    InMux I__15225 (
            .O(N__70606),
            .I(N__70593));
    InMux I__15224 (
            .O(N__70605),
            .I(N__70590));
    InMux I__15223 (
            .O(N__70604),
            .I(N__70587));
    InMux I__15222 (
            .O(N__70601),
            .I(N__70584));
    LocalMux I__15221 (
            .O(N__70596),
            .I(N__70581));
    LocalMux I__15220 (
            .O(N__70593),
            .I(N__70578));
    LocalMux I__15219 (
            .O(N__70590),
            .I(N__70575));
    LocalMux I__15218 (
            .O(N__70587),
            .I(N__70572));
    LocalMux I__15217 (
            .O(N__70584),
            .I(N__70569));
    Span4Mux_h I__15216 (
            .O(N__70581),
            .I(N__70566));
    Span4Mux_h I__15215 (
            .O(N__70578),
            .I(N__70563));
    Span4Mux_v I__15214 (
            .O(N__70575),
            .I(N__70560));
    Sp12to4 I__15213 (
            .O(N__70572),
            .I(N__70554));
    Span4Mux_v I__15212 (
            .O(N__70569),
            .I(N__70551));
    Span4Mux_h I__15211 (
            .O(N__70566),
            .I(N__70544));
    Span4Mux_h I__15210 (
            .O(N__70563),
            .I(N__70544));
    Span4Mux_v I__15209 (
            .O(N__70560),
            .I(N__70544));
    InMux I__15208 (
            .O(N__70559),
            .I(N__70537));
    InMux I__15207 (
            .O(N__70558),
            .I(N__70537));
    InMux I__15206 (
            .O(N__70557),
            .I(N__70537));
    Span12Mux_v I__15205 (
            .O(N__70554),
            .I(N__70534));
    Odrv4 I__15204 (
            .O(N__70551),
            .I(\pid_front.stateZ0Z_0 ));
    Odrv4 I__15203 (
            .O(N__70544),
            .I(\pid_front.stateZ0Z_0 ));
    LocalMux I__15202 (
            .O(N__70537),
            .I(\pid_front.stateZ0Z_0 ));
    Odrv12 I__15201 (
            .O(N__70534),
            .I(\pid_front.stateZ0Z_0 ));
    CascadeMux I__15200 (
            .O(N__70525),
            .I(\pid_front.N_382_cascade_ ));
    InMux I__15199 (
            .O(N__70522),
            .I(N__70502));
    InMux I__15198 (
            .O(N__70521),
            .I(N__70502));
    InMux I__15197 (
            .O(N__70520),
            .I(N__70502));
    InMux I__15196 (
            .O(N__70519),
            .I(N__70502));
    InMux I__15195 (
            .O(N__70518),
            .I(N__70502));
    InMux I__15194 (
            .O(N__70517),
            .I(N__70502));
    CascadeMux I__15193 (
            .O(N__70516),
            .I(N__70499));
    InMux I__15192 (
            .O(N__70515),
            .I(N__70492));
    LocalMux I__15191 (
            .O(N__70502),
            .I(N__70489));
    InMux I__15190 (
            .O(N__70499),
            .I(N__70486));
    InMux I__15189 (
            .O(N__70498),
            .I(N__70483));
    InMux I__15188 (
            .O(N__70497),
            .I(N__70479));
    InMux I__15187 (
            .O(N__70496),
            .I(N__70476));
    InMux I__15186 (
            .O(N__70495),
            .I(N__70473));
    LocalMux I__15185 (
            .O(N__70492),
            .I(N__70470));
    Span4Mux_v I__15184 (
            .O(N__70489),
            .I(N__70462));
    LocalMux I__15183 (
            .O(N__70486),
            .I(N__70462));
    LocalMux I__15182 (
            .O(N__70483),
            .I(N__70462));
    CascadeMux I__15181 (
            .O(N__70482),
            .I(N__70458));
    LocalMux I__15180 (
            .O(N__70479),
            .I(N__70451));
    LocalMux I__15179 (
            .O(N__70476),
            .I(N__70451));
    LocalMux I__15178 (
            .O(N__70473),
            .I(N__70451));
    Span4Mux_h I__15177 (
            .O(N__70470),
            .I(N__70448));
    CascadeMux I__15176 (
            .O(N__70469),
            .I(N__70444));
    Span4Mux_v I__15175 (
            .O(N__70462),
            .I(N__70441));
    InMux I__15174 (
            .O(N__70461),
            .I(N__70436));
    InMux I__15173 (
            .O(N__70458),
            .I(N__70436));
    Span4Mux_v I__15172 (
            .O(N__70451),
            .I(N__70433));
    Span4Mux_v I__15171 (
            .O(N__70448),
            .I(N__70430));
    InMux I__15170 (
            .O(N__70447),
            .I(N__70425));
    InMux I__15169 (
            .O(N__70444),
            .I(N__70425));
    Span4Mux_v I__15168 (
            .O(N__70441),
            .I(N__70422));
    LocalMux I__15167 (
            .O(N__70436),
            .I(\pid_front.stateZ0Z_1 ));
    Odrv4 I__15166 (
            .O(N__70433),
            .I(\pid_front.stateZ0Z_1 ));
    Odrv4 I__15165 (
            .O(N__70430),
            .I(\pid_front.stateZ0Z_1 ));
    LocalMux I__15164 (
            .O(N__70425),
            .I(\pid_front.stateZ0Z_1 ));
    Odrv4 I__15163 (
            .O(N__70422),
            .I(\pid_front.stateZ0Z_1 ));
    InMux I__15162 (
            .O(N__70411),
            .I(N__70407));
    InMux I__15161 (
            .O(N__70410),
            .I(N__70404));
    LocalMux I__15160 (
            .O(N__70407),
            .I(\pid_front.N_217 ));
    LocalMux I__15159 (
            .O(N__70404),
            .I(\pid_front.N_217 ));
    InMux I__15158 (
            .O(N__70399),
            .I(N__70396));
    LocalMux I__15157 (
            .O(N__70396),
            .I(N__70391));
    InMux I__15156 (
            .O(N__70395),
            .I(N__70386));
    InMux I__15155 (
            .O(N__70394),
            .I(N__70386));
    Span4Mux_v I__15154 (
            .O(N__70391),
            .I(N__70383));
    LocalMux I__15153 (
            .O(N__70386),
            .I(N__70380));
    Odrv4 I__15152 (
            .O(N__70383),
            .I(\pid_front.error_p_regZ0Z_10 ));
    Odrv4 I__15151 (
            .O(N__70380),
            .I(\pid_front.error_p_regZ0Z_10 ));
    CascadeMux I__15150 (
            .O(N__70375),
            .I(\pid_front.N_2382_i_cascade_ ));
    CascadeMux I__15149 (
            .O(N__70372),
            .I(\pid_front.error_p_reg_esr_RNIFM3D1Z0Z_10_cascade_ ));
    CascadeMux I__15148 (
            .O(N__70369),
            .I(N__70366));
    InMux I__15147 (
            .O(N__70366),
            .I(N__70362));
    InMux I__15146 (
            .O(N__70365),
            .I(N__70359));
    LocalMux I__15145 (
            .O(N__70362),
            .I(N__70356));
    LocalMux I__15144 (
            .O(N__70359),
            .I(N__70353));
    Span4Mux_h I__15143 (
            .O(N__70356),
            .I(N__70350));
    Odrv4 I__15142 (
            .O(N__70353),
            .I(\pid_front.error_p_reg_esr_RNI6R6D1Z0Z_8 ));
    Odrv4 I__15141 (
            .O(N__70350),
            .I(\pid_front.error_p_reg_esr_RNI6R6D1Z0Z_8 ));
    InMux I__15140 (
            .O(N__70345),
            .I(N__70342));
    LocalMux I__15139 (
            .O(N__70342),
            .I(N__70339));
    Span4Mux_v I__15138 (
            .O(N__70339),
            .I(N__70336));
    Odrv4 I__15137 (
            .O(N__70336),
            .I(\pid_front.error_p_reg_esr_RNIS5CU3Z0Z_9 ));
    InMux I__15136 (
            .O(N__70333),
            .I(N__70327));
    InMux I__15135 (
            .O(N__70332),
            .I(N__70327));
    LocalMux I__15134 (
            .O(N__70327),
            .I(\pid_front.error_p_reg_esr_RNILQ6FZ0Z_9 ));
    CascadeMux I__15133 (
            .O(N__70324),
            .I(N__70321));
    InMux I__15132 (
            .O(N__70321),
            .I(N__70318));
    LocalMux I__15131 (
            .O(N__70318),
            .I(N__70315));
    Span4Mux_v I__15130 (
            .O(N__70315),
            .I(N__70311));
    InMux I__15129 (
            .O(N__70314),
            .I(N__70308));
    Odrv4 I__15128 (
            .O(N__70311),
            .I(\pid_front.error_d_reg_prev_esr_RNI1K4E5_0Z0Z_10 ));
    LocalMux I__15127 (
            .O(N__70308),
            .I(\pid_front.error_d_reg_prev_esr_RNI1K4E5_0Z0Z_10 ));
    InMux I__15126 (
            .O(N__70303),
            .I(N__70300));
    LocalMux I__15125 (
            .O(N__70300),
            .I(\pid_front.error_p_reg_esr_RNIFM3D1Z0Z_10 ));
    CascadeMux I__15124 (
            .O(N__70297),
            .I(N__70294));
    InMux I__15123 (
            .O(N__70294),
            .I(N__70291));
    LocalMux I__15122 (
            .O(N__70291),
            .I(N__70288));
    Span4Mux_h I__15121 (
            .O(N__70288),
            .I(N__70285));
    Odrv4 I__15120 (
            .O(N__70285),
            .I(\pid_front.error_p_reg_esr_RNINU9V7Z0Z_9 ));
    CascadeMux I__15119 (
            .O(N__70282),
            .I(N__70278));
    InMux I__15118 (
            .O(N__70281),
            .I(N__70274));
    InMux I__15117 (
            .O(N__70278),
            .I(N__70269));
    InMux I__15116 (
            .O(N__70277),
            .I(N__70269));
    LocalMux I__15115 (
            .O(N__70274),
            .I(N__70263));
    LocalMux I__15114 (
            .O(N__70269),
            .I(N__70263));
    InMux I__15113 (
            .O(N__70268),
            .I(N__70260));
    Span4Mux_h I__15112 (
            .O(N__70263),
            .I(N__70257));
    LocalMux I__15111 (
            .O(N__70260),
            .I(\pid_front.error_d_reg_prevZ0Z_10 ));
    Odrv4 I__15110 (
            .O(N__70257),
            .I(\pid_front.error_d_reg_prevZ0Z_10 ));
    InMux I__15109 (
            .O(N__70252),
            .I(N__70249));
    LocalMux I__15108 (
            .O(N__70249),
            .I(N__70246));
    Span4Mux_h I__15107 (
            .O(N__70246),
            .I(N__70243));
    Odrv4 I__15106 (
            .O(N__70243),
            .I(\pid_side.N_109 ));
    CascadeMux I__15105 (
            .O(N__70240),
            .I(N__70237));
    InMux I__15104 (
            .O(N__70237),
            .I(N__70231));
    InMux I__15103 (
            .O(N__70236),
            .I(N__70231));
    LocalMux I__15102 (
            .O(N__70231),
            .I(N__70228));
    Odrv4 I__15101 (
            .O(N__70228),
            .I(\pid_front.error_d_reg_prevZ0Z_19 ));
    InMux I__15100 (
            .O(N__70225),
            .I(N__70219));
    InMux I__15099 (
            .O(N__70224),
            .I(N__70219));
    LocalMux I__15098 (
            .O(N__70219),
            .I(N__70216));
    Sp12to4 I__15097 (
            .O(N__70216),
            .I(N__70213));
    Span12Mux_v I__15096 (
            .O(N__70213),
            .I(N__70210));
    Span12Mux_h I__15095 (
            .O(N__70210),
            .I(N__70207));
    Odrv12 I__15094 (
            .O(N__70207),
            .I(\pid_front.error_p_regZ0Z_19 ));
    InMux I__15093 (
            .O(N__70204),
            .I(N__70198));
    InMux I__15092 (
            .O(N__70203),
            .I(N__70198));
    LocalMux I__15091 (
            .O(N__70198),
            .I(N__70195));
    Span4Mux_v I__15090 (
            .O(N__70195),
            .I(N__70192));
    Span4Mux_h I__15089 (
            .O(N__70192),
            .I(N__70189));
    Odrv4 I__15088 (
            .O(N__70189),
            .I(\pid_front.error_p_reg_esr_RNI0GC61Z0Z_19 ));
    CascadeMux I__15087 (
            .O(N__70186),
            .I(\pid_front.N_531_cascade_ ));
    InMux I__15086 (
            .O(N__70183),
            .I(N__70177));
    InMux I__15085 (
            .O(N__70182),
            .I(N__70177));
    LocalMux I__15084 (
            .O(N__70177),
            .I(\pid_front.N_255 ));
    InMux I__15083 (
            .O(N__70174),
            .I(N__70171));
    LocalMux I__15082 (
            .O(N__70171),
            .I(N__70166));
    InMux I__15081 (
            .O(N__70170),
            .I(N__70161));
    InMux I__15080 (
            .O(N__70169),
            .I(N__70161));
    Span4Mux_h I__15079 (
            .O(N__70166),
            .I(N__70158));
    LocalMux I__15078 (
            .O(N__70161),
            .I(N__70155));
    Odrv4 I__15077 (
            .O(N__70158),
            .I(\pid_front.error_i_acumm_preregZ0Z_9 ));
    Odrv4 I__15076 (
            .O(N__70155),
            .I(\pid_front.error_i_acumm_preregZ0Z_9 ));
    CascadeMux I__15075 (
            .O(N__70150),
            .I(N__70146));
    InMux I__15074 (
            .O(N__70149),
            .I(N__70140));
    InMux I__15073 (
            .O(N__70146),
            .I(N__70140));
    InMux I__15072 (
            .O(N__70145),
            .I(N__70137));
    LocalMux I__15071 (
            .O(N__70140),
            .I(\pid_front.N_633 ));
    LocalMux I__15070 (
            .O(N__70137),
            .I(\pid_front.N_633 ));
    CascadeMux I__15069 (
            .O(N__70132),
            .I(\pid_front.N_255_cascade_ ));
    InMux I__15068 (
            .O(N__70129),
            .I(N__70126));
    LocalMux I__15067 (
            .O(N__70126),
            .I(N__70123));
    Span4Mux_h I__15066 (
            .O(N__70123),
            .I(N__70120));
    Odrv4 I__15065 (
            .O(N__70120),
            .I(\pid_front.error_i_acummZ0Z_9 ));
    InMux I__15064 (
            .O(N__70117),
            .I(N__70113));
    InMux I__15063 (
            .O(N__70116),
            .I(N__70110));
    LocalMux I__15062 (
            .O(N__70113),
            .I(N__70107));
    LocalMux I__15061 (
            .O(N__70110),
            .I(N__70104));
    Odrv12 I__15060 (
            .O(N__70107),
            .I(\pid_front.N_276 ));
    Odrv4 I__15059 (
            .O(N__70104),
            .I(\pid_front.N_276 ));
    CascadeMux I__15058 (
            .O(N__70099),
            .I(\pid_front.N_276_cascade_ ));
    CascadeMux I__15057 (
            .O(N__70096),
            .I(N__70092));
    InMux I__15056 (
            .O(N__70095),
            .I(N__70084));
    InMux I__15055 (
            .O(N__70092),
            .I(N__70084));
    InMux I__15054 (
            .O(N__70091),
            .I(N__70084));
    LocalMux I__15053 (
            .O(N__70084),
            .I(N__70081));
    Odrv4 I__15052 (
            .O(N__70081),
            .I(\pid_front.N_632 ));
    InMux I__15051 (
            .O(N__70078),
            .I(N__70075));
    LocalMux I__15050 (
            .O(N__70075),
            .I(N__70072));
    Span12Mux_s11_h I__15049 (
            .O(N__70072),
            .I(N__70069));
    Odrv12 I__15048 (
            .O(N__70069),
            .I(pid_side_N_382_4));
    InMux I__15047 (
            .O(N__70066),
            .I(N__70062));
    InMux I__15046 (
            .O(N__70065),
            .I(N__70058));
    LocalMux I__15045 (
            .O(N__70062),
            .I(N__70054));
    InMux I__15044 (
            .O(N__70061),
            .I(N__70051));
    LocalMux I__15043 (
            .O(N__70058),
            .I(N__70048));
    CascadeMux I__15042 (
            .O(N__70057),
            .I(N__70045));
    Span4Mux_v I__15041 (
            .O(N__70054),
            .I(N__70042));
    LocalMux I__15040 (
            .O(N__70051),
            .I(N__70037));
    Sp12to4 I__15039 (
            .O(N__70048),
            .I(N__70037));
    InMux I__15038 (
            .O(N__70045),
            .I(N__70034));
    Odrv4 I__15037 (
            .O(N__70042),
            .I(xy_ki_7));
    Odrv12 I__15036 (
            .O(N__70037),
            .I(xy_ki_7));
    LocalMux I__15035 (
            .O(N__70034),
            .I(xy_ki_7));
    InMux I__15034 (
            .O(N__70027),
            .I(N__70024));
    LocalMux I__15033 (
            .O(N__70024),
            .I(N__70019));
    InMux I__15032 (
            .O(N__70023),
            .I(N__70016));
    InMux I__15031 (
            .O(N__70022),
            .I(N__70013));
    Span4Mux_v I__15030 (
            .O(N__70019),
            .I(N__70008));
    LocalMux I__15029 (
            .O(N__70016),
            .I(N__70008));
    LocalMux I__15028 (
            .O(N__70013),
            .I(N__70005));
    Span4Mux_v I__15027 (
            .O(N__70008),
            .I(N__70002));
    Span4Mux_v I__15026 (
            .O(N__70005),
            .I(N__69998));
    Span4Mux_v I__15025 (
            .O(N__70002),
            .I(N__69995));
    InMux I__15024 (
            .O(N__70001),
            .I(N__69992));
    Odrv4 I__15023 (
            .O(N__69998),
            .I(xy_ki_6));
    Odrv4 I__15022 (
            .O(N__69995),
            .I(xy_ki_6));
    LocalMux I__15021 (
            .O(N__69992),
            .I(xy_ki_6));
    CascadeMux I__15020 (
            .O(N__69985),
            .I(\pid_front.N_446_cascade_ ));
    InMux I__15019 (
            .O(N__69982),
            .I(N__69979));
    LocalMux I__15018 (
            .O(N__69979),
            .I(\pid_front.m20_2_03_0_2 ));
    InMux I__15017 (
            .O(N__69976),
            .I(N__69967));
    InMux I__15016 (
            .O(N__69975),
            .I(N__69967));
    InMux I__15015 (
            .O(N__69974),
            .I(N__69967));
    LocalMux I__15014 (
            .O(N__69967),
            .I(\pid_front.N_515 ));
    CascadeMux I__15013 (
            .O(N__69964),
            .I(\pid_front.N_438_cascade_ ));
    InMux I__15012 (
            .O(N__69961),
            .I(N__69958));
    LocalMux I__15011 (
            .O(N__69958),
            .I(N__69954));
    InMux I__15010 (
            .O(N__69957),
            .I(N__69951));
    Span4Mux_h I__15009 (
            .O(N__69954),
            .I(N__69945));
    LocalMux I__15008 (
            .O(N__69951),
            .I(N__69945));
    InMux I__15007 (
            .O(N__69950),
            .I(N__69942));
    Span4Mux_v I__15006 (
            .O(N__69945),
            .I(N__69939));
    LocalMux I__15005 (
            .O(N__69942),
            .I(N__69934));
    Span4Mux_v I__15004 (
            .O(N__69939),
            .I(N__69934));
    Odrv4 I__15003 (
            .O(N__69934),
            .I(\pid_front.error_i_reg_esr_RNI4CCUZ0Z_14 ));
    CascadeMux I__15002 (
            .O(N__69931),
            .I(N__69927));
    InMux I__15001 (
            .O(N__69930),
            .I(N__69924));
    InMux I__15000 (
            .O(N__69927),
            .I(N__69921));
    LocalMux I__14999 (
            .O(N__69924),
            .I(\pid_front.error_i_acumm_preregZ0Z_14 ));
    LocalMux I__14998 (
            .O(N__69921),
            .I(\pid_front.error_i_acumm_preregZ0Z_14 ));
    InMux I__14997 (
            .O(N__69916),
            .I(N__69913));
    LocalMux I__14996 (
            .O(N__69913),
            .I(N__69910));
    Span4Mux_h I__14995 (
            .O(N__69910),
            .I(N__69905));
    InMux I__14994 (
            .O(N__69909),
            .I(N__69900));
    InMux I__14993 (
            .O(N__69908),
            .I(N__69900));
    Odrv4 I__14992 (
            .O(N__69905),
            .I(\pid_front.error_i_reg_esr_RNI2BEVZ0Z_22 ));
    LocalMux I__14991 (
            .O(N__69900),
            .I(\pid_front.error_i_reg_esr_RNI2BEVZ0Z_22 ));
    InMux I__14990 (
            .O(N__69895),
            .I(N__69891));
    InMux I__14989 (
            .O(N__69894),
            .I(N__69888));
    LocalMux I__14988 (
            .O(N__69891),
            .I(\pid_front.error_i_acumm_preregZ0Z_22 ));
    LocalMux I__14987 (
            .O(N__69888),
            .I(\pid_front.error_i_acumm_preregZ0Z_22 ));
    CascadeMux I__14986 (
            .O(N__69883),
            .I(N__69879));
    InMux I__14985 (
            .O(N__69882),
            .I(N__69876));
    InMux I__14984 (
            .O(N__69879),
            .I(N__69873));
    LocalMux I__14983 (
            .O(N__69876),
            .I(N__69870));
    LocalMux I__14982 (
            .O(N__69873),
            .I(N__69867));
    Span4Mux_v I__14981 (
            .O(N__69870),
            .I(N__69863));
    Span4Mux_v I__14980 (
            .O(N__69867),
            .I(N__69860));
    InMux I__14979 (
            .O(N__69866),
            .I(N__69857));
    Odrv4 I__14978 (
            .O(N__69863),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_26_c_RNICQJV ));
    Odrv4 I__14977 (
            .O(N__69860),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_26_c_RNICQJV ));
    LocalMux I__14976 (
            .O(N__69857),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_26_c_RNICQJV ));
    InMux I__14975 (
            .O(N__69850),
            .I(N__69846));
    InMux I__14974 (
            .O(N__69849),
            .I(N__69843));
    LocalMux I__14973 (
            .O(N__69846),
            .I(\pid_front.error_i_acumm_preregZ0Z_27 ));
    LocalMux I__14972 (
            .O(N__69843),
            .I(\pid_front.error_i_acumm_preregZ0Z_27 ));
    InMux I__14971 (
            .O(N__69838),
            .I(N__69835));
    LocalMux I__14970 (
            .O(N__69835),
            .I(\pid_front.N_439 ));
    CascadeMux I__14969 (
            .O(N__69832),
            .I(\pid_front.error_i_reg_esr_RNO_5Z0Z_16_cascade_ ));
    CascadeMux I__14968 (
            .O(N__69829),
            .I(\pid_front.error_i_reg_9_rn_0_16_cascade_ ));
    CascadeMux I__14967 (
            .O(N__69826),
            .I(N__69823));
    InMux I__14966 (
            .O(N__69823),
            .I(N__69820));
    LocalMux I__14965 (
            .O(N__69820),
            .I(N__69817));
    Span4Mux_h I__14964 (
            .O(N__69817),
            .I(N__69814));
    Odrv4 I__14963 (
            .O(N__69814),
            .I(\pid_front.error_i_regZ0Z_16 ));
    InMux I__14962 (
            .O(N__69811),
            .I(N__69808));
    LocalMux I__14961 (
            .O(N__69808),
            .I(\pid_front.error_i_reg_9_sn_16 ));
    InMux I__14960 (
            .O(N__69805),
            .I(N__69802));
    LocalMux I__14959 (
            .O(N__69802),
            .I(N__69799));
    Span4Mux_h I__14958 (
            .O(N__69799),
            .I(N__69796));
    Odrv4 I__14957 (
            .O(N__69796),
            .I(\pid_front.N_188 ));
    InMux I__14956 (
            .O(N__69793),
            .I(N__69790));
    LocalMux I__14955 (
            .O(N__69790),
            .I(\pid_front.N_259 ));
    CascadeMux I__14954 (
            .O(N__69787),
            .I(\pid_front.N_259_cascade_ ));
    InMux I__14953 (
            .O(N__69784),
            .I(N__69781));
    LocalMux I__14952 (
            .O(N__69781),
            .I(N__69778));
    Span4Mux_v I__14951 (
            .O(N__69778),
            .I(N__69775));
    Span4Mux_h I__14950 (
            .O(N__69775),
            .I(N__69772));
    Odrv4 I__14949 (
            .O(N__69772),
            .I(\pid_front.N_111 ));
    InMux I__14948 (
            .O(N__69769),
            .I(N__69766));
    LocalMux I__14947 (
            .O(N__69766),
            .I(\pid_front.error_i_reg_9_1_14 ));
    CascadeMux I__14946 (
            .O(N__69763),
            .I(N__69760));
    InMux I__14945 (
            .O(N__69760),
            .I(N__69757));
    LocalMux I__14944 (
            .O(N__69757),
            .I(N__69754));
    Odrv4 I__14943 (
            .O(N__69754),
            .I(\pid_front.N_454 ));
    CascadeMux I__14942 (
            .O(N__69751),
            .I(\pid_front.N_515_cascade_ ));
    CascadeMux I__14941 (
            .O(N__69748),
            .I(\pid_front.N_450_cascade_ ));
    CascadeMux I__14940 (
            .O(N__69745),
            .I(\pid_front.m16_2_03_4_0_cascade_ ));
    CascadeMux I__14939 (
            .O(N__69742),
            .I(\pid_front.m16_2_03_4_cascade_ ));
    CascadeMux I__14938 (
            .O(N__69739),
            .I(N__69736));
    InMux I__14937 (
            .O(N__69736),
            .I(N__69733));
    LocalMux I__14936 (
            .O(N__69733),
            .I(N__69730));
    Span4Mux_h I__14935 (
            .O(N__69730),
            .I(N__69727));
    Odrv4 I__14934 (
            .O(N__69727),
            .I(\pid_front.error_i_regZ0Z_12 ));
    CascadeMux I__14933 (
            .O(N__69724),
            .I(\pid_front.m18_2_03_4_1_cascade_ ));
    InMux I__14932 (
            .O(N__69721),
            .I(N__69718));
    LocalMux I__14931 (
            .O(N__69718),
            .I(N__69715));
    Span4Mux_v I__14930 (
            .O(N__69715),
            .I(N__69712));
    Odrv4 I__14929 (
            .O(N__69712),
            .I(\pid_front.error_i_regZ0Z_14 ));
    InMux I__14928 (
            .O(N__69709),
            .I(N__69706));
    LocalMux I__14927 (
            .O(N__69706),
            .I(\pid_front.N_580 ));
    InMux I__14926 (
            .O(N__69703),
            .I(N__69696));
    InMux I__14925 (
            .O(N__69702),
            .I(N__69696));
    InMux I__14924 (
            .O(N__69701),
            .I(N__69693));
    LocalMux I__14923 (
            .O(N__69696),
            .I(N__69690));
    LocalMux I__14922 (
            .O(N__69693),
            .I(N__69687));
    Span4Mux_v I__14921 (
            .O(N__69690),
            .I(N__69684));
    Span4Mux_v I__14920 (
            .O(N__69687),
            .I(N__69681));
    Odrv4 I__14919 (
            .O(N__69684),
            .I(\pid_front.N_187 ));
    Odrv4 I__14918 (
            .O(N__69681),
            .I(\pid_front.N_187 ));
    InMux I__14917 (
            .O(N__69676),
            .I(N__69670));
    InMux I__14916 (
            .O(N__69675),
            .I(N__69670));
    LocalMux I__14915 (
            .O(N__69670),
            .I(\pid_front.N_263 ));
    InMux I__14914 (
            .O(N__69667),
            .I(N__69664));
    LocalMux I__14913 (
            .O(N__69664),
            .I(\pid_front.N_54_i_1 ));
    CascadeMux I__14912 (
            .O(N__69661),
            .I(\pid_front.N_54_i_1_cascade_ ));
    InMux I__14911 (
            .O(N__69658),
            .I(N__69654));
    InMux I__14910 (
            .O(N__69657),
            .I(N__69651));
    LocalMux I__14909 (
            .O(N__69654),
            .I(N__69648));
    LocalMux I__14908 (
            .O(N__69651),
            .I(N__69645));
    Span4Mux_v I__14907 (
            .O(N__69648),
            .I(N__69640));
    Span4Mux_v I__14906 (
            .O(N__69645),
            .I(N__69640));
    Odrv4 I__14905 (
            .O(N__69640),
            .I(\pid_side.N_2601_i ));
    InMux I__14904 (
            .O(N__69637),
            .I(N__69634));
    LocalMux I__14903 (
            .O(N__69634),
            .I(\pid_front.N_429 ));
    CascadeMux I__14902 (
            .O(N__69631),
            .I(\pid_front.N_332_cascade_ ));
    InMux I__14901 (
            .O(N__69628),
            .I(N__69625));
    LocalMux I__14900 (
            .O(N__69625),
            .I(\pid_front.N_262 ));
    CascadeMux I__14899 (
            .O(N__69622),
            .I(\pid_front.error_i_reg_esr_RNO_0Z0Z_17_cascade_ ));
    InMux I__14898 (
            .O(N__69619),
            .I(N__69616));
    LocalMux I__14897 (
            .O(N__69616),
            .I(N__69613));
    Span4Mux_v I__14896 (
            .O(N__69613),
            .I(N__69610));
    Span4Mux_v I__14895 (
            .O(N__69610),
            .I(N__69607));
    Sp12to4 I__14894 (
            .O(N__69607),
            .I(N__69604));
    Odrv12 I__14893 (
            .O(N__69604),
            .I(\pid_front.error_i_regZ0Z_17 ));
    InMux I__14892 (
            .O(N__69601),
            .I(N__69598));
    LocalMux I__14891 (
            .O(N__69598),
            .I(N__69595));
    Span4Mux_v I__14890 (
            .O(N__69595),
            .I(N__69591));
    InMux I__14889 (
            .O(N__69594),
            .I(N__69588));
    Odrv4 I__14888 (
            .O(N__69591),
            .I(\pid_front.N_6 ));
    LocalMux I__14887 (
            .O(N__69588),
            .I(\pid_front.N_6 ));
    InMux I__14886 (
            .O(N__69583),
            .I(N__69577));
    InMux I__14885 (
            .O(N__69582),
            .I(N__69574));
    InMux I__14884 (
            .O(N__69581),
            .I(N__69571));
    InMux I__14883 (
            .O(N__69580),
            .I(N__69568));
    LocalMux I__14882 (
            .O(N__69577),
            .I(N__69565));
    LocalMux I__14881 (
            .O(N__69574),
            .I(N__69562));
    LocalMux I__14880 (
            .O(N__69571),
            .I(N__69559));
    LocalMux I__14879 (
            .O(N__69568),
            .I(N__69556));
    Span4Mux_v I__14878 (
            .O(N__69565),
            .I(N__69553));
    Span4Mux_v I__14877 (
            .O(N__69562),
            .I(N__69545));
    Span4Mux_h I__14876 (
            .O(N__69559),
            .I(N__69545));
    Span4Mux_v I__14875 (
            .O(N__69556),
            .I(N__69545));
    Span4Mux_h I__14874 (
            .O(N__69553),
            .I(N__69542));
    InMux I__14873 (
            .O(N__69552),
            .I(N__69539));
    Odrv4 I__14872 (
            .O(N__69545),
            .I(\pid_front.m1_0_03 ));
    Odrv4 I__14871 (
            .O(N__69542),
            .I(\pid_front.m1_0_03 ));
    LocalMux I__14870 (
            .O(N__69539),
            .I(\pid_front.m1_0_03 ));
    InMux I__14869 (
            .O(N__69532),
            .I(N__69529));
    LocalMux I__14868 (
            .O(N__69529),
            .I(\pid_front.error_i_reg_esr_RNO_1Z0Z_17 ));
    InMux I__14867 (
            .O(N__69526),
            .I(N__69523));
    LocalMux I__14866 (
            .O(N__69523),
            .I(N__69520));
    Odrv4 I__14865 (
            .O(N__69520),
            .I(\pid_side.N_580 ));
    CascadeMux I__14864 (
            .O(N__69517),
            .I(\pid_side.N_156_cascade_ ));
    InMux I__14863 (
            .O(N__69514),
            .I(N__69511));
    LocalMux I__14862 (
            .O(N__69511),
            .I(\pid_side.N_182 ));
    CascadeMux I__14861 (
            .O(N__69508),
            .I(N__69505));
    InMux I__14860 (
            .O(N__69505),
            .I(N__69501));
    CascadeMux I__14859 (
            .O(N__69504),
            .I(N__69498));
    LocalMux I__14858 (
            .O(N__69501),
            .I(N__69495));
    InMux I__14857 (
            .O(N__69498),
            .I(N__69492));
    Span4Mux_h I__14856 (
            .O(N__69495),
            .I(N__69486));
    LocalMux I__14855 (
            .O(N__69492),
            .I(N__69486));
    InMux I__14854 (
            .O(N__69491),
            .I(N__69483));
    Span4Mux_v I__14853 (
            .O(N__69486),
            .I(N__69478));
    LocalMux I__14852 (
            .O(N__69483),
            .I(N__69475));
    InMux I__14851 (
            .O(N__69482),
            .I(N__69470));
    InMux I__14850 (
            .O(N__69481),
            .I(N__69470));
    Span4Mux_h I__14849 (
            .O(N__69478),
            .I(N__69467));
    Span4Mux_v I__14848 (
            .O(N__69475),
            .I(N__69464));
    LocalMux I__14847 (
            .O(N__69470),
            .I(N__69461));
    Span4Mux_v I__14846 (
            .O(N__69467),
            .I(N__69458));
    Odrv4 I__14845 (
            .O(N__69464),
            .I(pid_side_m10_2_03_3_i_0_a2_1_0));
    Odrv4 I__14844 (
            .O(N__69461),
            .I(pid_side_m10_2_03_3_i_0_a2_1_0));
    Odrv4 I__14843 (
            .O(N__69458),
            .I(pid_side_m10_2_03_3_i_0_a2_1_0));
    InMux I__14842 (
            .O(N__69451),
            .I(N__69448));
    LocalMux I__14841 (
            .O(N__69448),
            .I(\pid_side.N_549 ));
    CascadeMux I__14840 (
            .O(N__69445),
            .I(\pid_side.N_182_cascade_ ));
    InMux I__14839 (
            .O(N__69442),
            .I(N__69438));
    InMux I__14838 (
            .O(N__69441),
            .I(N__69435));
    LocalMux I__14837 (
            .O(N__69438),
            .I(N__69432));
    LocalMux I__14836 (
            .O(N__69435),
            .I(N__69429));
    Span4Mux_h I__14835 (
            .O(N__69432),
            .I(N__69424));
    Span4Mux_h I__14834 (
            .O(N__69429),
            .I(N__69424));
    Span4Mux_h I__14833 (
            .O(N__69424),
            .I(N__69421));
    Odrv4 I__14832 (
            .O(N__69421),
            .I(\Commands_frame_decoder.source_CH3data_1_sqmuxa ));
    InMux I__14831 (
            .O(N__69418),
            .I(N__69411));
    InMux I__14830 (
            .O(N__69417),
            .I(N__69411));
    InMux I__14829 (
            .O(N__69416),
            .I(N__69405));
    LocalMux I__14828 (
            .O(N__69411),
            .I(N__69402));
    InMux I__14827 (
            .O(N__69410),
            .I(N__69397));
    InMux I__14826 (
            .O(N__69409),
            .I(N__69397));
    InMux I__14825 (
            .O(N__69408),
            .I(N__69394));
    LocalMux I__14824 (
            .O(N__69405),
            .I(N__69389));
    Span4Mux_h I__14823 (
            .O(N__69402),
            .I(N__69386));
    LocalMux I__14822 (
            .O(N__69397),
            .I(N__69381));
    LocalMux I__14821 (
            .O(N__69394),
            .I(N__69381));
    InMux I__14820 (
            .O(N__69393),
            .I(N__69376));
    InMux I__14819 (
            .O(N__69392),
            .I(N__69376));
    Span4Mux_h I__14818 (
            .O(N__69389),
            .I(N__69368));
    Span4Mux_v I__14817 (
            .O(N__69386),
            .I(N__69361));
    Span4Mux_h I__14816 (
            .O(N__69381),
            .I(N__69361));
    LocalMux I__14815 (
            .O(N__69376),
            .I(N__69361));
    InMux I__14814 (
            .O(N__69375),
            .I(N__69350));
    InMux I__14813 (
            .O(N__69374),
            .I(N__69350));
    InMux I__14812 (
            .O(N__69373),
            .I(N__69350));
    InMux I__14811 (
            .O(N__69372),
            .I(N__69350));
    InMux I__14810 (
            .O(N__69371),
            .I(N__69350));
    Odrv4 I__14809 (
            .O(N__69368),
            .I(\Commands_frame_decoder.N_403 ));
    Odrv4 I__14808 (
            .O(N__69361),
            .I(\Commands_frame_decoder.N_403 ));
    LocalMux I__14807 (
            .O(N__69350),
            .I(\Commands_frame_decoder.N_403 ));
    InMux I__14806 (
            .O(N__69343),
            .I(N__69339));
    InMux I__14805 (
            .O(N__69342),
            .I(N__69336));
    LocalMux I__14804 (
            .O(N__69339),
            .I(N__69333));
    LocalMux I__14803 (
            .O(N__69336),
            .I(N__69330));
    Span4Mux_h I__14802 (
            .O(N__69333),
            .I(N__69327));
    Odrv4 I__14801 (
            .O(N__69330),
            .I(\Commands_frame_decoder.stateZ0Z_5 ));
    Odrv4 I__14800 (
            .O(N__69327),
            .I(\Commands_frame_decoder.stateZ0Z_5 ));
    InMux I__14799 (
            .O(N__69322),
            .I(N__69319));
    LocalMux I__14798 (
            .O(N__69319),
            .I(N__69316));
    Span4Mux_h I__14797 (
            .O(N__69316),
            .I(N__69312));
    InMux I__14796 (
            .O(N__69315),
            .I(N__69309));
    Sp12to4 I__14795 (
            .O(N__69312),
            .I(N__69304));
    LocalMux I__14794 (
            .O(N__69309),
            .I(N__69304));
    Span12Mux_h I__14793 (
            .O(N__69304),
            .I(N__69301));
    Odrv12 I__14792 (
            .O(N__69301),
            .I(\dron_frame_decoder_1.state_RNI6P6KZ0Z_4 ));
    InMux I__14791 (
            .O(N__69298),
            .I(N__69295));
    LocalMux I__14790 (
            .O(N__69295),
            .I(N__69292));
    Span4Mux_v I__14789 (
            .O(N__69292),
            .I(N__69287));
    InMux I__14788 (
            .O(N__69291),
            .I(N__69282));
    InMux I__14787 (
            .O(N__69290),
            .I(N__69282));
    Span4Mux_h I__14786 (
            .O(N__69287),
            .I(N__69279));
    LocalMux I__14785 (
            .O(N__69282),
            .I(N__69276));
    Span4Mux_h I__14784 (
            .O(N__69279),
            .I(N__69269));
    Span4Mux_v I__14783 (
            .O(N__69276),
            .I(N__69266));
    InMux I__14782 (
            .O(N__69275),
            .I(N__69261));
    InMux I__14781 (
            .O(N__69274),
            .I(N__69261));
    InMux I__14780 (
            .O(N__69273),
            .I(N__69256));
    InMux I__14779 (
            .O(N__69272),
            .I(N__69256));
    Odrv4 I__14778 (
            .O(N__69269),
            .I(\dron_frame_decoder_1.N_218 ));
    Odrv4 I__14777 (
            .O(N__69266),
            .I(\dron_frame_decoder_1.N_218 ));
    LocalMux I__14776 (
            .O(N__69261),
            .I(\dron_frame_decoder_1.N_218 ));
    LocalMux I__14775 (
            .O(N__69256),
            .I(\dron_frame_decoder_1.N_218 ));
    CascadeMux I__14774 (
            .O(N__69247),
            .I(N__69243));
    CascadeMux I__14773 (
            .O(N__69246),
            .I(N__69240));
    InMux I__14772 (
            .O(N__69243),
            .I(N__69237));
    InMux I__14771 (
            .O(N__69240),
            .I(N__69234));
    LocalMux I__14770 (
            .O(N__69237),
            .I(N__69231));
    LocalMux I__14769 (
            .O(N__69234),
            .I(N__69228));
    Span4Mux_v I__14768 (
            .O(N__69231),
            .I(N__69223));
    Span4Mux_v I__14767 (
            .O(N__69228),
            .I(N__69223));
    Span4Mux_h I__14766 (
            .O(N__69223),
            .I(N__69219));
    InMux I__14765 (
            .O(N__69222),
            .I(N__69216));
    Span4Mux_h I__14764 (
            .O(N__69219),
            .I(N__69213));
    LocalMux I__14763 (
            .O(N__69216),
            .I(N__69210));
    Span4Mux_v I__14762 (
            .O(N__69213),
            .I(N__69207));
    Odrv4 I__14761 (
            .O(N__69210),
            .I(\dron_frame_decoder_1.stateZ0Z_7 ));
    Odrv4 I__14760 (
            .O(N__69207),
            .I(\dron_frame_decoder_1.stateZ0Z_7 ));
    IoInMux I__14759 (
            .O(N__69202),
            .I(N__69199));
    LocalMux I__14758 (
            .O(N__69199),
            .I(N__69195));
    InMux I__14757 (
            .O(N__69198),
            .I(N__69192));
    Span4Mux_s3_v I__14756 (
            .O(N__69195),
            .I(N__69187));
    LocalMux I__14755 (
            .O(N__69192),
            .I(N__69184));
    CascadeMux I__14754 (
            .O(N__69191),
            .I(N__69179));
    CascadeMux I__14753 (
            .O(N__69190),
            .I(N__69174));
    Span4Mux_v I__14752 (
            .O(N__69187),
            .I(N__69171));
    Span4Mux_v I__14751 (
            .O(N__69184),
            .I(N__69168));
    InMux I__14750 (
            .O(N__69183),
            .I(N__69165));
    InMux I__14749 (
            .O(N__69182),
            .I(N__69162));
    InMux I__14748 (
            .O(N__69179),
            .I(N__69159));
    InMux I__14747 (
            .O(N__69178),
            .I(N__69156));
    InMux I__14746 (
            .O(N__69177),
            .I(N__69151));
    InMux I__14745 (
            .O(N__69174),
            .I(N__69151));
    Span4Mux_v I__14744 (
            .O(N__69171),
            .I(N__69147));
    Span4Mux_h I__14743 (
            .O(N__69168),
            .I(N__69142));
    LocalMux I__14742 (
            .O(N__69165),
            .I(N__69142));
    LocalMux I__14741 (
            .O(N__69162),
            .I(N__69139));
    LocalMux I__14740 (
            .O(N__69159),
            .I(N__69132));
    LocalMux I__14739 (
            .O(N__69156),
            .I(N__69132));
    LocalMux I__14738 (
            .O(N__69151),
            .I(N__69132));
    InMux I__14737 (
            .O(N__69150),
            .I(N__69129));
    Span4Mux_h I__14736 (
            .O(N__69147),
            .I(N__69124));
    Span4Mux_h I__14735 (
            .O(N__69142),
            .I(N__69124));
    Span4Mux_v I__14734 (
            .O(N__69139),
            .I(N__69121));
    Span4Mux_h I__14733 (
            .O(N__69132),
            .I(N__69118));
    LocalMux I__14732 (
            .O(N__69129),
            .I(N__69115));
    Span4Mux_v I__14731 (
            .O(N__69124),
            .I(N__69112));
    Span4Mux_v I__14730 (
            .O(N__69121),
            .I(N__69109));
    Span4Mux_v I__14729 (
            .O(N__69118),
            .I(N__69106));
    Span4Mux_h I__14728 (
            .O(N__69115),
            .I(N__69101));
    Span4Mux_v I__14727 (
            .O(N__69112),
            .I(N__69098));
    Span4Mux_h I__14726 (
            .O(N__69109),
            .I(N__69093));
    Span4Mux_v I__14725 (
            .O(N__69106),
            .I(N__69093));
    InMux I__14724 (
            .O(N__69105),
            .I(N__69088));
    InMux I__14723 (
            .O(N__69104),
            .I(N__69088));
    Odrv4 I__14722 (
            .O(N__69101),
            .I(debug_CH1_0A_c));
    Odrv4 I__14721 (
            .O(N__69098),
            .I(debug_CH1_0A_c));
    Odrv4 I__14720 (
            .O(N__69093),
            .I(debug_CH1_0A_c));
    LocalMux I__14719 (
            .O(N__69088),
            .I(debug_CH1_0A_c));
    CascadeMux I__14718 (
            .O(N__69079),
            .I(N__69074));
    InMux I__14717 (
            .O(N__69078),
            .I(N__69071));
    InMux I__14716 (
            .O(N__69077),
            .I(N__69068));
    InMux I__14715 (
            .O(N__69074),
            .I(N__69065));
    LocalMux I__14714 (
            .O(N__69071),
            .I(N__69062));
    LocalMux I__14713 (
            .O(N__69068),
            .I(N__69059));
    LocalMux I__14712 (
            .O(N__69065),
            .I(N__69056));
    Span4Mux_v I__14711 (
            .O(N__69062),
            .I(N__69053));
    Span4Mux_v I__14710 (
            .O(N__69059),
            .I(N__69050));
    Span4Mux_v I__14709 (
            .O(N__69056),
            .I(N__69047));
    Span4Mux_h I__14708 (
            .O(N__69053),
            .I(N__69038));
    Span4Mux_v I__14707 (
            .O(N__69050),
            .I(N__69038));
    Span4Mux_v I__14706 (
            .O(N__69047),
            .I(N__69038));
    InMux I__14705 (
            .O(N__69046),
            .I(N__69033));
    InMux I__14704 (
            .O(N__69045),
            .I(N__69033));
    Span4Mux_h I__14703 (
            .O(N__69038),
            .I(N__69030));
    LocalMux I__14702 (
            .O(N__69033),
            .I(\pid_alt.stateZ0Z_0 ));
    Odrv4 I__14701 (
            .O(N__69030),
            .I(\pid_alt.stateZ0Z_0 ));
    CascadeMux I__14700 (
            .O(N__69025),
            .I(N__69015));
    CascadeMux I__14699 (
            .O(N__69024),
            .I(N__69005));
    InMux I__14698 (
            .O(N__69023),
            .I(N__68985));
    InMux I__14697 (
            .O(N__69022),
            .I(N__68985));
    InMux I__14696 (
            .O(N__69021),
            .I(N__68985));
    InMux I__14695 (
            .O(N__69020),
            .I(N__68985));
    InMux I__14694 (
            .O(N__69019),
            .I(N__68985));
    InMux I__14693 (
            .O(N__69018),
            .I(N__68985));
    InMux I__14692 (
            .O(N__69015),
            .I(N__68985));
    InMux I__14691 (
            .O(N__69014),
            .I(N__68985));
    InMux I__14690 (
            .O(N__69013),
            .I(N__68980));
    InMux I__14689 (
            .O(N__69012),
            .I(N__68980));
    InMux I__14688 (
            .O(N__69011),
            .I(N__68976));
    InMux I__14687 (
            .O(N__69010),
            .I(N__68961));
    InMux I__14686 (
            .O(N__69009),
            .I(N__68961));
    InMux I__14685 (
            .O(N__69008),
            .I(N__68961));
    InMux I__14684 (
            .O(N__69005),
            .I(N__68961));
    InMux I__14683 (
            .O(N__69004),
            .I(N__68961));
    InMux I__14682 (
            .O(N__69003),
            .I(N__68961));
    InMux I__14681 (
            .O(N__69002),
            .I(N__68961));
    LocalMux I__14680 (
            .O(N__68985),
            .I(N__68955));
    LocalMux I__14679 (
            .O(N__68980),
            .I(N__68952));
    InMux I__14678 (
            .O(N__68979),
            .I(N__68949));
    LocalMux I__14677 (
            .O(N__68976),
            .I(N__68946));
    LocalMux I__14676 (
            .O(N__68961),
            .I(N__68943));
    InMux I__14675 (
            .O(N__68960),
            .I(N__68936));
    InMux I__14674 (
            .O(N__68959),
            .I(N__68936));
    InMux I__14673 (
            .O(N__68958),
            .I(N__68936));
    Span4Mux_h I__14672 (
            .O(N__68955),
            .I(N__68931));
    Span4Mux_v I__14671 (
            .O(N__68952),
            .I(N__68931));
    LocalMux I__14670 (
            .O(N__68949),
            .I(N__68928));
    Span4Mux_v I__14669 (
            .O(N__68946),
            .I(N__68921));
    Span4Mux_h I__14668 (
            .O(N__68943),
            .I(N__68921));
    LocalMux I__14667 (
            .O(N__68936),
            .I(N__68921));
    Span4Mux_h I__14666 (
            .O(N__68931),
            .I(N__68916));
    Span4Mux_v I__14665 (
            .O(N__68928),
            .I(N__68916));
    Span4Mux_v I__14664 (
            .O(N__68921),
            .I(N__68913));
    Span4Mux_v I__14663 (
            .O(N__68916),
            .I(N__68907));
    Span4Mux_h I__14662 (
            .O(N__68913),
            .I(N__68907));
    InMux I__14661 (
            .O(N__68912),
            .I(N__68904));
    Span4Mux_h I__14660 (
            .O(N__68907),
            .I(N__68901));
    LocalMux I__14659 (
            .O(N__68904),
            .I(\pid_alt.N_72_i ));
    Odrv4 I__14658 (
            .O(N__68901),
            .I(\pid_alt.N_72_i ));
    InMux I__14657 (
            .O(N__68896),
            .I(N__68893));
    LocalMux I__14656 (
            .O(N__68893),
            .I(N__68890));
    Span4Mux_v I__14655 (
            .O(N__68890),
            .I(N__68887));
    Span4Mux_h I__14654 (
            .O(N__68887),
            .I(N__68884));
    Span4Mux_v I__14653 (
            .O(N__68884),
            .I(N__68881));
    Odrv4 I__14652 (
            .O(N__68881),
            .I(\pid_front.error_p_reg_esr_RNICMVCGZ0Z_14 ));
    InMux I__14651 (
            .O(N__68878),
            .I(N__68875));
    LocalMux I__14650 (
            .O(N__68875),
            .I(\pid_side.error_i_reg_esr_RNO_1_0_17 ));
    InMux I__14649 (
            .O(N__68872),
            .I(N__68869));
    LocalMux I__14648 (
            .O(N__68869),
            .I(N__68866));
    Span4Mux_h I__14647 (
            .O(N__68866),
            .I(N__68863));
    Odrv4 I__14646 (
            .O(N__68863),
            .I(\pid_side.error_i_regZ0Z_17 ));
    InMux I__14645 (
            .O(N__68860),
            .I(N__68857));
    LocalMux I__14644 (
            .O(N__68857),
            .I(\pid_side.m16_2_03_4 ));
    CascadeMux I__14643 (
            .O(N__68854),
            .I(\pid_side.m0_2_03_cascade_ ));
    CascadeMux I__14642 (
            .O(N__68851),
            .I(N__68848));
    InMux I__14641 (
            .O(N__68848),
            .I(N__68845));
    LocalMux I__14640 (
            .O(N__68845),
            .I(N__68842));
    Span4Mux_h I__14639 (
            .O(N__68842),
            .I(N__68839));
    Odrv4 I__14638 (
            .O(N__68839),
            .I(\pid_side.error_i_regZ0Z_12 ));
    CascadeMux I__14637 (
            .O(N__68836),
            .I(\pid_side.m1_0_03_cascade_ ));
    InMux I__14636 (
            .O(N__68833),
            .I(N__68830));
    LocalMux I__14635 (
            .O(N__68830),
            .I(N__68827));
    Odrv4 I__14634 (
            .O(N__68827),
            .I(\pid_side.error_i_reg_9_rn_1_13 ));
    CascadeMux I__14633 (
            .O(N__68824),
            .I(\pid_side.N_232_cascade_ ));
    CascadeMux I__14632 (
            .O(N__68821),
            .I(\pid_side.N_549_cascade_ ));
    CascadeMux I__14631 (
            .O(N__68818),
            .I(\pid_side.error_i_reg_esr_RNO_0_0_6_cascade_ ));
    CascadeMux I__14630 (
            .O(N__68815),
            .I(N__68812));
    InMux I__14629 (
            .O(N__68812),
            .I(N__68809));
    LocalMux I__14628 (
            .O(N__68809),
            .I(N__68806));
    Span4Mux_h I__14627 (
            .O(N__68806),
            .I(N__68803));
    Sp12to4 I__14626 (
            .O(N__68803),
            .I(N__68800));
    Odrv12 I__14625 (
            .O(N__68800),
            .I(\pid_side.error_i_regZ0Z_6 ));
    InMux I__14624 (
            .O(N__68797),
            .I(N__68794));
    LocalMux I__14623 (
            .O(N__68794),
            .I(\pid_side.m78_0_1 ));
    CascadeMux I__14622 (
            .O(N__68791),
            .I(\pid_side.m78_0_0_cascade_ ));
    CascadeMux I__14621 (
            .O(N__68788),
            .I(N__68785));
    InMux I__14620 (
            .O(N__68785),
            .I(N__68782));
    LocalMux I__14619 (
            .O(N__68782),
            .I(N__68779));
    Span4Mux_h I__14618 (
            .O(N__68779),
            .I(N__68776));
    Odrv4 I__14617 (
            .O(N__68776),
            .I(\pid_side.error_i_regZ0Z_11 ));
    InMux I__14616 (
            .O(N__68773),
            .I(N__68770));
    LocalMux I__14615 (
            .O(N__68770),
            .I(\pid_side.N_626 ));
    CascadeMux I__14614 (
            .O(N__68767),
            .I(\pid_side.N_626_cascade_ ));
    InMux I__14613 (
            .O(N__68764),
            .I(N__68761));
    LocalMux I__14612 (
            .O(N__68761),
            .I(\pid_side.N_398 ));
    CascadeMux I__14611 (
            .O(N__68758),
            .I(\pid_side.N_161_cascade_ ));
    InMux I__14610 (
            .O(N__68755),
            .I(N__68752));
    LocalMux I__14609 (
            .O(N__68752),
            .I(\pid_side.m13_2_03_4_i_0_o2_2_1 ));
    InMux I__14608 (
            .O(N__68749),
            .I(N__68746));
    LocalMux I__14607 (
            .O(N__68746),
            .I(N__68742));
    InMux I__14606 (
            .O(N__68745),
            .I(N__68739));
    Odrv4 I__14605 (
            .O(N__68742),
            .I(\pid_side.N_594 ));
    LocalMux I__14604 (
            .O(N__68739),
            .I(\pid_side.N_594 ));
    CascadeMux I__14603 (
            .O(N__68734),
            .I(\pid_side.N_594_cascade_ ));
    CascadeMux I__14602 (
            .O(N__68731),
            .I(\pid_side.error_i_reg_9_sn_13_cascade_ ));
    CascadeMux I__14601 (
            .O(N__68728),
            .I(N__68725));
    InMux I__14600 (
            .O(N__68725),
            .I(N__68722));
    LocalMux I__14599 (
            .O(N__68722),
            .I(N__68719));
    Span4Mux_h I__14598 (
            .O(N__68719),
            .I(N__68716));
    Odrv4 I__14597 (
            .O(N__68716),
            .I(\pid_side.error_i_regZ0Z_13 ));
    InMux I__14596 (
            .O(N__68713),
            .I(N__68709));
    InMux I__14595 (
            .O(N__68712),
            .I(N__68706));
    LocalMux I__14594 (
            .O(N__68709),
            .I(N__68703));
    LocalMux I__14593 (
            .O(N__68706),
            .I(N__68700));
    Span4Mux_v I__14592 (
            .O(N__68703),
            .I(N__68696));
    Span4Mux_v I__14591 (
            .O(N__68700),
            .I(N__68693));
    InMux I__14590 (
            .O(N__68699),
            .I(N__68690));
    Odrv4 I__14589 (
            .O(N__68696),
            .I(xy_ki_5));
    Odrv4 I__14588 (
            .O(N__68693),
            .I(xy_ki_5));
    LocalMux I__14587 (
            .O(N__68690),
            .I(xy_ki_5));
    CascadeMux I__14586 (
            .O(N__68683),
            .I(pid_side_N_490_cascade_));
    CascadeMux I__14585 (
            .O(N__68680),
            .I(\pid_side.m78_0_a2_sx_cascade_ ));
    InMux I__14584 (
            .O(N__68677),
            .I(N__68674));
    LocalMux I__14583 (
            .O(N__68674),
            .I(\pid_side.N_394 ));
    InMux I__14582 (
            .O(N__68671),
            .I(N__68667));
    InMux I__14581 (
            .O(N__68670),
            .I(N__68664));
    LocalMux I__14580 (
            .O(N__68667),
            .I(N__68661));
    LocalMux I__14579 (
            .O(N__68664),
            .I(N__68658));
    Span4Mux_h I__14578 (
            .O(N__68661),
            .I(N__68655));
    Odrv12 I__14577 (
            .O(N__68658),
            .I(pid_side_m78_0_a2_0_0));
    Odrv4 I__14576 (
            .O(N__68655),
            .I(pid_side_m78_0_a2_0_0));
    InMux I__14575 (
            .O(N__68650),
            .I(N__68646));
    InMux I__14574 (
            .O(N__68649),
            .I(N__68643));
    LocalMux I__14573 (
            .O(N__68646),
            .I(N__68640));
    LocalMux I__14572 (
            .O(N__68643),
            .I(N__68637));
    Span4Mux_h I__14571 (
            .O(N__68640),
            .I(N__68634));
    Span4Mux_h I__14570 (
            .O(N__68637),
            .I(N__68629));
    Span4Mux_v I__14569 (
            .O(N__68634),
            .I(N__68629));
    Odrv4 I__14568 (
            .O(N__68629),
            .I(\pid_side.error_d_reg_prev_esr_RNI9LLC4Z0Z_12 ));
    CascadeMux I__14567 (
            .O(N__68626),
            .I(\pid_side.error_d_reg_prev_esr_RNID3GT3Z0Z_10_cascade_ ));
    InMux I__14566 (
            .O(N__68623),
            .I(N__68619));
    InMux I__14565 (
            .O(N__68622),
            .I(N__68616));
    LocalMux I__14564 (
            .O(N__68619),
            .I(\pid_side.error_p_reg_esr_RNIL0VP1Z0Z_12 ));
    LocalMux I__14563 (
            .O(N__68616),
            .I(\pid_side.error_p_reg_esr_RNIL0VP1Z0Z_12 ));
    CascadeMux I__14562 (
            .O(N__68611),
            .I(N__68608));
    InMux I__14561 (
            .O(N__68608),
            .I(N__68605));
    LocalMux I__14560 (
            .O(N__68605),
            .I(N__68602));
    Span4Mux_v I__14559 (
            .O(N__68602),
            .I(N__68599));
    Odrv4 I__14558 (
            .O(N__68599),
            .I(\pid_side.error_d_reg_prev_esr_RNIUOPVAZ0Z_10 ));
    CascadeMux I__14557 (
            .O(N__68596),
            .I(\pid_side.un1_pid_prereg_167_0_cascade_ ));
    InMux I__14556 (
            .O(N__68593),
            .I(N__68590));
    LocalMux I__14555 (
            .O(N__68590),
            .I(N__68585));
    InMux I__14554 (
            .O(N__68589),
            .I(N__68580));
    InMux I__14553 (
            .O(N__68588),
            .I(N__68580));
    Span4Mux_h I__14552 (
            .O(N__68585),
            .I(N__68577));
    LocalMux I__14551 (
            .O(N__68580),
            .I(N__68574));
    Odrv4 I__14550 (
            .O(N__68577),
            .I(\pid_side.error_d_reg_prev_esr_RNI59QR8Z0Z_12 ));
    Odrv12 I__14549 (
            .O(N__68574),
            .I(\pid_side.error_d_reg_prev_esr_RNI59QR8Z0Z_12 ));
    InMux I__14548 (
            .O(N__68569),
            .I(N__68566));
    LocalMux I__14547 (
            .O(N__68566),
            .I(\pid_side.un1_pid_prereg_167_0_1 ));
    InMux I__14546 (
            .O(N__68563),
            .I(N__68558));
    InMux I__14545 (
            .O(N__68562),
            .I(N__68553));
    InMux I__14544 (
            .O(N__68561),
            .I(N__68553));
    LocalMux I__14543 (
            .O(N__68558),
            .I(\pid_side.un1_pid_prereg_79 ));
    LocalMux I__14542 (
            .O(N__68553),
            .I(\pid_side.un1_pid_prereg_79 ));
    CascadeMux I__14541 (
            .O(N__68548),
            .I(\pid_side.error_d_reg_fast_esr_RNIPEC11Z0Z_12_cascade_ ));
    CascadeMux I__14540 (
            .O(N__68545),
            .I(\pid_side.error_d_reg_fast_esr_RNIEIJH2Z0Z_12_cascade_ ));
    InMux I__14539 (
            .O(N__68542),
            .I(N__68539));
    LocalMux I__14538 (
            .O(N__68539),
            .I(N__68535));
    InMux I__14537 (
            .O(N__68538),
            .I(N__68532));
    Span4Mux_h I__14536 (
            .O(N__68535),
            .I(N__68529));
    LocalMux I__14535 (
            .O(N__68532),
            .I(\pid_side.error_d_reg_prev_esr_RNIJHVG3Z0Z_12 ));
    Odrv4 I__14534 (
            .O(N__68529),
            .I(\pid_side.error_d_reg_prev_esr_RNIJHVG3Z0Z_12 ));
    InMux I__14533 (
            .O(N__68524),
            .I(N__68521));
    LocalMux I__14532 (
            .O(N__68521),
            .I(\pid_side.error_d_reg_fast_esr_RNIPHKNZ0Z_12 ));
    InMux I__14531 (
            .O(N__68518),
            .I(N__68512));
    InMux I__14530 (
            .O(N__68517),
            .I(N__68512));
    LocalMux I__14529 (
            .O(N__68512),
            .I(N__68509));
    Span4Mux_h I__14528 (
            .O(N__68509),
            .I(N__68506));
    Odrv4 I__14527 (
            .O(N__68506),
            .I(\pid_side.error_d_reg_esr_RNI2OIOZ0Z_13 ));
    CascadeMux I__14526 (
            .O(N__68503),
            .I(N__68499));
    InMux I__14525 (
            .O(N__68502),
            .I(N__68491));
    InMux I__14524 (
            .O(N__68499),
            .I(N__68491));
    InMux I__14523 (
            .O(N__68498),
            .I(N__68491));
    LocalMux I__14522 (
            .O(N__68491),
            .I(N__68488));
    Odrv4 I__14521 (
            .O(N__68488),
            .I(\pid_side.error_d_reg_fast_esr_RNIFGGE_0Z0Z_13 ));
    CascadeMux I__14520 (
            .O(N__68485),
            .I(N__68481));
    InMux I__14519 (
            .O(N__68484),
            .I(N__68478));
    InMux I__14518 (
            .O(N__68481),
            .I(N__68475));
    LocalMux I__14517 (
            .O(N__68478),
            .I(N__68470));
    LocalMux I__14516 (
            .O(N__68475),
            .I(N__68470));
    Span4Mux_h I__14515 (
            .O(N__68470),
            .I(N__68467));
    Odrv4 I__14514 (
            .O(N__68467),
            .I(\pid_side.error_d_reg_prev_esr_RNI5RIO_0Z0Z_14 ));
    InMux I__14513 (
            .O(N__68464),
            .I(N__68461));
    LocalMux I__14512 (
            .O(N__68461),
            .I(\pid_side.error_d_reg_fast_esr_RNIEIJH2Z0Z_12 ));
    InMux I__14511 (
            .O(N__68458),
            .I(N__68455));
    LocalMux I__14510 (
            .O(N__68455),
            .I(\pid_side.error_d_reg_prev_esr_RNI4M9H4Z0Z_14 ));
    InMux I__14509 (
            .O(N__68452),
            .I(N__68449));
    LocalMux I__14508 (
            .O(N__68449),
            .I(N__68446));
    Odrv4 I__14507 (
            .O(N__68446),
            .I(\pid_side.error_d_reg_prev_esr_RNIOVFK9Z0Z_17 ));
    InMux I__14506 (
            .O(N__68443),
            .I(N__68440));
    LocalMux I__14505 (
            .O(N__68440),
            .I(N__68437));
    Span4Mux_h I__14504 (
            .O(N__68437),
            .I(N__68433));
    InMux I__14503 (
            .O(N__68436),
            .I(N__68430));
    Odrv4 I__14502 (
            .O(N__68433),
            .I(\pid_side.un1_pid_prereg_0_18 ));
    LocalMux I__14501 (
            .O(N__68430),
            .I(\pid_side.un1_pid_prereg_0_18 ));
    CascadeMux I__14500 (
            .O(N__68425),
            .I(N__68422));
    InMux I__14499 (
            .O(N__68422),
            .I(N__68419));
    LocalMux I__14498 (
            .O(N__68419),
            .I(N__68416));
    Odrv4 I__14497 (
            .O(N__68416),
            .I(\pid_side.error_d_reg_prev_esr_RNII83B3Z0Z_21 ));
    CascadeMux I__14496 (
            .O(N__68413),
            .I(\pid_side.error_p_reg_esr_RNI4O091_0Z0Z_10_cascade_ ));
    CascadeMux I__14495 (
            .O(N__68410),
            .I(\pid_side.error_d_reg_prev_esr_RNIV62K2Z0Z_10_cascade_ ));
    InMux I__14494 (
            .O(N__68407),
            .I(N__68404));
    LocalMux I__14493 (
            .O(N__68404),
            .I(\pid_side.error_p_reg_esr_RNI4O091Z0Z_10 ));
    CascadeMux I__14492 (
            .O(N__68401),
            .I(\pid_side.un1_pid_prereg_153_0_cascade_ ));
    InMux I__14491 (
            .O(N__68398),
            .I(N__68395));
    LocalMux I__14490 (
            .O(N__68395),
            .I(N__68392));
    Span4Mux_h I__14489 (
            .O(N__68392),
            .I(N__68389));
    Odrv4 I__14488 (
            .O(N__68389),
            .I(\pid_side.error_d_reg_prev_esr_RNII28CBZ0Z_10 ));
    InMux I__14487 (
            .O(N__68386),
            .I(N__68383));
    LocalMux I__14486 (
            .O(N__68383),
            .I(\pid_side.error_d_reg_prev_esr_RNIV62K2Z0Z_10 ));
    InMux I__14485 (
            .O(N__68380),
            .I(N__68377));
    LocalMux I__14484 (
            .O(N__68377),
            .I(\pid_side.error_d_reg_prev_esr_RNID3GT3Z0Z_10 ));
    InMux I__14483 (
            .O(N__68374),
            .I(N__68371));
    LocalMux I__14482 (
            .O(N__68371),
            .I(N__68366));
    InMux I__14481 (
            .O(N__68370),
            .I(N__68361));
    InMux I__14480 (
            .O(N__68369),
            .I(N__68361));
    Span4Mux_h I__14479 (
            .O(N__68366),
            .I(N__68358));
    LocalMux I__14478 (
            .O(N__68361),
            .I(N__68355));
    Odrv4 I__14477 (
            .O(N__68358),
            .I(\pid_side.error_i_reg_esr_RNIJVKRZ0Z_12 ));
    Odrv4 I__14476 (
            .O(N__68355),
            .I(\pid_side.error_i_reg_esr_RNIJVKRZ0Z_12 ));
    InMux I__14475 (
            .O(N__68350),
            .I(N__68347));
    LocalMux I__14474 (
            .O(N__68347),
            .I(N__68344));
    Span4Mux_h I__14473 (
            .O(N__68344),
            .I(N__68341));
    Span4Mux_h I__14472 (
            .O(N__68341),
            .I(N__68337));
    InMux I__14471 (
            .O(N__68340),
            .I(N__68334));
    Odrv4 I__14470 (
            .O(N__68337),
            .I(\pid_side.un1_pid_prereg_0_22 ));
    LocalMux I__14469 (
            .O(N__68334),
            .I(\pid_side.un1_pid_prereg_0_22 ));
    CascadeMux I__14468 (
            .O(N__68329),
            .I(\pid_side.un1_pid_prereg_0_24_cascade_ ));
    InMux I__14467 (
            .O(N__68326),
            .I(N__68323));
    LocalMux I__14466 (
            .O(N__68323),
            .I(N__68320));
    Span4Mux_h I__14465 (
            .O(N__68320),
            .I(N__68315));
    InMux I__14464 (
            .O(N__68319),
            .I(N__68310));
    InMux I__14463 (
            .O(N__68318),
            .I(N__68310));
    Odrv4 I__14462 (
            .O(N__68315),
            .I(\pid_side.un1_pid_prereg_0_23 ));
    LocalMux I__14461 (
            .O(N__68310),
            .I(\pid_side.un1_pid_prereg_0_23 ));
    InMux I__14460 (
            .O(N__68305),
            .I(N__68302));
    LocalMux I__14459 (
            .O(N__68302),
            .I(\pid_side.error_d_reg_prev_esr_RNINEHM6Z0Z_21 ));
    InMux I__14458 (
            .O(N__68299),
            .I(N__68296));
    LocalMux I__14457 (
            .O(N__68296),
            .I(\pid_side.error_d_reg_prev_esr_RNIRLKM6Z0Z_21 ));
    InMux I__14456 (
            .O(N__68293),
            .I(N__68289));
    InMux I__14455 (
            .O(N__68292),
            .I(N__68286));
    LocalMux I__14454 (
            .O(N__68289),
            .I(\pid_side.un1_pid_prereg_0_15 ));
    LocalMux I__14453 (
            .O(N__68286),
            .I(\pid_side.un1_pid_prereg_0_15 ));
    InMux I__14452 (
            .O(N__68281),
            .I(N__68276));
    InMux I__14451 (
            .O(N__68280),
            .I(N__68271));
    InMux I__14450 (
            .O(N__68279),
            .I(N__68271));
    LocalMux I__14449 (
            .O(N__68276),
            .I(\pid_side.un1_pid_prereg_0_14 ));
    LocalMux I__14448 (
            .O(N__68271),
            .I(\pid_side.un1_pid_prereg_0_14 ));
    CascadeMux I__14447 (
            .O(N__68266),
            .I(\pid_side.un1_pid_prereg_0_17_cascade_ ));
    CascadeMux I__14446 (
            .O(N__68263),
            .I(N__68260));
    InMux I__14445 (
            .O(N__68260),
            .I(N__68257));
    LocalMux I__14444 (
            .O(N__68257),
            .I(\pid_side.error_d_reg_prev_esr_RNIOUVL6Z0Z_21 ));
    InMux I__14443 (
            .O(N__68254),
            .I(N__68249));
    InMux I__14442 (
            .O(N__68253),
            .I(N__68246));
    InMux I__14441 (
            .O(N__68252),
            .I(N__68243));
    LocalMux I__14440 (
            .O(N__68249),
            .I(N__68240));
    LocalMux I__14439 (
            .O(N__68246),
            .I(N__68235));
    LocalMux I__14438 (
            .O(N__68243),
            .I(N__68235));
    Span4Mux_v I__14437 (
            .O(N__68240),
            .I(N__68232));
    Span4Mux_h I__14436 (
            .O(N__68235),
            .I(N__68229));
    Odrv4 I__14435 (
            .O(N__68232),
            .I(\pid_side.error_i_reg_esr_RNIO8QSZ0Z_23 ));
    Odrv4 I__14434 (
            .O(N__68229),
            .I(\pid_side.error_i_reg_esr_RNIO8QSZ0Z_23 ));
    InMux I__14433 (
            .O(N__68224),
            .I(N__68221));
    LocalMux I__14432 (
            .O(N__68221),
            .I(N__68218));
    Span4Mux_v I__14431 (
            .O(N__68218),
            .I(N__68214));
    InMux I__14430 (
            .O(N__68217),
            .I(N__68211));
    Odrv4 I__14429 (
            .O(N__68214),
            .I(\pid_side.un1_pid_prereg_0_4 ));
    LocalMux I__14428 (
            .O(N__68211),
            .I(\pid_side.un1_pid_prereg_0_4 ));
    CascadeMux I__14427 (
            .O(N__68206),
            .I(N__68203));
    InMux I__14426 (
            .O(N__68203),
            .I(N__68200));
    LocalMux I__14425 (
            .O(N__68200),
            .I(N__68197));
    Span4Mux_v I__14424 (
            .O(N__68197),
            .I(N__68193));
    InMux I__14423 (
            .O(N__68196),
            .I(N__68190));
    Odrv4 I__14422 (
            .O(N__68193),
            .I(\pid_side.un1_pid_prereg_0_5 ));
    LocalMux I__14421 (
            .O(N__68190),
            .I(\pid_side.un1_pid_prereg_0_5 ));
    InMux I__14420 (
            .O(N__68185),
            .I(N__68182));
    LocalMux I__14419 (
            .O(N__68182),
            .I(N__68179));
    Odrv4 I__14418 (
            .O(N__68179),
            .I(\pid_side.error_d_reg_prev_esr_RNISR7K9Z0Z_16 ));
    InMux I__14417 (
            .O(N__68176),
            .I(N__68170));
    InMux I__14416 (
            .O(N__68175),
            .I(N__68170));
    LocalMux I__14415 (
            .O(N__68170),
            .I(N__68166));
    InMux I__14414 (
            .O(N__68169),
            .I(N__68163));
    Span4Mux_h I__14413 (
            .O(N__68166),
            .I(N__68160));
    LocalMux I__14412 (
            .O(N__68163),
            .I(\pid_side.error_i_reg_esr_RNIQBRSZ0Z_24 ));
    Odrv4 I__14411 (
            .O(N__68160),
            .I(\pid_side.error_i_reg_esr_RNIQBRSZ0Z_24 ));
    InMux I__14410 (
            .O(N__68155),
            .I(N__68151));
    InMux I__14409 (
            .O(N__68154),
            .I(N__68148));
    LocalMux I__14408 (
            .O(N__68151),
            .I(\pid_side.un1_pid_prereg_0_17 ));
    LocalMux I__14407 (
            .O(N__68148),
            .I(\pid_side.un1_pid_prereg_0_17 ));
    InMux I__14406 (
            .O(N__68143),
            .I(N__68138));
    InMux I__14405 (
            .O(N__68142),
            .I(N__68133));
    InMux I__14404 (
            .O(N__68141),
            .I(N__68133));
    LocalMux I__14403 (
            .O(N__68138),
            .I(\pid_side.un1_pid_prereg_0_16 ));
    LocalMux I__14402 (
            .O(N__68133),
            .I(\pid_side.un1_pid_prereg_0_16 ));
    CascadeMux I__14401 (
            .O(N__68128),
            .I(\pid_side.un1_pid_prereg_0_18_cascade_ ));
    InMux I__14400 (
            .O(N__68125),
            .I(N__68122));
    LocalMux I__14399 (
            .O(N__68122),
            .I(\pid_side.error_d_reg_prev_esr_RNI0B4M6Z0Z_21 ));
    InMux I__14398 (
            .O(N__68119),
            .I(N__68113));
    InMux I__14397 (
            .O(N__68118),
            .I(N__68113));
    LocalMux I__14396 (
            .O(N__68113),
            .I(\pid_side.un1_pid_prereg_0_7 ));
    CascadeMux I__14395 (
            .O(N__68110),
            .I(N__68107));
    InMux I__14394 (
            .O(N__68107),
            .I(N__68104));
    LocalMux I__14393 (
            .O(N__68104),
            .I(N__68101));
    Span4Mux_h I__14392 (
            .O(N__68101),
            .I(N__68097));
    InMux I__14391 (
            .O(N__68100),
            .I(N__68094));
    Odrv4 I__14390 (
            .O(N__68097),
            .I(\pid_side.un1_pid_prereg_0_9 ));
    LocalMux I__14389 (
            .O(N__68094),
            .I(\pid_side.un1_pid_prereg_0_9 ));
    CascadeMux I__14388 (
            .O(N__68089),
            .I(N__68086));
    InMux I__14387 (
            .O(N__68086),
            .I(N__68079));
    InMux I__14386 (
            .O(N__68085),
            .I(N__68079));
    InMux I__14385 (
            .O(N__68084),
            .I(N__68076));
    LocalMux I__14384 (
            .O(N__68079),
            .I(\pid_side.un1_pid_prereg_0_6 ));
    LocalMux I__14383 (
            .O(N__68076),
            .I(\pid_side.un1_pid_prereg_0_6 ));
    InMux I__14382 (
            .O(N__68071),
            .I(N__68068));
    LocalMux I__14381 (
            .O(N__68068),
            .I(N__68065));
    Span4Mux_v I__14380 (
            .O(N__68065),
            .I(N__68060));
    InMux I__14379 (
            .O(N__68064),
            .I(N__68057));
    InMux I__14378 (
            .O(N__68063),
            .I(N__68054));
    Odrv4 I__14377 (
            .O(N__68060),
            .I(\pid_side.un1_pid_prereg_0_8 ));
    LocalMux I__14376 (
            .O(N__68057),
            .I(\pid_side.un1_pid_prereg_0_8 ));
    LocalMux I__14375 (
            .O(N__68054),
            .I(\pid_side.un1_pid_prereg_0_8 ));
    InMux I__14374 (
            .O(N__68047),
            .I(N__68044));
    LocalMux I__14373 (
            .O(N__68044),
            .I(\pid_side.error_d_reg_prev_esr_RNIGI4KKZ0Z_12 ));
    CascadeMux I__14372 (
            .O(N__68041),
            .I(N__68037));
    InMux I__14371 (
            .O(N__68040),
            .I(N__68033));
    InMux I__14370 (
            .O(N__68037),
            .I(N__68028));
    InMux I__14369 (
            .O(N__68036),
            .I(N__68028));
    LocalMux I__14368 (
            .O(N__68033),
            .I(N__68025));
    LocalMux I__14367 (
            .O(N__68028),
            .I(N__68022));
    Span4Mux_h I__14366 (
            .O(N__68025),
            .I(N__68017));
    Span4Mux_h I__14365 (
            .O(N__68022),
            .I(N__68017));
    Span4Mux_v I__14364 (
            .O(N__68017),
            .I(N__68014));
    Odrv4 I__14363 (
            .O(N__68014),
            .I(\pid_side.error_d_reg_prev_esr_RNI73UC2_0Z0Z_14 ));
    InMux I__14362 (
            .O(N__68011),
            .I(N__68008));
    LocalMux I__14361 (
            .O(N__68008),
            .I(\pid_side.error_d_reg_prev_esr_RNICCO8BZ0Z_12 ));
    InMux I__14360 (
            .O(N__68005),
            .I(N__68002));
    LocalMux I__14359 (
            .O(N__68002),
            .I(\pid_side.error_d_reg_prev_esr_RNIBNLL9Z0Z_18 ));
    InMux I__14358 (
            .O(N__67999),
            .I(N__67996));
    LocalMux I__14357 (
            .O(N__67996),
            .I(N__67993));
    Odrv4 I__14356 (
            .O(N__67993),
            .I(\pid_side.error_d_reg_prev_esr_RNI2BI34Z0Z_21 ));
    InMux I__14355 (
            .O(N__67990),
            .I(N__67986));
    InMux I__14354 (
            .O(N__67989),
            .I(N__67983));
    LocalMux I__14353 (
            .O(N__67986),
            .I(N__67980));
    LocalMux I__14352 (
            .O(N__67983),
            .I(N__67976));
    Span12Mux_s3_v I__14351 (
            .O(N__67980),
            .I(N__67973));
    InMux I__14350 (
            .O(N__67979),
            .I(N__67970));
    Span4Mux_h I__14349 (
            .O(N__67976),
            .I(N__67967));
    Odrv12 I__14348 (
            .O(N__67973),
            .I(\pid_side.error_i_reg_esr_RNIM5PSZ0Z_22 ));
    LocalMux I__14347 (
            .O(N__67970),
            .I(\pid_side.error_i_reg_esr_RNIM5PSZ0Z_22 ));
    Odrv4 I__14346 (
            .O(N__67967),
            .I(\pid_side.error_i_reg_esr_RNIM5PSZ0Z_22 ));
    CascadeMux I__14345 (
            .O(N__67960),
            .I(N__67957));
    InMux I__14344 (
            .O(N__67957),
            .I(N__67953));
    InMux I__14343 (
            .O(N__67956),
            .I(N__67950));
    LocalMux I__14342 (
            .O(N__67953),
            .I(\pid_side.un1_pid_prereg_0_13 ));
    LocalMux I__14341 (
            .O(N__67950),
            .I(\pid_side.un1_pid_prereg_0_13 ));
    InMux I__14340 (
            .O(N__67945),
            .I(N__67940));
    InMux I__14339 (
            .O(N__67944),
            .I(N__67935));
    InMux I__14338 (
            .O(N__67943),
            .I(N__67935));
    LocalMux I__14337 (
            .O(N__67940),
            .I(\pid_side.un1_pid_prereg_0_10 ));
    LocalMux I__14336 (
            .O(N__67935),
            .I(\pid_side.un1_pid_prereg_0_10 ));
    InMux I__14335 (
            .O(N__67930),
            .I(N__67924));
    InMux I__14334 (
            .O(N__67929),
            .I(N__67924));
    LocalMux I__14333 (
            .O(N__67924),
            .I(\pid_side.un1_pid_prereg_0_11 ));
    CascadeMux I__14332 (
            .O(N__67921),
            .I(\pid_side.un1_pid_prereg_0_13_cascade_ ));
    InMux I__14331 (
            .O(N__67918),
            .I(N__67913));
    InMux I__14330 (
            .O(N__67917),
            .I(N__67908));
    InMux I__14329 (
            .O(N__67916),
            .I(N__67908));
    LocalMux I__14328 (
            .O(N__67913),
            .I(\pid_side.un1_pid_prereg_0_12 ));
    LocalMux I__14327 (
            .O(N__67908),
            .I(\pid_side.un1_pid_prereg_0_12 ));
    InMux I__14326 (
            .O(N__67903),
            .I(N__67900));
    LocalMux I__14325 (
            .O(N__67900),
            .I(\pid_side.error_d_reg_prev_esr_RNIR9TU8Z0Z_21 ));
    InMux I__14324 (
            .O(N__67897),
            .I(N__67894));
    LocalMux I__14323 (
            .O(N__67894),
            .I(\pid_side.un1_pid_prereg_0_axb_30 ));
    InMux I__14322 (
            .O(N__67891),
            .I(N__67887));
    InMux I__14321 (
            .O(N__67890),
            .I(N__67884));
    LocalMux I__14320 (
            .O(N__67887),
            .I(N__67881));
    LocalMux I__14319 (
            .O(N__67884),
            .I(N__67877));
    Span4Mux_h I__14318 (
            .O(N__67881),
            .I(N__67874));
    InMux I__14317 (
            .O(N__67880),
            .I(N__67871));
    Odrv12 I__14316 (
            .O(N__67877),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_26_c_RNI0LUS ));
    Odrv4 I__14315 (
            .O(N__67874),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_26_c_RNI0LUS ));
    LocalMux I__14314 (
            .O(N__67871),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_26_c_RNI0LUS ));
    CascadeMux I__14313 (
            .O(N__67864),
            .I(\pid_side.error_d_reg_prev_esr_RNIOUJE2Z0Z_6_cascade_ ));
    CascadeMux I__14312 (
            .O(N__67861),
            .I(\pid_side.un1_pid_prereg_66_0_cascade_ ));
    InMux I__14311 (
            .O(N__67858),
            .I(N__67855));
    LocalMux I__14310 (
            .O(N__67855),
            .I(\pid_side.error_p_reg_esr_RNIRH187Z0Z_5 ));
    InMux I__14309 (
            .O(N__67852),
            .I(N__67847));
    InMux I__14308 (
            .O(N__67851),
            .I(N__67842));
    InMux I__14307 (
            .O(N__67850),
            .I(N__67842));
    LocalMux I__14306 (
            .O(N__67847),
            .I(N__67839));
    LocalMux I__14305 (
            .O(N__67842),
            .I(N__67836));
    Span4Mux_h I__14304 (
            .O(N__67839),
            .I(N__67833));
    Span4Mux_h I__14303 (
            .O(N__67836),
            .I(N__67830));
    Odrv4 I__14302 (
            .O(N__67833),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_5_c_RNIC5QN ));
    Odrv4 I__14301 (
            .O(N__67830),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_5_c_RNIC5QN ));
    InMux I__14300 (
            .O(N__67825),
            .I(N__67822));
    LocalMux I__14299 (
            .O(N__67822),
            .I(\pid_side.error_d_reg_prev_esr_RNIOUJE2Z0Z_6 ));
    CascadeMux I__14298 (
            .O(N__67819),
            .I(N__67816));
    InMux I__14297 (
            .O(N__67816),
            .I(N__67813));
    LocalMux I__14296 (
            .O(N__67813),
            .I(\pid_side.error_p_reg_esr_RNIBABR4Z0Z_5 ));
    InMux I__14295 (
            .O(N__67810),
            .I(N__67806));
    InMux I__14294 (
            .O(N__67809),
            .I(N__67803));
    LocalMux I__14293 (
            .O(N__67806),
            .I(N__67800));
    LocalMux I__14292 (
            .O(N__67803),
            .I(N__67795));
    Span4Mux_v I__14291 (
            .O(N__67800),
            .I(N__67795));
    Odrv4 I__14290 (
            .O(N__67795),
            .I(\pid_side.error_d_reg_prev_esr_RNI8UIO_0Z0Z_15 ));
    InMux I__14289 (
            .O(N__67792),
            .I(N__67786));
    InMux I__14288 (
            .O(N__67791),
            .I(N__67786));
    LocalMux I__14287 (
            .O(N__67786),
            .I(\pid_side.error_d_reg_prevZ0Z_15 ));
    InMux I__14286 (
            .O(N__67783),
            .I(N__67777));
    InMux I__14285 (
            .O(N__67782),
            .I(N__67777));
    LocalMux I__14284 (
            .O(N__67777),
            .I(N__67774));
    Odrv4 I__14283 (
            .O(N__67774),
            .I(\pid_side.error_d_reg_prev_esr_RNI8UIOZ0Z_15 ));
    InMux I__14282 (
            .O(N__67771),
            .I(N__67767));
    InMux I__14281 (
            .O(N__67770),
            .I(N__67764));
    LocalMux I__14280 (
            .O(N__67767),
            .I(N__67759));
    LocalMux I__14279 (
            .O(N__67764),
            .I(N__67759));
    Span4Mux_v I__14278 (
            .O(N__67759),
            .I(N__67756));
    Odrv4 I__14277 (
            .O(N__67756),
            .I(\pid_side.error_d_reg_prev_esr_RNIE4JOZ0Z_17 ));
    InMux I__14276 (
            .O(N__67753),
            .I(N__67750));
    LocalMux I__14275 (
            .O(N__67750),
            .I(N__67746));
    InMux I__14274 (
            .O(N__67749),
            .I(N__67743));
    Span4Mux_v I__14273 (
            .O(N__67746),
            .I(N__67740));
    LocalMux I__14272 (
            .O(N__67743),
            .I(\pid_side.error_d_reg_prevZ0Z_17 ));
    Odrv4 I__14271 (
            .O(N__67740),
            .I(\pid_side.error_d_reg_prevZ0Z_17 ));
    InMux I__14270 (
            .O(N__67735),
            .I(N__67732));
    LocalMux I__14269 (
            .O(N__67732),
            .I(N__67729));
    Sp12to4 I__14268 (
            .O(N__67729),
            .I(N__67726));
    Span12Mux_v I__14267 (
            .O(N__67726),
            .I(N__67723));
    Span12Mux_h I__14266 (
            .O(N__67723),
            .I(N__67720));
    Odrv12 I__14265 (
            .O(N__67720),
            .I(\pid_front.O_0_19 ));
    InMux I__14264 (
            .O(N__67717),
            .I(N__67711));
    InMux I__14263 (
            .O(N__67716),
            .I(N__67711));
    LocalMux I__14262 (
            .O(N__67711),
            .I(N__67708));
    Span4Mux_h I__14261 (
            .O(N__67708),
            .I(N__67705));
    Odrv4 I__14260 (
            .O(N__67705),
            .I(\pid_front.error_p_regZ0Z_15 ));
    CascadeMux I__14259 (
            .O(N__67702),
            .I(N__67699));
    InMux I__14258 (
            .O(N__67699),
            .I(N__67693));
    InMux I__14257 (
            .O(N__67698),
            .I(N__67693));
    LocalMux I__14256 (
            .O(N__67693),
            .I(N__67689));
    InMux I__14255 (
            .O(N__67692),
            .I(N__67681));
    Span4Mux_v I__14254 (
            .O(N__67689),
            .I(N__67678));
    InMux I__14253 (
            .O(N__67688),
            .I(N__67675));
    InMux I__14252 (
            .O(N__67687),
            .I(N__67672));
    InMux I__14251 (
            .O(N__67686),
            .I(N__67669));
    InMux I__14250 (
            .O(N__67685),
            .I(N__67664));
    InMux I__14249 (
            .O(N__67684),
            .I(N__67664));
    LocalMux I__14248 (
            .O(N__67681),
            .I(N__67659));
    Span4Mux_v I__14247 (
            .O(N__67678),
            .I(N__67659));
    LocalMux I__14246 (
            .O(N__67675),
            .I(\pid_front.error_p_regZ0Z_13 ));
    LocalMux I__14245 (
            .O(N__67672),
            .I(\pid_front.error_p_regZ0Z_13 ));
    LocalMux I__14244 (
            .O(N__67669),
            .I(\pid_front.error_p_regZ0Z_13 ));
    LocalMux I__14243 (
            .O(N__67664),
            .I(\pid_front.error_p_regZ0Z_13 ));
    Odrv4 I__14242 (
            .O(N__67659),
            .I(\pid_front.error_p_regZ0Z_13 ));
    InMux I__14241 (
            .O(N__67648),
            .I(N__67642));
    InMux I__14240 (
            .O(N__67647),
            .I(N__67642));
    LocalMux I__14239 (
            .O(N__67642),
            .I(N__67636));
    InMux I__14238 (
            .O(N__67641),
            .I(N__67630));
    InMux I__14237 (
            .O(N__67640),
            .I(N__67627));
    InMux I__14236 (
            .O(N__67639),
            .I(N__67624));
    Span12Mux_h I__14235 (
            .O(N__67636),
            .I(N__67621));
    InMux I__14234 (
            .O(N__67635),
            .I(N__67616));
    InMux I__14233 (
            .O(N__67634),
            .I(N__67616));
    InMux I__14232 (
            .O(N__67633),
            .I(N__67613));
    LocalMux I__14231 (
            .O(N__67630),
            .I(\pid_front.error_d_reg_prevZ0Z_13 ));
    LocalMux I__14230 (
            .O(N__67627),
            .I(\pid_front.error_d_reg_prevZ0Z_13 ));
    LocalMux I__14229 (
            .O(N__67624),
            .I(\pid_front.error_d_reg_prevZ0Z_13 ));
    Odrv12 I__14228 (
            .O(N__67621),
            .I(\pid_front.error_d_reg_prevZ0Z_13 ));
    LocalMux I__14227 (
            .O(N__67616),
            .I(\pid_front.error_d_reg_prevZ0Z_13 ));
    LocalMux I__14226 (
            .O(N__67613),
            .I(\pid_front.error_d_reg_prevZ0Z_13 ));
    InMux I__14225 (
            .O(N__67600),
            .I(N__67596));
    InMux I__14224 (
            .O(N__67599),
            .I(N__67593));
    LocalMux I__14223 (
            .O(N__67596),
            .I(\pid_front.error_d_reg_fastZ0Z_13 ));
    LocalMux I__14222 (
            .O(N__67593),
            .I(\pid_front.error_d_reg_fastZ0Z_13 ));
    CascadeMux I__14221 (
            .O(N__67588),
            .I(N__67584));
    InMux I__14220 (
            .O(N__67587),
            .I(N__67580));
    InMux I__14219 (
            .O(N__67584),
            .I(N__67574));
    InMux I__14218 (
            .O(N__67583),
            .I(N__67574));
    LocalMux I__14217 (
            .O(N__67580),
            .I(N__67571));
    InMux I__14216 (
            .O(N__67579),
            .I(N__67568));
    LocalMux I__14215 (
            .O(N__67574),
            .I(N__67565));
    Odrv4 I__14214 (
            .O(N__67571),
            .I(\pid_front.error_p_regZ0Z_14 ));
    LocalMux I__14213 (
            .O(N__67568),
            .I(\pid_front.error_p_regZ0Z_14 ));
    Odrv4 I__14212 (
            .O(N__67565),
            .I(\pid_front.error_p_regZ0Z_14 ));
    InMux I__14211 (
            .O(N__67558),
            .I(N__67554));
    InMux I__14210 (
            .O(N__67557),
            .I(N__67551));
    LocalMux I__14209 (
            .O(N__67554),
            .I(N__67546));
    LocalMux I__14208 (
            .O(N__67551),
            .I(N__67546));
    Span4Mux_v I__14207 (
            .O(N__67546),
            .I(N__67541));
    InMux I__14206 (
            .O(N__67545),
            .I(N__67536));
    InMux I__14205 (
            .O(N__67544),
            .I(N__67536));
    Odrv4 I__14204 (
            .O(N__67541),
            .I(\pid_front.error_d_reg_prevZ0Z_14 ));
    LocalMux I__14203 (
            .O(N__67536),
            .I(\pid_front.error_d_reg_prevZ0Z_14 ));
    CascadeMux I__14202 (
            .O(N__67531),
            .I(\pid_front.N_2401_0_0_0_cascade_ ));
    InMux I__14201 (
            .O(N__67528),
            .I(N__67525));
    LocalMux I__14200 (
            .O(N__67525),
            .I(N__67522));
    Odrv4 I__14199 (
            .O(N__67522),
            .I(\pid_front.N_4_1_1_1 ));
    CascadeMux I__14198 (
            .O(N__67519),
            .I(\pid_front.g0_2_0_cascade_ ));
    InMux I__14197 (
            .O(N__67516),
            .I(N__67513));
    LocalMux I__14196 (
            .O(N__67513),
            .I(\pid_front.error_p_reg_esr_RNIBIFG6Z0Z_12 ));
    InMux I__14195 (
            .O(N__67510),
            .I(N__67506));
    InMux I__14194 (
            .O(N__67509),
            .I(N__67503));
    LocalMux I__14193 (
            .O(N__67506),
            .I(N__67498));
    LocalMux I__14192 (
            .O(N__67503),
            .I(N__67498));
    Span4Mux_v I__14191 (
            .O(N__67498),
            .I(N__67495));
    Odrv4 I__14190 (
            .O(N__67495),
            .I(\pid_side.error_d_reg_prev_esr_RNISKLO_0Z0Z_20 ));
    InMux I__14189 (
            .O(N__67492),
            .I(N__67486));
    InMux I__14188 (
            .O(N__67491),
            .I(N__67486));
    LocalMux I__14187 (
            .O(N__67486),
            .I(\pid_side.error_d_reg_prevZ0Z_20 ));
    InMux I__14186 (
            .O(N__67483),
            .I(N__67477));
    InMux I__14185 (
            .O(N__67482),
            .I(N__67477));
    LocalMux I__14184 (
            .O(N__67477),
            .I(N__67474));
    Span4Mux_v I__14183 (
            .O(N__67474),
            .I(N__67471));
    Odrv4 I__14182 (
            .O(N__67471),
            .I(\pid_side.error_d_reg_prev_esr_RNISKLOZ0Z_20 ));
    InMux I__14181 (
            .O(N__67468),
            .I(N__67460));
    InMux I__14180 (
            .O(N__67467),
            .I(N__67460));
    InMux I__14179 (
            .O(N__67466),
            .I(N__67455));
    InMux I__14178 (
            .O(N__67465),
            .I(N__67455));
    LocalMux I__14177 (
            .O(N__67460),
            .I(\pid_front.un1_pid_prereg_79 ));
    LocalMux I__14176 (
            .O(N__67455),
            .I(\pid_front.un1_pid_prereg_79 ));
    InMux I__14175 (
            .O(N__67450),
            .I(N__67442));
    InMux I__14174 (
            .O(N__67449),
            .I(N__67442));
    InMux I__14173 (
            .O(N__67448),
            .I(N__67437));
    InMux I__14172 (
            .O(N__67447),
            .I(N__67437));
    LocalMux I__14171 (
            .O(N__67442),
            .I(\pid_front.un1_pid_prereg_135_0 ));
    LocalMux I__14170 (
            .O(N__67437),
            .I(\pid_front.un1_pid_prereg_135_0 ));
    InMux I__14169 (
            .O(N__67432),
            .I(N__67429));
    LocalMux I__14168 (
            .O(N__67429),
            .I(N__67423));
    InMux I__14167 (
            .O(N__67428),
            .I(N__67418));
    InMux I__14166 (
            .O(N__67427),
            .I(N__67418));
    InMux I__14165 (
            .O(N__67426),
            .I(N__67415));
    Odrv4 I__14164 (
            .O(N__67423),
            .I(\pid_front.error_d_reg_prev_fastZ0Z_12 ));
    LocalMux I__14163 (
            .O(N__67418),
            .I(\pid_front.error_d_reg_prev_fastZ0Z_12 ));
    LocalMux I__14162 (
            .O(N__67415),
            .I(\pid_front.error_d_reg_prev_fastZ0Z_12 ));
    InMux I__14161 (
            .O(N__67408),
            .I(N__67405));
    LocalMux I__14160 (
            .O(N__67405),
            .I(N__67402));
    Span12Mux_v I__14159 (
            .O(N__67402),
            .I(N__67399));
    Span12Mux_h I__14158 (
            .O(N__67399),
            .I(N__67396));
    Odrv12 I__14157 (
            .O(N__67396),
            .I(\pid_front.O_0_4 ));
    CascadeMux I__14156 (
            .O(N__67393),
            .I(N__67390));
    InMux I__14155 (
            .O(N__67390),
            .I(N__67386));
    InMux I__14154 (
            .O(N__67389),
            .I(N__67383));
    LocalMux I__14153 (
            .O(N__67386),
            .I(N__67380));
    LocalMux I__14152 (
            .O(N__67383),
            .I(N__67377));
    Span4Mux_h I__14151 (
            .O(N__67380),
            .I(N__67372));
    Span4Mux_h I__14150 (
            .O(N__67377),
            .I(N__67372));
    Odrv4 I__14149 (
            .O(N__67372),
            .I(\pid_front.error_p_regZ0Z_0 ));
    InMux I__14148 (
            .O(N__67369),
            .I(N__67366));
    LocalMux I__14147 (
            .O(N__67366),
            .I(N__67363));
    Span4Mux_v I__14146 (
            .O(N__67363),
            .I(N__67360));
    Sp12to4 I__14145 (
            .O(N__67360),
            .I(N__67357));
    Span12Mux_h I__14144 (
            .O(N__67357),
            .I(N__67354));
    Span12Mux_v I__14143 (
            .O(N__67354),
            .I(N__67351));
    Odrv12 I__14142 (
            .O(N__67351),
            .I(\pid_front.O_0_14 ));
    InMux I__14141 (
            .O(N__67348),
            .I(N__67345));
    LocalMux I__14140 (
            .O(N__67345),
            .I(N__67342));
    Span4Mux_h I__14139 (
            .O(N__67342),
            .I(N__67339));
    Span4Mux_h I__14138 (
            .O(N__67339),
            .I(N__67336));
    Sp12to4 I__14137 (
            .O(N__67336),
            .I(N__67333));
    Span12Mux_v I__14136 (
            .O(N__67333),
            .I(N__67330));
    Odrv12 I__14135 (
            .O(N__67330),
            .I(\pid_front.O_0_15 ));
    InMux I__14134 (
            .O(N__67327),
            .I(N__67324));
    LocalMux I__14133 (
            .O(N__67324),
            .I(N__67321));
    Span4Mux_v I__14132 (
            .O(N__67321),
            .I(N__67318));
    Span4Mux_h I__14131 (
            .O(N__67318),
            .I(N__67315));
    Sp12to4 I__14130 (
            .O(N__67315),
            .I(N__67312));
    Span12Mux_h I__14129 (
            .O(N__67312),
            .I(N__67309));
    Odrv12 I__14128 (
            .O(N__67309),
            .I(\pid_front.O_0_16 ));
    InMux I__14127 (
            .O(N__67306),
            .I(N__67303));
    LocalMux I__14126 (
            .O(N__67303),
            .I(N__67300));
    Span4Mux_h I__14125 (
            .O(N__67300),
            .I(N__67297));
    Sp12to4 I__14124 (
            .O(N__67297),
            .I(N__67294));
    Span12Mux_h I__14123 (
            .O(N__67294),
            .I(N__67291));
    Odrv12 I__14122 (
            .O(N__67291),
            .I(\pid_front.O_0_18 ));
    CascadeMux I__14121 (
            .O(N__67288),
            .I(\pid_front.error_d_reg_fast_esr_RNIQSG63Z0Z_12_cascade_ ));
    InMux I__14120 (
            .O(N__67285),
            .I(N__67279));
    InMux I__14119 (
            .O(N__67284),
            .I(N__67279));
    LocalMux I__14118 (
            .O(N__67279),
            .I(N__67276));
    Span4Mux_v I__14117 (
            .O(N__67276),
            .I(N__67273));
    Odrv4 I__14116 (
            .O(N__67273),
            .I(\pid_front.error_d_reg_esr_RNIETB61Z0Z_13 ));
    InMux I__14115 (
            .O(N__67270),
            .I(N__67264));
    InMux I__14114 (
            .O(N__67269),
            .I(N__67264));
    LocalMux I__14113 (
            .O(N__67264),
            .I(\pid_front.error_p_reg_esr_RNIH0C61_0Z0Z_14 ));
    CascadeMux I__14112 (
            .O(N__67261),
            .I(\pid_front.error_p_reg_esr_RNIK42C6Z0Z_14_cascade_ ));
    CascadeMux I__14111 (
            .O(N__67258),
            .I(\pid_front.un1_pid_prereg_167_0_1_cascade_ ));
    InMux I__14110 (
            .O(N__67255),
            .I(N__67252));
    LocalMux I__14109 (
            .O(N__67252),
            .I(\pid_front.un1_pid_prereg_167_0 ));
    InMux I__14108 (
            .O(N__67249),
            .I(N__67240));
    InMux I__14107 (
            .O(N__67248),
            .I(N__67240));
    InMux I__14106 (
            .O(N__67247),
            .I(N__67240));
    LocalMux I__14105 (
            .O(N__67240),
            .I(N__67237));
    Odrv4 I__14104 (
            .O(N__67237),
            .I(\pid_front.error_d_reg_fast_esr_RNIR9PO_0Z0Z_13 ));
    InMux I__14103 (
            .O(N__67234),
            .I(N__67231));
    LocalMux I__14102 (
            .O(N__67231),
            .I(\pid_front.error_d_reg_fast_esr_RNIQSG63Z0Z_12 ));
    InMux I__14101 (
            .O(N__67228),
            .I(N__67225));
    LocalMux I__14100 (
            .O(N__67225),
            .I(N__67222));
    Span4Mux_h I__14099 (
            .O(N__67222),
            .I(N__67218));
    InMux I__14098 (
            .O(N__67221),
            .I(N__67215));
    Odrv4 I__14097 (
            .O(N__67218),
            .I(\pid_front.error_d_reg_prev_esr_RNIJVGT4Z0Z_12 ));
    LocalMux I__14096 (
            .O(N__67215),
            .I(\pid_front.error_d_reg_prev_esr_RNIJVGT4Z0Z_12 ));
    InMux I__14095 (
            .O(N__67210),
            .I(N__67206));
    InMux I__14094 (
            .O(N__67209),
            .I(N__67203));
    LocalMux I__14093 (
            .O(N__67206),
            .I(N__67198));
    LocalMux I__14092 (
            .O(N__67203),
            .I(N__67198));
    Odrv4 I__14091 (
            .O(N__67198),
            .I(\pid_front.error_p_reg_esr_RNILTVH2Z0Z_12 ));
    InMux I__14090 (
            .O(N__67195),
            .I(N__67191));
    InMux I__14089 (
            .O(N__67194),
            .I(N__67188));
    LocalMux I__14088 (
            .O(N__67191),
            .I(\pid_front.N_2394_i ));
    LocalMux I__14087 (
            .O(N__67188),
            .I(\pid_front.N_2394_i ));
    CascadeMux I__14086 (
            .O(N__67183),
            .I(\pid_front.N_3_i_1_1_cascade_ ));
    InMux I__14085 (
            .O(N__67180),
            .I(N__67177));
    LocalMux I__14084 (
            .O(N__67177),
            .I(N__67174));
    Span4Mux_v I__14083 (
            .O(N__67174),
            .I(N__67171));
    Odrv4 I__14082 (
            .O(N__67171),
            .I(\pid_front.N_3_i_1 ));
    InMux I__14081 (
            .O(N__67168),
            .I(N__67165));
    LocalMux I__14080 (
            .O(N__67165),
            .I(N__67162));
    Span4Mux_v I__14079 (
            .O(N__67162),
            .I(N__67159));
    Odrv4 I__14078 (
            .O(N__67159),
            .I(\pid_front.g0_1_0 ));
    InMux I__14077 (
            .O(N__67156),
            .I(N__67150));
    InMux I__14076 (
            .O(N__67155),
            .I(N__67150));
    LocalMux I__14075 (
            .O(N__67150),
            .I(\pid_front.error_p_reg_esr_RNI8NB61_1Z0Z_11 ));
    CascadeMux I__14074 (
            .O(N__67147),
            .I(N__67144));
    InMux I__14073 (
            .O(N__67144),
            .I(N__67138));
    InMux I__14072 (
            .O(N__67143),
            .I(N__67138));
    LocalMux I__14071 (
            .O(N__67138),
            .I(\pid_front.error_d_reg_prevZ0Z_15 ));
    InMux I__14070 (
            .O(N__67135),
            .I(N__67129));
    InMux I__14069 (
            .O(N__67134),
            .I(N__67129));
    LocalMux I__14068 (
            .O(N__67129),
            .I(N__67126));
    Odrv4 I__14067 (
            .O(N__67126),
            .I(\pid_front.error_p_reg_esr_RNIK3C61Z0Z_15 ));
    InMux I__14066 (
            .O(N__67123),
            .I(N__67120));
    LocalMux I__14065 (
            .O(N__67120),
            .I(\pid_front.error_d_reg_fast_esr_RNI5VGKZ0Z_12 ));
    CascadeMux I__14064 (
            .O(N__67117),
            .I(\pid_front.error_d_reg_fast_esr_RNID6KB1Z0Z_12_cascade_ ));
    InMux I__14063 (
            .O(N__67114),
            .I(N__67108));
    InMux I__14062 (
            .O(N__67113),
            .I(N__67108));
    LocalMux I__14061 (
            .O(N__67108),
            .I(N__67105));
    Span4Mux_v I__14060 (
            .O(N__67105),
            .I(N__67102));
    Odrv4 I__14059 (
            .O(N__67102),
            .I(\pid_front.error_d_reg_prevZ0Z_20 ));
    CascadeMux I__14058 (
            .O(N__67099),
            .I(N__67094));
    CascadeMux I__14057 (
            .O(N__67098),
            .I(N__67085));
    CascadeMux I__14056 (
            .O(N__67097),
            .I(N__67082));
    InMux I__14055 (
            .O(N__67094),
            .I(N__67079));
    CascadeMux I__14054 (
            .O(N__67093),
            .I(N__67075));
    CascadeMux I__14053 (
            .O(N__67092),
            .I(N__67072));
    InMux I__14052 (
            .O(N__67091),
            .I(N__67063));
    InMux I__14051 (
            .O(N__67090),
            .I(N__67063));
    InMux I__14050 (
            .O(N__67089),
            .I(N__67063));
    InMux I__14049 (
            .O(N__67088),
            .I(N__67060));
    InMux I__14048 (
            .O(N__67085),
            .I(N__67055));
    InMux I__14047 (
            .O(N__67082),
            .I(N__67055));
    LocalMux I__14046 (
            .O(N__67079),
            .I(N__67052));
    InMux I__14045 (
            .O(N__67078),
            .I(N__67045));
    InMux I__14044 (
            .O(N__67075),
            .I(N__67045));
    InMux I__14043 (
            .O(N__67072),
            .I(N__67045));
    CascadeMux I__14042 (
            .O(N__67071),
            .I(N__67040));
    CascadeMux I__14041 (
            .O(N__67070),
            .I(N__67036));
    LocalMux I__14040 (
            .O(N__67063),
            .I(N__67027));
    LocalMux I__14039 (
            .O(N__67060),
            .I(N__67027));
    LocalMux I__14038 (
            .O(N__67055),
            .I(N__67027));
    Span4Mux_s3_v I__14037 (
            .O(N__67052),
            .I(N__67027));
    LocalMux I__14036 (
            .O(N__67045),
            .I(N__67024));
    InMux I__14035 (
            .O(N__67044),
            .I(N__67015));
    InMux I__14034 (
            .O(N__67043),
            .I(N__67015));
    InMux I__14033 (
            .O(N__67040),
            .I(N__67015));
    InMux I__14032 (
            .O(N__67039),
            .I(N__67015));
    InMux I__14031 (
            .O(N__67036),
            .I(N__67012));
    Span4Mux_v I__14030 (
            .O(N__67027),
            .I(N__67009));
    Span4Mux_h I__14029 (
            .O(N__67024),
            .I(N__67004));
    LocalMux I__14028 (
            .O(N__67015),
            .I(N__67004));
    LocalMux I__14027 (
            .O(N__67012),
            .I(\pid_front.error_d_reg_prevZ0Z_21 ));
    Odrv4 I__14026 (
            .O(N__67009),
            .I(\pid_front.error_d_reg_prevZ0Z_21 ));
    Odrv4 I__14025 (
            .O(N__67004),
            .I(\pid_front.error_d_reg_prevZ0Z_21 ));
    InMux I__14024 (
            .O(N__66997),
            .I(N__66994));
    LocalMux I__14023 (
            .O(N__66994),
            .I(N__66991));
    Span4Mux_v I__14022 (
            .O(N__66991),
            .I(N__66987));
    InMux I__14021 (
            .O(N__66990),
            .I(N__66984));
    Span4Mux_h I__14020 (
            .O(N__66987),
            .I(N__66981));
    LocalMux I__14019 (
            .O(N__66984),
            .I(N__66978));
    Span4Mux_v I__14018 (
            .O(N__66981),
            .I(N__66974));
    Span4Mux_v I__14017 (
            .O(N__66978),
            .I(N__66971));
    InMux I__14016 (
            .O(N__66977),
            .I(N__66968));
    Odrv4 I__14015 (
            .O(N__66974),
            .I(\pid_front.error_d_regZ0Z_4 ));
    Odrv4 I__14014 (
            .O(N__66971),
            .I(\pid_front.error_d_regZ0Z_4 ));
    LocalMux I__14013 (
            .O(N__66968),
            .I(\pid_front.error_d_regZ0Z_4 ));
    InMux I__14012 (
            .O(N__66961),
            .I(N__66957));
    InMux I__14011 (
            .O(N__66960),
            .I(N__66954));
    LocalMux I__14010 (
            .O(N__66957),
            .I(N__66951));
    LocalMux I__14009 (
            .O(N__66954),
            .I(N__66948));
    Span4Mux_h I__14008 (
            .O(N__66951),
            .I(N__66945));
    Span4Mux_h I__14007 (
            .O(N__66948),
            .I(N__66942));
    Span4Mux_v I__14006 (
            .O(N__66945),
            .I(N__66939));
    Odrv4 I__14005 (
            .O(N__66942),
            .I(\pid_front.error_d_reg_prevZ0Z_4 ));
    Odrv4 I__14004 (
            .O(N__66939),
            .I(\pid_front.error_d_reg_prevZ0Z_4 ));
    InMux I__14003 (
            .O(N__66934),
            .I(N__66931));
    LocalMux I__14002 (
            .O(N__66931),
            .I(N__66928));
    Span4Mux_h I__14001 (
            .O(N__66928),
            .I(N__66925));
    Odrv4 I__14000 (
            .O(N__66925),
            .I(\pid_front.error_p_reg_esr_RNIGL6FZ0Z_8 ));
    InMux I__13999 (
            .O(N__66922),
            .I(N__66915));
    InMux I__13998 (
            .O(N__66921),
            .I(N__66915));
    InMux I__13997 (
            .O(N__66920),
            .I(N__66912));
    LocalMux I__13996 (
            .O(N__66915),
            .I(N__66909));
    LocalMux I__13995 (
            .O(N__66912),
            .I(N__66906));
    Span4Mux_v I__13994 (
            .O(N__66909),
            .I(N__66901));
    Span4Mux_v I__13993 (
            .O(N__66906),
            .I(N__66901));
    Odrv4 I__13992 (
            .O(N__66901),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_8_c_RNI1BPE ));
    InMux I__13991 (
            .O(N__66898),
            .I(N__66889));
    InMux I__13990 (
            .O(N__66897),
            .I(N__66889));
    InMux I__13989 (
            .O(N__66896),
            .I(N__66889));
    LocalMux I__13988 (
            .O(N__66889),
            .I(N__66886));
    Span4Mux_h I__13987 (
            .O(N__66886),
            .I(N__66883));
    Odrv4 I__13986 (
            .O(N__66883),
            .I(\pid_front.N_483 ));
    CascadeMux I__13985 (
            .O(N__66880),
            .I(\pid_front.un1_pid_prereg_0_25_cascade_ ));
    CascadeMux I__13984 (
            .O(N__66877),
            .I(N__66874));
    InMux I__13983 (
            .O(N__66874),
            .I(N__66871));
    LocalMux I__13982 (
            .O(N__66871),
            .I(N__66868));
    Span4Mux_h I__13981 (
            .O(N__66868),
            .I(N__66865));
    Span4Mux_v I__13980 (
            .O(N__66865),
            .I(N__66862));
    Odrv4 I__13979 (
            .O(N__66862),
            .I(\pid_front.error_d_reg_prev_esr_RNIDF6C4Z0Z_21 ));
    InMux I__13978 (
            .O(N__66859),
            .I(N__66856));
    LocalMux I__13977 (
            .O(N__66856),
            .I(N__66853));
    Span4Mux_v I__13976 (
            .O(N__66853),
            .I(N__66850));
    Odrv4 I__13975 (
            .O(N__66850),
            .I(\pid_front.un1_pid_prereg_0_axb_30 ));
    InMux I__13974 (
            .O(N__66847),
            .I(N__66844));
    LocalMux I__13973 (
            .O(N__66844),
            .I(N__66841));
    Span4Mux_v I__13972 (
            .O(N__66841),
            .I(N__66838));
    Odrv4 I__13971 (
            .O(N__66838),
            .I(\pid_front.error_d_reg_prev_esr_RNIR0EO8Z0Z_21 ));
    InMux I__13970 (
            .O(N__66835),
            .I(N__66830));
    InMux I__13969 (
            .O(N__66834),
            .I(N__66825));
    InMux I__13968 (
            .O(N__66833),
            .I(N__66825));
    LocalMux I__13967 (
            .O(N__66830),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_27_c_RNIDSKV ));
    LocalMux I__13966 (
            .O(N__66825),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_27_c_RNIDSKV ));
    CascadeMux I__13965 (
            .O(N__66820),
            .I(N__66816));
    CascadeMux I__13964 (
            .O(N__66819),
            .I(N__66812));
    InMux I__13963 (
            .O(N__66816),
            .I(N__66807));
    InMux I__13962 (
            .O(N__66815),
            .I(N__66807));
    InMux I__13961 (
            .O(N__66812),
            .I(N__66804));
    LocalMux I__13960 (
            .O(N__66807),
            .I(\pid_front.un1_pid_prereg_0_26 ));
    LocalMux I__13959 (
            .O(N__66804),
            .I(\pid_front.un1_pid_prereg_0_26 ));
    InMux I__13958 (
            .O(N__66799),
            .I(N__66795));
    InMux I__13957 (
            .O(N__66798),
            .I(N__66792));
    LocalMux I__13956 (
            .O(N__66795),
            .I(\pid_front.un1_pid_prereg_0_24 ));
    LocalMux I__13955 (
            .O(N__66792),
            .I(\pid_front.un1_pid_prereg_0_24 ));
    InMux I__13954 (
            .O(N__66787),
            .I(N__66784));
    LocalMux I__13953 (
            .O(N__66784),
            .I(N__66781));
    Span4Mux_v I__13952 (
            .O(N__66781),
            .I(N__66778));
    Span4Mux_v I__13951 (
            .O(N__66778),
            .I(N__66774));
    InMux I__13950 (
            .O(N__66777),
            .I(N__66771));
    Odrv4 I__13949 (
            .O(N__66774),
            .I(\pid_front.un1_pid_prereg_0_23 ));
    LocalMux I__13948 (
            .O(N__66771),
            .I(\pid_front.un1_pid_prereg_0_23 ));
    InMux I__13947 (
            .O(N__66766),
            .I(N__66763));
    LocalMux I__13946 (
            .O(N__66763),
            .I(N__66760));
    Span4Mux_v I__13945 (
            .O(N__66760),
            .I(N__66757));
    Span4Mux_v I__13944 (
            .O(N__66757),
            .I(N__66753));
    InMux I__13943 (
            .O(N__66756),
            .I(N__66750));
    Odrv4 I__13942 (
            .O(N__66753),
            .I(\pid_front.un1_pid_prereg_0_22 ));
    LocalMux I__13941 (
            .O(N__66750),
            .I(\pid_front.un1_pid_prereg_0_22 ));
    CascadeMux I__13940 (
            .O(N__66745),
            .I(\pid_front.un1_pid_prereg_0_24_cascade_ ));
    InMux I__13939 (
            .O(N__66742),
            .I(N__66733));
    InMux I__13938 (
            .O(N__66741),
            .I(N__66733));
    InMux I__13937 (
            .O(N__66740),
            .I(N__66726));
    InMux I__13936 (
            .O(N__66739),
            .I(N__66726));
    InMux I__13935 (
            .O(N__66738),
            .I(N__66726));
    LocalMux I__13934 (
            .O(N__66733),
            .I(\pid_front.un1_pid_prereg_0_25 ));
    LocalMux I__13933 (
            .O(N__66726),
            .I(\pid_front.un1_pid_prereg_0_25 ));
    InMux I__13932 (
            .O(N__66721),
            .I(N__66718));
    LocalMux I__13931 (
            .O(N__66718),
            .I(N__66715));
    Span4Mux_v I__13930 (
            .O(N__66715),
            .I(N__66712));
    Odrv4 I__13929 (
            .O(N__66712),
            .I(\pid_front.error_d_reg_prev_esr_RNINPAO8Z0Z_21 ));
    InMux I__13928 (
            .O(N__66709),
            .I(N__66696));
    InMux I__13927 (
            .O(N__66708),
            .I(N__66696));
    InMux I__13926 (
            .O(N__66707),
            .I(N__66696));
    InMux I__13925 (
            .O(N__66706),
            .I(N__66684));
    InMux I__13924 (
            .O(N__66705),
            .I(N__66684));
    InMux I__13923 (
            .O(N__66704),
            .I(N__66684));
    InMux I__13922 (
            .O(N__66703),
            .I(N__66681));
    LocalMux I__13921 (
            .O(N__66696),
            .I(N__66678));
    InMux I__13920 (
            .O(N__66695),
            .I(N__66669));
    InMux I__13919 (
            .O(N__66694),
            .I(N__66669));
    InMux I__13918 (
            .O(N__66693),
            .I(N__66669));
    InMux I__13917 (
            .O(N__66692),
            .I(N__66669));
    CascadeMux I__13916 (
            .O(N__66691),
            .I(N__66664));
    LocalMux I__13915 (
            .O(N__66684),
            .I(N__66658));
    LocalMux I__13914 (
            .O(N__66681),
            .I(N__66651));
    Span4Mux_h I__13913 (
            .O(N__66678),
            .I(N__66651));
    LocalMux I__13912 (
            .O(N__66669),
            .I(N__66651));
    InMux I__13911 (
            .O(N__66668),
            .I(N__66644));
    InMux I__13910 (
            .O(N__66667),
            .I(N__66644));
    InMux I__13909 (
            .O(N__66664),
            .I(N__66644));
    InMux I__13908 (
            .O(N__66663),
            .I(N__66641));
    InMux I__13907 (
            .O(N__66662),
            .I(N__66636));
    InMux I__13906 (
            .O(N__66661),
            .I(N__66636));
    Span4Mux_h I__13905 (
            .O(N__66658),
            .I(N__66631));
    Span4Mux_v I__13904 (
            .O(N__66651),
            .I(N__66631));
    LocalMux I__13903 (
            .O(N__66644),
            .I(\pid_front.error_p_regZ0Z_20 ));
    LocalMux I__13902 (
            .O(N__66641),
            .I(\pid_front.error_p_regZ0Z_20 ));
    LocalMux I__13901 (
            .O(N__66636),
            .I(\pid_front.error_p_regZ0Z_20 ));
    Odrv4 I__13900 (
            .O(N__66631),
            .I(\pid_front.error_p_regZ0Z_20 ));
    InMux I__13899 (
            .O(N__66622),
            .I(N__66618));
    InMux I__13898 (
            .O(N__66621),
            .I(N__66615));
    LocalMux I__13897 (
            .O(N__66618),
            .I(N__66612));
    LocalMux I__13896 (
            .O(N__66615),
            .I(N__66609));
    Span4Mux_h I__13895 (
            .O(N__66612),
            .I(N__66606));
    Span4Mux_v I__13894 (
            .O(N__66609),
            .I(N__66603));
    Odrv4 I__13893 (
            .O(N__66606),
            .I(\pid_front.un1_pid_prereg_370_1 ));
    Odrv4 I__13892 (
            .O(N__66603),
            .I(\pid_front.un1_pid_prereg_370_1 ));
    InMux I__13891 (
            .O(N__66598),
            .I(N__66595));
    LocalMux I__13890 (
            .O(N__66595),
            .I(\pid_front.error_i_acummZ0Z_7 ));
    InMux I__13889 (
            .O(N__66592),
            .I(N__66589));
    LocalMux I__13888 (
            .O(N__66589),
            .I(\pid_front.error_i_acummZ0Z_8 ));
    CascadeMux I__13887 (
            .O(N__66586),
            .I(\pid_front.N_62_i_1_cascade_ ));
    CascadeMux I__13886 (
            .O(N__66583),
            .I(N__66580));
    InMux I__13885 (
            .O(N__66580),
            .I(N__66577));
    LocalMux I__13884 (
            .O(N__66577),
            .I(N__66574));
    Odrv4 I__13883 (
            .O(N__66574),
            .I(\pid_front.error_i_acummZ0Z_3 ));
    InMux I__13882 (
            .O(N__66571),
            .I(N__66568));
    LocalMux I__13881 (
            .O(N__66568),
            .I(\pid_front.N_177 ));
    CascadeMux I__13880 (
            .O(N__66565),
            .I(\pid_front.N_177_cascade_ ));
    CascadeMux I__13879 (
            .O(N__66562),
            .I(\pid_front.N_158_cascade_ ));
    InMux I__13878 (
            .O(N__66559),
            .I(N__66552));
    InMux I__13877 (
            .O(N__66558),
            .I(N__66545));
    InMux I__13876 (
            .O(N__66557),
            .I(N__66545));
    InMux I__13875 (
            .O(N__66556),
            .I(N__66545));
    InMux I__13874 (
            .O(N__66555),
            .I(N__66542));
    LocalMux I__13873 (
            .O(N__66552),
            .I(N__66539));
    LocalMux I__13872 (
            .O(N__66545),
            .I(\pid_front.N_601 ));
    LocalMux I__13871 (
            .O(N__66542),
            .I(\pid_front.N_601 ));
    Odrv12 I__13870 (
            .O(N__66539),
            .I(\pid_front.N_601 ));
    InMux I__13869 (
            .O(N__66532),
            .I(N__66529));
    LocalMux I__13868 (
            .O(N__66529),
            .I(\pid_front.N_208 ));
    InMux I__13867 (
            .O(N__66526),
            .I(N__66520));
    InMux I__13866 (
            .O(N__66525),
            .I(N__66520));
    LocalMux I__13865 (
            .O(N__66520),
            .I(\pid_front.N_181 ));
    InMux I__13864 (
            .O(N__66517),
            .I(N__66514));
    LocalMux I__13863 (
            .O(N__66514),
            .I(\pid_front.error_i_acummZ0Z_1 ));
    InMux I__13862 (
            .O(N__66511),
            .I(N__66505));
    InMux I__13861 (
            .O(N__66510),
            .I(N__66505));
    LocalMux I__13860 (
            .O(N__66505),
            .I(\pid_front.error_i_acumm_13_0_tz_1_0 ));
    InMux I__13859 (
            .O(N__66502),
            .I(N__66499));
    LocalMux I__13858 (
            .O(N__66499),
            .I(\pid_front.error_i_acummZ0Z_2 ));
    CascadeMux I__13857 (
            .O(N__66496),
            .I(N__66493));
    InMux I__13856 (
            .O(N__66493),
            .I(N__66490));
    LocalMux I__13855 (
            .O(N__66490),
            .I(\pid_front.error_i_acummZ0Z_6 ));
    InMux I__13854 (
            .O(N__66487),
            .I(N__66484));
    LocalMux I__13853 (
            .O(N__66484),
            .I(\pid_front.error_i_acummZ0Z_5 ));
    CascadeMux I__13852 (
            .O(N__66481),
            .I(\pid_front.N_633_cascade_ ));
    InMux I__13851 (
            .O(N__66478),
            .I(N__66475));
    LocalMux I__13850 (
            .O(N__66475),
            .I(\pid_front.N_530 ));
    InMux I__13849 (
            .O(N__66472),
            .I(N__66466));
    InMux I__13848 (
            .O(N__66471),
            .I(N__66466));
    LocalMux I__13847 (
            .O(N__66466),
            .I(\pid_front.N_251 ));
    CascadeMux I__13846 (
            .O(N__66463),
            .I(\pid_front.N_251_cascade_ ));
    CascadeMux I__13845 (
            .O(N__66460),
            .I(N__66457));
    InMux I__13844 (
            .O(N__66457),
            .I(N__66454));
    LocalMux I__13843 (
            .O(N__66454),
            .I(\pid_front.error_i_acummZ0Z_4 ));
    CascadeMux I__13842 (
            .O(N__66451),
            .I(pid_side_N_607_cascade_));
    InMux I__13841 (
            .O(N__66448),
            .I(N__66445));
    LocalMux I__13840 (
            .O(N__66445),
            .I(N__66442));
    Span4Mux_h I__13839 (
            .O(N__66442),
            .I(N__66439));
    Span4Mux_h I__13838 (
            .O(N__66439),
            .I(N__66436));
    Odrv4 I__13837 (
            .O(N__66436),
            .I(\pid_front.error_cry_1_0_c_RNINF5AZ0Z3 ));
    CascadeMux I__13836 (
            .O(N__66433),
            .I(N__66430));
    InMux I__13835 (
            .O(N__66430),
            .I(N__66427));
    LocalMux I__13834 (
            .O(N__66427),
            .I(\pid_front.error_i_regZ0Z_2 ));
    CascadeMux I__13833 (
            .O(N__66424),
            .I(N__66421));
    InMux I__13832 (
            .O(N__66421),
            .I(N__66418));
    LocalMux I__13831 (
            .O(N__66418),
            .I(\pid_front.error_i_regZ0Z_1 ));
    CascadeMux I__13830 (
            .O(N__66415),
            .I(pid_front_N_335_cascade_));
    CascadeMux I__13829 (
            .O(N__66412),
            .I(\pid_side.error_i_reg_9_1_rn_sx_16_cascade_ ));
    InMux I__13828 (
            .O(N__66409),
            .I(N__66406));
    LocalMux I__13827 (
            .O(N__66406),
            .I(N__66403));
    Odrv12 I__13826 (
            .O(N__66403),
            .I(\pid_side.error_i_reg_9_1_sn_16 ));
    CascadeMux I__13825 (
            .O(N__66400),
            .I(\pid_side.error_i_reg_9_1_rn_0_16_cascade_ ));
    InMux I__13824 (
            .O(N__66397),
            .I(N__66394));
    LocalMux I__13823 (
            .O(N__66394),
            .I(N__66391));
    Odrv12 I__13822 (
            .O(N__66391),
            .I(\pid_side.error_i_reg_9_1_16 ));
    CascadeMux I__13821 (
            .O(N__66388),
            .I(\pid_front.N_600_cascade_ ));
    InMux I__13820 (
            .O(N__66385),
            .I(N__66382));
    LocalMux I__13819 (
            .O(N__66382),
            .I(N__66379));
    Odrv12 I__13818 (
            .O(N__66379),
            .I(\pid_front.error_i_acumm_preregZ0Z_0 ));
    CascadeMux I__13817 (
            .O(N__66376),
            .I(\pid_front.error_i_acumm_13_0_tz_1_0_cascade_ ));
    InMux I__13816 (
            .O(N__66373),
            .I(N__66370));
    LocalMux I__13815 (
            .O(N__66370),
            .I(N__66367));
    Span4Mux_h I__13814 (
            .O(N__66367),
            .I(N__66363));
    InMux I__13813 (
            .O(N__66366),
            .I(N__66360));
    Odrv4 I__13812 (
            .O(N__66363),
            .I(\pid_front.error_i_acummZ0Z_0 ));
    LocalMux I__13811 (
            .O(N__66360),
            .I(\pid_front.error_i_acummZ0Z_0 ));
    InMux I__13810 (
            .O(N__66355),
            .I(N__66352));
    LocalMux I__13809 (
            .O(N__66352),
            .I(\pid_front.error_i_reg_9_rn_0_27 ));
    InMux I__13808 (
            .O(N__66349),
            .I(N__66346));
    LocalMux I__13807 (
            .O(N__66346),
            .I(\pid_front.N_458 ));
    CascadeMux I__13806 (
            .O(N__66343),
            .I(\pid_front.N_314_cascade_ ));
    InMux I__13805 (
            .O(N__66340),
            .I(N__66337));
    LocalMux I__13804 (
            .O(N__66337),
            .I(N__66334));
    Span4Mux_v I__13803 (
            .O(N__66334),
            .I(N__66329));
    InMux I__13802 (
            .O(N__66333),
            .I(N__66326));
    InMux I__13801 (
            .O(N__66332),
            .I(N__66323));
    Odrv4 I__13800 (
            .O(N__66329),
            .I(\pid_front.N_225 ));
    LocalMux I__13799 (
            .O(N__66326),
            .I(\pid_front.N_225 ));
    LocalMux I__13798 (
            .O(N__66323),
            .I(\pid_front.N_225 ));
    CascadeMux I__13797 (
            .O(N__66316),
            .I(\pid_front.m24_2_03_0_0_cascade_ ));
    InMux I__13796 (
            .O(N__66313),
            .I(N__66310));
    LocalMux I__13795 (
            .O(N__66310),
            .I(\pid_front.m24_2_03_0_1 ));
    CascadeMux I__13794 (
            .O(N__66307),
            .I(\pid_front.m24_2_03_0_cascade_ ));
    CascadeMux I__13793 (
            .O(N__66304),
            .I(N__66301));
    InMux I__13792 (
            .O(N__66301),
            .I(N__66298));
    LocalMux I__13791 (
            .O(N__66298),
            .I(N__66295));
    Span4Mux_v I__13790 (
            .O(N__66295),
            .I(N__66292));
    Odrv4 I__13789 (
            .O(N__66292),
            .I(\pid_front.error_i_regZ0Z_20 ));
    InMux I__13788 (
            .O(N__66289),
            .I(N__66286));
    LocalMux I__13787 (
            .O(N__66286),
            .I(N__66283));
    Span4Mux_h I__13786 (
            .O(N__66283),
            .I(N__66279));
    CascadeMux I__13785 (
            .O(N__66282),
            .I(N__66276));
    Span4Mux_h I__13784 (
            .O(N__66279),
            .I(N__66273));
    InMux I__13783 (
            .O(N__66276),
            .I(N__66270));
    Odrv4 I__13782 (
            .O(N__66273),
            .I(\pid_front.error_i_regZ0Z_0 ));
    LocalMux I__13781 (
            .O(N__66270),
            .I(\pid_front.error_i_regZ0Z_0 ));
    InMux I__13780 (
            .O(N__66265),
            .I(N__66261));
    InMux I__13779 (
            .O(N__66264),
            .I(N__66258));
    LocalMux I__13778 (
            .O(N__66261),
            .I(N__66255));
    LocalMux I__13777 (
            .O(N__66258),
            .I(N__66252));
    Span4Mux_v I__13776 (
            .O(N__66255),
            .I(N__66249));
    Span4Mux_v I__13775 (
            .O(N__66252),
            .I(N__66246));
    Odrv4 I__13774 (
            .O(N__66249),
            .I(\pid_front.error_cry_1_c_RNILQ1FZ0Z2 ));
    Odrv4 I__13773 (
            .O(N__66246),
            .I(\pid_front.error_cry_1_c_RNILQ1FZ0Z2 ));
    InMux I__13772 (
            .O(N__66241),
            .I(N__66238));
    LocalMux I__13771 (
            .O(N__66238),
            .I(\pid_side.N_259 ));
    CascadeMux I__13770 (
            .O(N__66235),
            .I(\pid_side.N_259_cascade_ ));
    InMux I__13769 (
            .O(N__66232),
            .I(N__66229));
    LocalMux I__13768 (
            .O(N__66229),
            .I(N__66226));
    Span4Mux_h I__13767 (
            .O(N__66226),
            .I(N__66223));
    Odrv4 I__13766 (
            .O(N__66223),
            .I(\pid_side.error_i_reg_esr_RNO_2Z0Z_14 ));
    InMux I__13765 (
            .O(N__66220),
            .I(N__66217));
    LocalMux I__13764 (
            .O(N__66217),
            .I(N__66213));
    InMux I__13763 (
            .O(N__66216),
            .I(N__66210));
    Span4Mux_v I__13762 (
            .O(N__66213),
            .I(N__66204));
    LocalMux I__13761 (
            .O(N__66210),
            .I(N__66204));
    InMux I__13760 (
            .O(N__66209),
            .I(N__66201));
    Odrv4 I__13759 (
            .O(N__66204),
            .I(\pid_front.N_156 ));
    LocalMux I__13758 (
            .O(N__66201),
            .I(\pid_front.N_156 ));
    CascadeMux I__13757 (
            .O(N__66196),
            .I(\pid_front.N_163_cascade_ ));
    InMux I__13756 (
            .O(N__66193),
            .I(N__66190));
    LocalMux I__13755 (
            .O(N__66190),
            .I(N__66187));
    Odrv4 I__13754 (
            .O(N__66187),
            .I(\pid_front.N_186 ));
    CascadeMux I__13753 (
            .O(N__66184),
            .I(\pid_front.N_186_cascade_ ));
    InMux I__13752 (
            .O(N__66181),
            .I(N__66178));
    LocalMux I__13751 (
            .O(N__66178),
            .I(\pid_front.N_338 ));
    InMux I__13750 (
            .O(N__66175),
            .I(N__66172));
    LocalMux I__13749 (
            .O(N__66172),
            .I(N__66169));
    Odrv4 I__13748 (
            .O(N__66169),
            .I(\pid_front.N_339 ));
    CascadeMux I__13747 (
            .O(N__66166),
            .I(\pid_front.N_42_i_i_0_cascade_ ));
    InMux I__13746 (
            .O(N__66163),
            .I(N__66160));
    LocalMux I__13745 (
            .O(N__66160),
            .I(\pid_front.error_i_reg_9_sn_27 ));
    InMux I__13744 (
            .O(N__66157),
            .I(N__66151));
    InMux I__13743 (
            .O(N__66156),
            .I(N__66151));
    LocalMux I__13742 (
            .O(N__66151),
            .I(N__66148));
    Sp12to4 I__13741 (
            .O(N__66148),
            .I(N__66145));
    Odrv12 I__13740 (
            .O(N__66145),
            .I(\pid_front.error_i_regZ0Z_27 ));
    CascadeMux I__13739 (
            .O(N__66142),
            .I(\pid_side.N_189_cascade_ ));
    InMux I__13738 (
            .O(N__66139),
            .I(N__66136));
    LocalMux I__13737 (
            .O(N__66136),
            .I(\pid_side.m5_0_03_4_i_i_0 ));
    InMux I__13736 (
            .O(N__66133),
            .I(N__66130));
    LocalMux I__13735 (
            .O(N__66130),
            .I(N__66127));
    Odrv4 I__13734 (
            .O(N__66127),
            .I(\pid_side.N_6 ));
    CascadeMux I__13733 (
            .O(N__66124),
            .I(\pid_side.N_6_cascade_ ));
    CascadeMux I__13732 (
            .O(N__66121),
            .I(\pid_side.error_i_reg_esr_RNO_2Z0Z_16_cascade_ ));
    CascadeMux I__13731 (
            .O(N__66118),
            .I(N__66115));
    InMux I__13730 (
            .O(N__66115),
            .I(N__66112));
    LocalMux I__13729 (
            .O(N__66112),
            .I(N__66109));
    Span4Mux_h I__13728 (
            .O(N__66109),
            .I(N__66106));
    Span4Mux_v I__13727 (
            .O(N__66106),
            .I(N__66103));
    Odrv4 I__13726 (
            .O(N__66103),
            .I(\pid_side.error_i_regZ0Z_16 ));
    InMux I__13725 (
            .O(N__66100),
            .I(N__66097));
    LocalMux I__13724 (
            .O(N__66097),
            .I(\pid_side.m4_2_01 ));
    InMux I__13723 (
            .O(N__66094),
            .I(N__66091));
    LocalMux I__13722 (
            .O(N__66091),
            .I(\pid_side.error_i_reg_esr_RNO_1Z0Z_16 ));
    CascadeMux I__13721 (
            .O(N__66088),
            .I(\pid_side.N_263_cascade_ ));
    InMux I__13720 (
            .O(N__66085),
            .I(N__66082));
    LocalMux I__13719 (
            .O(N__66082),
            .I(\pid_side.error_i_reg_esr_RNO_1Z0Z_14 ));
    InMux I__13718 (
            .O(N__66079),
            .I(N__66076));
    LocalMux I__13717 (
            .O(N__66076),
            .I(\pid_side.m18_2_03_4_o3_1_1 ));
    InMux I__13716 (
            .O(N__66073),
            .I(N__66068));
    InMux I__13715 (
            .O(N__66072),
            .I(N__66065));
    InMux I__13714 (
            .O(N__66071),
            .I(N__66061));
    LocalMux I__13713 (
            .O(N__66068),
            .I(N__66058));
    LocalMux I__13712 (
            .O(N__66065),
            .I(N__66055));
    InMux I__13711 (
            .O(N__66064),
            .I(N__66052));
    LocalMux I__13710 (
            .O(N__66061),
            .I(N__66047));
    Span4Mux_h I__13709 (
            .O(N__66058),
            .I(N__66047));
    Span4Mux_h I__13708 (
            .O(N__66055),
            .I(N__66042));
    LocalMux I__13707 (
            .O(N__66052),
            .I(N__66042));
    Span4Mux_v I__13706 (
            .O(N__66047),
            .I(N__66039));
    Span4Mux_v I__13705 (
            .O(N__66042),
            .I(N__66036));
    Odrv4 I__13704 (
            .O(N__66039),
            .I(\pid_front.N_629 ));
    Odrv4 I__13703 (
            .O(N__66036),
            .I(\pid_front.N_629 ));
    InMux I__13702 (
            .O(N__66031),
            .I(N__66028));
    LocalMux I__13701 (
            .O(N__66028),
            .I(N__66025));
    Span4Mux_h I__13700 (
            .O(N__66025),
            .I(N__66022));
    Span4Mux_v I__13699 (
            .O(N__66022),
            .I(N__66019));
    Odrv4 I__13698 (
            .O(N__66019),
            .I(\pid_side.N_228_0 ));
    CascadeMux I__13697 (
            .O(N__66016),
            .I(\pid_side.m16_2_03_4_0_cascade_ ));
    InMux I__13696 (
            .O(N__66013),
            .I(N__66010));
    LocalMux I__13695 (
            .O(N__66010),
            .I(\pid_side.N_263 ));
    InMux I__13694 (
            .O(N__66007),
            .I(N__66004));
    LocalMux I__13693 (
            .O(N__66004),
            .I(N__66001));
    Span4Mux_v I__13692 (
            .O(N__66001),
            .I(N__65998));
    Odrv4 I__13691 (
            .O(N__65998),
            .I(\pid_front.N_394 ));
    CascadeMux I__13690 (
            .O(N__65995),
            .I(N__65992));
    InMux I__13689 (
            .O(N__65992),
            .I(N__65989));
    LocalMux I__13688 (
            .O(N__65989),
            .I(N__65986));
    Span4Mux_v I__13687 (
            .O(N__65986),
            .I(N__65983));
    Odrv4 I__13686 (
            .O(N__65983),
            .I(\pid_front.error_i_reg_9_rn_1_26 ));
    CascadeMux I__13685 (
            .O(N__65980),
            .I(pid_side_m10_2_03_3_i_0_a2_1_0_cascade_));
    CascadeMux I__13684 (
            .O(N__65977),
            .I(\pid_side.m13_2_03_4_i_0_o2_1_0_cascade_ ));
    InMux I__13683 (
            .O(N__65974),
            .I(N__65971));
    LocalMux I__13682 (
            .O(N__65971),
            .I(\pid_side.error_cry_3_0_c_RNIER8NCZ0 ));
    CascadeMux I__13681 (
            .O(N__65968),
            .I(\pid_side.m18_2_03_4_o3_1_cascade_ ));
    InMux I__13680 (
            .O(N__65965),
            .I(N__65962));
    LocalMux I__13679 (
            .O(N__65962),
            .I(N__65959));
    Odrv4 I__13678 (
            .O(N__65959),
            .I(\pid_side.N_543 ));
    InMux I__13677 (
            .O(N__65956),
            .I(N__65950));
    IoInMux I__13676 (
            .O(N__65955),
            .I(N__65945));
    InMux I__13675 (
            .O(N__65954),
            .I(N__65942));
    InMux I__13674 (
            .O(N__65953),
            .I(N__65938));
    LocalMux I__13673 (
            .O(N__65950),
            .I(N__65933));
    InMux I__13672 (
            .O(N__65949),
            .I(N__65930));
    InMux I__13671 (
            .O(N__65948),
            .I(N__65927));
    LocalMux I__13670 (
            .O(N__65945),
            .I(N__65924));
    LocalMux I__13669 (
            .O(N__65942),
            .I(N__65921));
    InMux I__13668 (
            .O(N__65941),
            .I(N__65918));
    LocalMux I__13667 (
            .O(N__65938),
            .I(N__65914));
    InMux I__13666 (
            .O(N__65937),
            .I(N__65911));
    InMux I__13665 (
            .O(N__65936),
            .I(N__65908));
    Span4Mux_s1_h I__13664 (
            .O(N__65933),
            .I(N__65904));
    LocalMux I__13663 (
            .O(N__65930),
            .I(N__65901));
    LocalMux I__13662 (
            .O(N__65927),
            .I(N__65898));
    IoSpan4Mux I__13661 (
            .O(N__65924),
            .I(N__65895));
    Span4Mux_v I__13660 (
            .O(N__65921),
            .I(N__65890));
    LocalMux I__13659 (
            .O(N__65918),
            .I(N__65890));
    InMux I__13658 (
            .O(N__65917),
            .I(N__65887));
    Span4Mux_v I__13657 (
            .O(N__65914),
            .I(N__65882));
    LocalMux I__13656 (
            .O(N__65911),
            .I(N__65882));
    LocalMux I__13655 (
            .O(N__65908),
            .I(N__65879));
    InMux I__13654 (
            .O(N__65907),
            .I(N__65875));
    Span4Mux_v I__13653 (
            .O(N__65904),
            .I(N__65869));
    Span4Mux_s1_h I__13652 (
            .O(N__65901),
            .I(N__65869));
    Span4Mux_s3_h I__13651 (
            .O(N__65898),
            .I(N__65855));
    IoSpan4Mux I__13650 (
            .O(N__65895),
            .I(N__65851));
    Span4Mux_v I__13649 (
            .O(N__65890),
            .I(N__65846));
    LocalMux I__13648 (
            .O(N__65887),
            .I(N__65846));
    Span4Mux_v I__13647 (
            .O(N__65882),
            .I(N__65842));
    Span4Mux_v I__13646 (
            .O(N__65879),
            .I(N__65839));
    InMux I__13645 (
            .O(N__65878),
            .I(N__65836));
    LocalMux I__13644 (
            .O(N__65875),
            .I(N__65833));
    InMux I__13643 (
            .O(N__65874),
            .I(N__65830));
    Span4Mux_h I__13642 (
            .O(N__65869),
            .I(N__65826));
    InMux I__13641 (
            .O(N__65868),
            .I(N__65823));
    CascadeMux I__13640 (
            .O(N__65867),
            .I(N__65819));
    CascadeMux I__13639 (
            .O(N__65866),
            .I(N__65816));
    CascadeMux I__13638 (
            .O(N__65865),
            .I(N__65813));
    CascadeMux I__13637 (
            .O(N__65864),
            .I(N__65810));
    CascadeMux I__13636 (
            .O(N__65863),
            .I(N__65807));
    CascadeMux I__13635 (
            .O(N__65862),
            .I(N__65804));
    CascadeMux I__13634 (
            .O(N__65861),
            .I(N__65801));
    CascadeMux I__13633 (
            .O(N__65860),
            .I(N__65798));
    CascadeMux I__13632 (
            .O(N__65859),
            .I(N__65795));
    CascadeMux I__13631 (
            .O(N__65858),
            .I(N__65789));
    Span4Mux_h I__13630 (
            .O(N__65855),
            .I(N__65785));
    CascadeMux I__13629 (
            .O(N__65854),
            .I(N__65781));
    Span4Mux_s3_v I__13628 (
            .O(N__65851),
            .I(N__65778));
    Span4Mux_v I__13627 (
            .O(N__65846),
            .I(N__65775));
    InMux I__13626 (
            .O(N__65845),
            .I(N__65772));
    Span4Mux_v I__13625 (
            .O(N__65842),
            .I(N__65765));
    Span4Mux_s1_h I__13624 (
            .O(N__65839),
            .I(N__65765));
    LocalMux I__13623 (
            .O(N__65836),
            .I(N__65765));
    Span4Mux_v I__13622 (
            .O(N__65833),
            .I(N__65762));
    LocalMux I__13621 (
            .O(N__65830),
            .I(N__65759));
    InMux I__13620 (
            .O(N__65829),
            .I(N__65756));
    Span4Mux_h I__13619 (
            .O(N__65826),
            .I(N__65751));
    LocalMux I__13618 (
            .O(N__65823),
            .I(N__65751));
    InMux I__13617 (
            .O(N__65822),
            .I(N__65744));
    InMux I__13616 (
            .O(N__65819),
            .I(N__65744));
    InMux I__13615 (
            .O(N__65816),
            .I(N__65744));
    InMux I__13614 (
            .O(N__65813),
            .I(N__65735));
    InMux I__13613 (
            .O(N__65810),
            .I(N__65735));
    InMux I__13612 (
            .O(N__65807),
            .I(N__65735));
    InMux I__13611 (
            .O(N__65804),
            .I(N__65735));
    InMux I__13610 (
            .O(N__65801),
            .I(N__65728));
    InMux I__13609 (
            .O(N__65798),
            .I(N__65728));
    InMux I__13608 (
            .O(N__65795),
            .I(N__65728));
    CascadeMux I__13607 (
            .O(N__65794),
            .I(N__65725));
    CascadeMux I__13606 (
            .O(N__65793),
            .I(N__65722));
    InMux I__13605 (
            .O(N__65792),
            .I(N__65719));
    InMux I__13604 (
            .O(N__65789),
            .I(N__65716));
    CascadeMux I__13603 (
            .O(N__65788),
            .I(N__65713));
    Span4Mux_v I__13602 (
            .O(N__65785),
            .I(N__65710));
    InMux I__13601 (
            .O(N__65784),
            .I(N__65707));
    InMux I__13600 (
            .O(N__65781),
            .I(N__65701));
    Sp12to4 I__13599 (
            .O(N__65778),
            .I(N__65696));
    Sp12to4 I__13598 (
            .O(N__65775),
            .I(N__65693));
    LocalMux I__13597 (
            .O(N__65772),
            .I(N__65690));
    Span4Mux_v I__13596 (
            .O(N__65765),
            .I(N__65681));
    Span4Mux_h I__13595 (
            .O(N__65762),
            .I(N__65681));
    Span4Mux_s1_h I__13594 (
            .O(N__65759),
            .I(N__65681));
    LocalMux I__13593 (
            .O(N__65756),
            .I(N__65681));
    Span4Mux_v I__13592 (
            .O(N__65751),
            .I(N__65678));
    LocalMux I__13591 (
            .O(N__65744),
            .I(N__65675));
    LocalMux I__13590 (
            .O(N__65735),
            .I(N__65670));
    LocalMux I__13589 (
            .O(N__65728),
            .I(N__65670));
    InMux I__13588 (
            .O(N__65725),
            .I(N__65667));
    InMux I__13587 (
            .O(N__65722),
            .I(N__65664));
    LocalMux I__13586 (
            .O(N__65719),
            .I(N__65661));
    LocalMux I__13585 (
            .O(N__65716),
            .I(N__65658));
    InMux I__13584 (
            .O(N__65713),
            .I(N__65655));
    Span4Mux_h I__13583 (
            .O(N__65710),
            .I(N__65652));
    LocalMux I__13582 (
            .O(N__65707),
            .I(N__65649));
    CascadeMux I__13581 (
            .O(N__65706),
            .I(N__65646));
    CascadeMux I__13580 (
            .O(N__65705),
            .I(N__65642));
    CascadeMux I__13579 (
            .O(N__65704),
            .I(N__65639));
    LocalMux I__13578 (
            .O(N__65701),
            .I(N__65635));
    CascadeMux I__13577 (
            .O(N__65700),
            .I(N__65632));
    CascadeMux I__13576 (
            .O(N__65699),
            .I(N__65629));
    Span12Mux_s10_v I__13575 (
            .O(N__65696),
            .I(N__65623));
    Span12Mux_h I__13574 (
            .O(N__65693),
            .I(N__65623));
    Span4Mux_v I__13573 (
            .O(N__65690),
            .I(N__65618));
    Span4Mux_v I__13572 (
            .O(N__65681),
            .I(N__65618));
    Span4Mux_h I__13571 (
            .O(N__65678),
            .I(N__65615));
    Span4Mux_h I__13570 (
            .O(N__65675),
            .I(N__65612));
    Span4Mux_h I__13569 (
            .O(N__65670),
            .I(N__65605));
    LocalMux I__13568 (
            .O(N__65667),
            .I(N__65605));
    LocalMux I__13567 (
            .O(N__65664),
            .I(N__65605));
    Span4Mux_h I__13566 (
            .O(N__65661),
            .I(N__65602));
    Span4Mux_h I__13565 (
            .O(N__65658),
            .I(N__65597));
    LocalMux I__13564 (
            .O(N__65655),
            .I(N__65597));
    Span4Mux_h I__13563 (
            .O(N__65652),
            .I(N__65592));
    Span4Mux_v I__13562 (
            .O(N__65649),
            .I(N__65592));
    InMux I__13561 (
            .O(N__65646),
            .I(N__65589));
    InMux I__13560 (
            .O(N__65645),
            .I(N__65582));
    InMux I__13559 (
            .O(N__65642),
            .I(N__65582));
    InMux I__13558 (
            .O(N__65639),
            .I(N__65582));
    CascadeMux I__13557 (
            .O(N__65638),
            .I(N__65579));
    Span4Mux_h I__13556 (
            .O(N__65635),
            .I(N__65576));
    InMux I__13555 (
            .O(N__65632),
            .I(N__65571));
    InMux I__13554 (
            .O(N__65629),
            .I(N__65571));
    CascadeMux I__13553 (
            .O(N__65628),
            .I(N__65568));
    Span12Mux_v I__13552 (
            .O(N__65623),
            .I(N__65563));
    Sp12to4 I__13551 (
            .O(N__65618),
            .I(N__65563));
    Span4Mux_v I__13550 (
            .O(N__65615),
            .I(N__65560));
    Span4Mux_h I__13549 (
            .O(N__65612),
            .I(N__65555));
    Span4Mux_v I__13548 (
            .O(N__65605),
            .I(N__65555));
    Span4Mux_v I__13547 (
            .O(N__65602),
            .I(N__65550));
    Span4Mux_v I__13546 (
            .O(N__65597),
            .I(N__65550));
    Span4Mux_v I__13545 (
            .O(N__65592),
            .I(N__65543));
    LocalMux I__13544 (
            .O(N__65589),
            .I(N__65543));
    LocalMux I__13543 (
            .O(N__65582),
            .I(N__65543));
    InMux I__13542 (
            .O(N__65579),
            .I(N__65540));
    Span4Mux_h I__13541 (
            .O(N__65576),
            .I(N__65535));
    LocalMux I__13540 (
            .O(N__65571),
            .I(N__65535));
    InMux I__13539 (
            .O(N__65568),
            .I(N__65532));
    Odrv12 I__13538 (
            .O(N__65563),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__13537 (
            .O(N__65560),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__13536 (
            .O(N__65555),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__13535 (
            .O(N__65550),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__13534 (
            .O(N__65543),
            .I(CONSTANT_ONE_NET));
    LocalMux I__13533 (
            .O(N__65540),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__13532 (
            .O(N__65535),
            .I(CONSTANT_ONE_NET));
    LocalMux I__13531 (
            .O(N__65532),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__13530 (
            .O(N__65515),
            .I(\pid_side.m13_2_03_4_i_0_o2_1_cascade_ ));
    InMux I__13529 (
            .O(N__65512),
            .I(N__65509));
    LocalMux I__13528 (
            .O(N__65509),
            .I(\pid_side.m13_2_03_4_i_3 ));
    CascadeMux I__13527 (
            .O(N__65506),
            .I(\pid_side.m13_2_03_4_i_3_cascade_ ));
    CascadeMux I__13526 (
            .O(N__65503),
            .I(N__65500));
    InMux I__13525 (
            .O(N__65500),
            .I(N__65496));
    InMux I__13524 (
            .O(N__65499),
            .I(N__65493));
    LocalMux I__13523 (
            .O(N__65496),
            .I(N__65490));
    LocalMux I__13522 (
            .O(N__65493),
            .I(\pid_side.error_i_regZ0Z_9 ));
    Odrv4 I__13521 (
            .O(N__65490),
            .I(\pid_side.error_i_regZ0Z_9 ));
    InMux I__13520 (
            .O(N__65485),
            .I(N__65477));
    InMux I__13519 (
            .O(N__65484),
            .I(N__65477));
    InMux I__13518 (
            .O(N__65483),
            .I(N__65472));
    InMux I__13517 (
            .O(N__65482),
            .I(N__65472));
    LocalMux I__13516 (
            .O(N__65477),
            .I(N__65469));
    LocalMux I__13515 (
            .O(N__65472),
            .I(N__65465));
    Span4Mux_v I__13514 (
            .O(N__65469),
            .I(N__65462));
    InMux I__13513 (
            .O(N__65468),
            .I(N__65459));
    Span4Mux_v I__13512 (
            .O(N__65465),
            .I(N__65456));
    Span4Mux_v I__13511 (
            .O(N__65462),
            .I(N__65453));
    LocalMux I__13510 (
            .O(N__65459),
            .I(\pid_side.state_ns_0 ));
    Odrv4 I__13509 (
            .O(N__65456),
            .I(\pid_side.state_ns_0 ));
    Odrv4 I__13508 (
            .O(N__65453),
            .I(\pid_side.state_ns_0 ));
    CascadeMux I__13507 (
            .O(N__65446),
            .I(N__65443));
    InMux I__13506 (
            .O(N__65443),
            .I(N__65439));
    InMux I__13505 (
            .O(N__65442),
            .I(N__65436));
    LocalMux I__13504 (
            .O(N__65439),
            .I(N__65431));
    LocalMux I__13503 (
            .O(N__65436),
            .I(N__65431));
    Odrv4 I__13502 (
            .O(N__65431),
            .I(\pid_side.error_i_regZ0Z_7 ));
    CascadeMux I__13501 (
            .O(N__65428),
            .I(N__65425));
    InMux I__13500 (
            .O(N__65425),
            .I(N__65422));
    LocalMux I__13499 (
            .O(N__65422),
            .I(\pid_side.N_163 ));
    CascadeMux I__13498 (
            .O(N__65419),
            .I(\pid_side.N_163_cascade_ ));
    CascadeMux I__13497 (
            .O(N__65416),
            .I(\pid_side.N_186_cascade_ ));
    InMux I__13496 (
            .O(N__65413),
            .I(N__65410));
    LocalMux I__13495 (
            .O(N__65410),
            .I(\pid_side.error_i_reg_9_sn_27 ));
    InMux I__13494 (
            .O(N__65407),
            .I(N__65404));
    LocalMux I__13493 (
            .O(N__65404),
            .I(N__65399));
    InMux I__13492 (
            .O(N__65403),
            .I(N__65394));
    InMux I__13491 (
            .O(N__65402),
            .I(N__65394));
    Odrv12 I__13490 (
            .O(N__65399),
            .I(\pid_side.error_i_reg_esr_RNI2MSRZ0Z_19 ));
    LocalMux I__13489 (
            .O(N__65394),
            .I(\pid_side.error_i_reg_esr_RNI2MSRZ0Z_19 ));
    CascadeMux I__13488 (
            .O(N__65389),
            .I(\pid_side.un1_pid_prereg_0_7_cascade_ ));
    CascadeMux I__13487 (
            .O(N__65386),
            .I(N__65383));
    InMux I__13486 (
            .O(N__65383),
            .I(N__65380));
    LocalMux I__13485 (
            .O(N__65380),
            .I(N__65377));
    Span4Mux_v I__13484 (
            .O(N__65377),
            .I(N__65374));
    Odrv4 I__13483 (
            .O(N__65374),
            .I(\pid_side.error_d_reg_prev_esr_RNI675Q4Z0Z_17 ));
    CascadeMux I__13482 (
            .O(N__65371),
            .I(\pid_side.N_3_i_1_1_cascade_ ));
    InMux I__13481 (
            .O(N__65368),
            .I(N__65365));
    LocalMux I__13480 (
            .O(N__65365),
            .I(N__65362));
    Span4Mux_h I__13479 (
            .O(N__65362),
            .I(N__65359));
    Odrv4 I__13478 (
            .O(N__65359),
            .I(\pid_side.N_5 ));
    CascadeMux I__13477 (
            .O(N__65356),
            .I(\pid_side.N_3_i_1_cascade_ ));
    CascadeMux I__13476 (
            .O(N__65353),
            .I(\pid_side.error_d_reg_prev_esr_RNIQTGL4Z0Z_12_cascade_ ));
    InMux I__13475 (
            .O(N__65350),
            .I(N__65347));
    LocalMux I__13474 (
            .O(N__65347),
            .I(N__65344));
    Span4Mux_h I__13473 (
            .O(N__65344),
            .I(N__65340));
    InMux I__13472 (
            .O(N__65343),
            .I(N__65337));
    Span4Mux_v I__13471 (
            .O(N__65340),
            .I(N__65334));
    LocalMux I__13470 (
            .O(N__65337),
            .I(N__65331));
    Odrv4 I__13469 (
            .O(N__65334),
            .I(\pid_side.un1_pid_prereg_0_axb_14 ));
    Odrv12 I__13468 (
            .O(N__65331),
            .I(\pid_side.un1_pid_prereg_0_axb_14 ));
    InMux I__13467 (
            .O(N__65326),
            .I(N__65323));
    LocalMux I__13466 (
            .O(N__65323),
            .I(\pid_side.N_5_0 ));
    CascadeMux I__13465 (
            .O(N__65320),
            .I(\pid_side.un1_pid_prereg_79_cascade_ ));
    CascadeMux I__13464 (
            .O(N__65317),
            .I(\pid_side.un1_pid_prereg_0_15_cascade_ ));
    InMux I__13463 (
            .O(N__65314),
            .I(N__65311));
    LocalMux I__13462 (
            .O(N__65311),
            .I(\pid_side.error_d_reg_prev_esr_RNIASUA3Z0Z_21 ));
    InMux I__13461 (
            .O(N__65308),
            .I(N__65305));
    LocalMux I__13460 (
            .O(N__65305),
            .I(N__65300));
    InMux I__13459 (
            .O(N__65304),
            .I(N__65295));
    InMux I__13458 (
            .O(N__65303),
            .I(N__65295));
    Span4Mux_v I__13457 (
            .O(N__65300),
            .I(N__65290));
    LocalMux I__13456 (
            .O(N__65295),
            .I(N__65290));
    Odrv4 I__13455 (
            .O(N__65290),
            .I(\pid_side.error_i_reg_esr_RNIK2OSZ0Z_21 ));
    InMux I__13454 (
            .O(N__65287),
            .I(N__65281));
    InMux I__13453 (
            .O(N__65286),
            .I(N__65281));
    LocalMux I__13452 (
            .O(N__65281),
            .I(\pid_side.un1_pid_prereg_370_1 ));
    InMux I__13451 (
            .O(N__65278),
            .I(N__65274));
    InMux I__13450 (
            .O(N__65277),
            .I(N__65270));
    LocalMux I__13449 (
            .O(N__65274),
            .I(N__65267));
    InMux I__13448 (
            .O(N__65273),
            .I(N__65264));
    LocalMux I__13447 (
            .O(N__65270),
            .I(N__65261));
    Odrv12 I__13446 (
            .O(N__65267),
            .I(\pid_side.error_i_reg_esr_RNIRGURZ0Z_20 ));
    LocalMux I__13445 (
            .O(N__65264),
            .I(\pid_side.error_i_reg_esr_RNIRGURZ0Z_20 ));
    Odrv4 I__13444 (
            .O(N__65261),
            .I(\pid_side.error_i_reg_esr_RNIRGURZ0Z_20 ));
    CascadeMux I__13443 (
            .O(N__65254),
            .I(\pid_side.un1_pid_prereg_0_9_cascade_ ));
    CascadeMux I__13442 (
            .O(N__65251),
            .I(N__65248));
    InMux I__13441 (
            .O(N__65248),
            .I(N__65245));
    LocalMux I__13440 (
            .O(N__65245),
            .I(N__65242));
    Span4Mux_h I__13439 (
            .O(N__65242),
            .I(N__65239));
    Odrv4 I__13438 (
            .O(N__65239),
            .I(\pid_side.error_d_reg_prev_esr_RNIIOAQ4Z0Z_18 ));
    InMux I__13437 (
            .O(N__65236),
            .I(N__65232));
    InMux I__13436 (
            .O(N__65235),
            .I(N__65229));
    LocalMux I__13435 (
            .O(N__65232),
            .I(N__65225));
    LocalMux I__13434 (
            .O(N__65229),
            .I(N__65222));
    InMux I__13433 (
            .O(N__65228),
            .I(N__65219));
    Odrv4 I__13432 (
            .O(N__65225),
            .I(\pid_side.error_i_reg_esr_RNI0JRRZ0Z_18 ));
    Odrv4 I__13431 (
            .O(N__65222),
            .I(\pid_side.error_i_reg_esr_RNI0JRRZ0Z_18 ));
    LocalMux I__13430 (
            .O(N__65219),
            .I(\pid_side.error_i_reg_esr_RNI0JRRZ0Z_18 ));
    CascadeMux I__13429 (
            .O(N__65212),
            .I(N__65209));
    InMux I__13428 (
            .O(N__65209),
            .I(N__65206));
    LocalMux I__13427 (
            .O(N__65206),
            .I(N__65203));
    Span12Mux_s10_v I__13426 (
            .O(N__65203),
            .I(N__65200));
    Odrv12 I__13425 (
            .O(N__65200),
            .I(\pid_side.error_d_reg_prev_esr_RNIME5B3Z0Z_21 ));
    CascadeMux I__13424 (
            .O(N__65197),
            .I(N__65194));
    InMux I__13423 (
            .O(N__65194),
            .I(N__65191));
    LocalMux I__13422 (
            .O(N__65191),
            .I(N__65188));
    Odrv4 I__13421 (
            .O(N__65188),
            .I(\pid_side.pid_preregZ0Z_27 ));
    InMux I__13420 (
            .O(N__65185),
            .I(\pid_side.un1_pid_prereg_0_cry_26 ));
    CascadeMux I__13419 (
            .O(N__65182),
            .I(N__65179));
    InMux I__13418 (
            .O(N__65179),
            .I(N__65176));
    LocalMux I__13417 (
            .O(N__65176),
            .I(N__65173));
    Span4Mux_h I__13416 (
            .O(N__65173),
            .I(N__65170));
    Span4Mux_v I__13415 (
            .O(N__65170),
            .I(N__65167));
    Odrv4 I__13414 (
            .O(N__65167),
            .I(\pid_side.error_d_reg_prev_esr_RNIQK7B3Z0Z_21 ));
    InMux I__13413 (
            .O(N__65164),
            .I(N__65161));
    LocalMux I__13412 (
            .O(N__65161),
            .I(N__65158));
    Odrv4 I__13411 (
            .O(N__65158),
            .I(\pid_side.pid_preregZ0Z_28 ));
    InMux I__13410 (
            .O(N__65155),
            .I(\pid_side.un1_pid_prereg_0_cry_27 ));
    InMux I__13409 (
            .O(N__65152),
            .I(N__65149));
    LocalMux I__13408 (
            .O(N__65149),
            .I(N__65146));
    Span4Mux_h I__13407 (
            .O(N__65146),
            .I(N__65143));
    Odrv4 I__13406 (
            .O(N__65143),
            .I(\pid_side.pid_preregZ0Z_29 ));
    InMux I__13405 (
            .O(N__65140),
            .I(\pid_side.un1_pid_prereg_0_cry_28 ));
    InMux I__13404 (
            .O(N__65137),
            .I(\pid_side.un1_pid_prereg_0_cry_29 ));
    CascadeMux I__13403 (
            .O(N__65134),
            .I(N__65131));
    InMux I__13402 (
            .O(N__65131),
            .I(N__65121));
    InMux I__13401 (
            .O(N__65130),
            .I(N__65121));
    InMux I__13400 (
            .O(N__65129),
            .I(N__65118));
    InMux I__13399 (
            .O(N__65128),
            .I(N__65115));
    InMux I__13398 (
            .O(N__65127),
            .I(N__65112));
    InMux I__13397 (
            .O(N__65126),
            .I(N__65109));
    LocalMux I__13396 (
            .O(N__65121),
            .I(N__65099));
    LocalMux I__13395 (
            .O(N__65118),
            .I(N__65099));
    LocalMux I__13394 (
            .O(N__65115),
            .I(N__65099));
    LocalMux I__13393 (
            .O(N__65112),
            .I(N__65099));
    LocalMux I__13392 (
            .O(N__65109),
            .I(N__65096));
    InMux I__13391 (
            .O(N__65108),
            .I(N__65093));
    Span4Mux_h I__13390 (
            .O(N__65099),
            .I(N__65090));
    Span4Mux_h I__13389 (
            .O(N__65096),
            .I(N__65085));
    LocalMux I__13388 (
            .O(N__65093),
            .I(N__65085));
    Odrv4 I__13387 (
            .O(N__65090),
            .I(\pid_side.pid_preregZ0Z_30 ));
    Odrv4 I__13386 (
            .O(N__65085),
            .I(\pid_side.pid_preregZ0Z_30 ));
    CEMux I__13385 (
            .O(N__65080),
            .I(N__65047));
    CEMux I__13384 (
            .O(N__65079),
            .I(N__65047));
    CEMux I__13383 (
            .O(N__65078),
            .I(N__65047));
    CEMux I__13382 (
            .O(N__65077),
            .I(N__65047));
    CEMux I__13381 (
            .O(N__65076),
            .I(N__65047));
    CEMux I__13380 (
            .O(N__65075),
            .I(N__65047));
    CEMux I__13379 (
            .O(N__65074),
            .I(N__65047));
    CEMux I__13378 (
            .O(N__65073),
            .I(N__65047));
    CEMux I__13377 (
            .O(N__65072),
            .I(N__65047));
    CEMux I__13376 (
            .O(N__65071),
            .I(N__65047));
    CEMux I__13375 (
            .O(N__65070),
            .I(N__65047));
    GlobalMux I__13374 (
            .O(N__65047),
            .I(N__65044));
    gio2CtrlBuf I__13373 (
            .O(N__65044),
            .I(\pid_side.state_0_g_0 ));
    CascadeMux I__13372 (
            .O(N__65041),
            .I(N__65038));
    InMux I__13371 (
            .O(N__65038),
            .I(N__65035));
    LocalMux I__13370 (
            .O(N__65035),
            .I(N__65032));
    Odrv4 I__13369 (
            .O(N__65032),
            .I(\pid_side.error_d_reg_prev_esr_RNIC7HE7Z0Z_21 ));
    CascadeMux I__13368 (
            .O(N__65029),
            .I(\pid_side.un1_pid_prereg_0_11_cascade_ ));
    CascadeMux I__13367 (
            .O(N__65026),
            .I(N__65023));
    InMux I__13366 (
            .O(N__65023),
            .I(N__65020));
    LocalMux I__13365 (
            .O(N__65020),
            .I(N__65017));
    Odrv4 I__13364 (
            .O(N__65017),
            .I(\pid_side.error_d_reg_prev_esr_RNIPUAR4Z0Z_19 ));
    CascadeMux I__13363 (
            .O(N__65014),
            .I(N__65011));
    InMux I__13362 (
            .O(N__65011),
            .I(N__65008));
    LocalMux I__13361 (
            .O(N__65008),
            .I(\pid_side.error_d_reg_prev_esr_RNIE21B3Z0Z_21 ));
    CascadeMux I__13360 (
            .O(N__65005),
            .I(N__65002));
    InMux I__13359 (
            .O(N__65002),
            .I(N__64999));
    LocalMux I__13358 (
            .O(N__64999),
            .I(\pid_side.error_d_reg_prev_esr_RNIMK2Q4Z0Z_16 ));
    CascadeMux I__13357 (
            .O(N__64996),
            .I(N__64993));
    InMux I__13356 (
            .O(N__64993),
            .I(N__64990));
    LocalMux I__13355 (
            .O(N__64990),
            .I(\pid_side.pid_preregZ0Z_19 ));
    InMux I__13354 (
            .O(N__64987),
            .I(\pid_side.un1_pid_prereg_0_cry_18 ));
    InMux I__13353 (
            .O(N__64984),
            .I(N__64981));
    LocalMux I__13352 (
            .O(N__64981),
            .I(\pid_side.pid_preregZ0Z_20 ));
    InMux I__13351 (
            .O(N__64978),
            .I(\pid_side.un1_pid_prereg_0_cry_19 ));
    InMux I__13350 (
            .O(N__64975),
            .I(N__64972));
    LocalMux I__13349 (
            .O(N__64972),
            .I(\pid_side.pid_preregZ0Z_21 ));
    InMux I__13348 (
            .O(N__64969),
            .I(\pid_side.un1_pid_prereg_0_cry_20 ));
    InMux I__13347 (
            .O(N__64966),
            .I(N__64963));
    LocalMux I__13346 (
            .O(N__64963),
            .I(\pid_side.pid_preregZ0Z_22 ));
    InMux I__13345 (
            .O(N__64960),
            .I(\pid_side.un1_pid_prereg_0_cry_21 ));
    CascadeMux I__13344 (
            .O(N__64957),
            .I(N__64954));
    InMux I__13343 (
            .O(N__64954),
            .I(N__64951));
    LocalMux I__13342 (
            .O(N__64951),
            .I(N__64948));
    Odrv4 I__13341 (
            .O(N__64948),
            .I(\pid_side.pid_preregZ0Z_23 ));
    InMux I__13340 (
            .O(N__64945),
            .I(bfn_16_7_0_));
    InMux I__13339 (
            .O(N__64942),
            .I(N__64939));
    LocalMux I__13338 (
            .O(N__64939),
            .I(N__64936));
    Odrv4 I__13337 (
            .O(N__64936),
            .I(\pid_side.pid_preregZ0Z_24 ));
    InMux I__13336 (
            .O(N__64933),
            .I(\pid_side.un1_pid_prereg_0_cry_23 ));
    InMux I__13335 (
            .O(N__64930),
            .I(N__64927));
    LocalMux I__13334 (
            .O(N__64927),
            .I(N__64924));
    Odrv4 I__13333 (
            .O(N__64924),
            .I(\pid_side.pid_preregZ0Z_25 ));
    InMux I__13332 (
            .O(N__64921),
            .I(\pid_side.un1_pid_prereg_0_cry_24 ));
    InMux I__13331 (
            .O(N__64918),
            .I(N__64915));
    LocalMux I__13330 (
            .O(N__64915),
            .I(N__64912));
    Span4Mux_h I__13329 (
            .O(N__64912),
            .I(N__64909));
    Odrv4 I__13328 (
            .O(N__64909),
            .I(\pid_side.error_d_reg_prev_esr_RNI8N8M6Z0Z_21 ));
    InMux I__13327 (
            .O(N__64906),
            .I(N__64903));
    LocalMux I__13326 (
            .O(N__64903),
            .I(N__64900));
    Odrv4 I__13325 (
            .O(N__64900),
            .I(\pid_side.pid_preregZ0Z_26 ));
    InMux I__13324 (
            .O(N__64897),
            .I(\pid_side.un1_pid_prereg_0_cry_25 ));
    InMux I__13323 (
            .O(N__64894),
            .I(N__64891));
    LocalMux I__13322 (
            .O(N__64891),
            .I(N__64888));
    Span4Mux_h I__13321 (
            .O(N__64888),
            .I(N__64885));
    Odrv4 I__13320 (
            .O(N__64885),
            .I(\pid_side.error_d_reg_prev_esr_RNIG3DM6Z0Z_21 ));
    InMux I__13319 (
            .O(N__64882),
            .I(N__64879));
    LocalMux I__13318 (
            .O(N__64879),
            .I(N__64874));
    InMux I__13317 (
            .O(N__64878),
            .I(N__64871));
    CascadeMux I__13316 (
            .O(N__64877),
            .I(N__64868));
    Span4Mux_v I__13315 (
            .O(N__64874),
            .I(N__64865));
    LocalMux I__13314 (
            .O(N__64871),
            .I(N__64862));
    InMux I__13313 (
            .O(N__64868),
            .I(N__64859));
    Span4Mux_h I__13312 (
            .O(N__64865),
            .I(N__64856));
    Span4Mux_v I__13311 (
            .O(N__64862),
            .I(N__64851));
    LocalMux I__13310 (
            .O(N__64859),
            .I(N__64851));
    Odrv4 I__13309 (
            .O(N__64856),
            .I(\pid_side.pid_preregZ0Z_11 ));
    Odrv4 I__13308 (
            .O(N__64851),
            .I(\pid_side.pid_preregZ0Z_11 ));
    InMux I__13307 (
            .O(N__64846),
            .I(\pid_side.un1_pid_prereg_0_cry_10 ));
    CascadeMux I__13306 (
            .O(N__64843),
            .I(N__64840));
    InMux I__13305 (
            .O(N__64840),
            .I(N__64836));
    InMux I__13304 (
            .O(N__64839),
            .I(N__64831));
    LocalMux I__13303 (
            .O(N__64836),
            .I(N__64828));
    InMux I__13302 (
            .O(N__64835),
            .I(N__64823));
    InMux I__13301 (
            .O(N__64834),
            .I(N__64823));
    LocalMux I__13300 (
            .O(N__64831),
            .I(N__64820));
    Span4Mux_h I__13299 (
            .O(N__64828),
            .I(N__64817));
    LocalMux I__13298 (
            .O(N__64823),
            .I(N__64814));
    Odrv12 I__13297 (
            .O(N__64820),
            .I(\pid_side.pid_preregZ0Z_12 ));
    Odrv4 I__13296 (
            .O(N__64817),
            .I(\pid_side.pid_preregZ0Z_12 ));
    Odrv4 I__13295 (
            .O(N__64814),
            .I(\pid_side.pid_preregZ0Z_12 ));
    InMux I__13294 (
            .O(N__64807),
            .I(\pid_side.un1_pid_prereg_0_cry_11 ));
    CascadeMux I__13293 (
            .O(N__64804),
            .I(N__64798));
    InMux I__13292 (
            .O(N__64803),
            .I(N__64792));
    InMux I__13291 (
            .O(N__64802),
            .I(N__64792));
    InMux I__13290 (
            .O(N__64801),
            .I(N__64789));
    InMux I__13289 (
            .O(N__64798),
            .I(N__64784));
    InMux I__13288 (
            .O(N__64797),
            .I(N__64784));
    LocalMux I__13287 (
            .O(N__64792),
            .I(N__64781));
    LocalMux I__13286 (
            .O(N__64789),
            .I(N__64776));
    LocalMux I__13285 (
            .O(N__64784),
            .I(N__64776));
    Odrv12 I__13284 (
            .O(N__64781),
            .I(\pid_side.pid_preregZ0Z_13 ));
    Odrv4 I__13283 (
            .O(N__64776),
            .I(\pid_side.pid_preregZ0Z_13 ));
    InMux I__13282 (
            .O(N__64771),
            .I(\pid_side.un1_pid_prereg_0_cry_12 ));
    InMux I__13281 (
            .O(N__64768),
            .I(N__64765));
    LocalMux I__13280 (
            .O(N__64765),
            .I(N__64762));
    Odrv4 I__13279 (
            .O(N__64762),
            .I(\pid_side.un1_pid_prereg_0_cry_13_THRU_CO ));
    InMux I__13278 (
            .O(N__64759),
            .I(\pid_side.un1_pid_prereg_0_cry_13 ));
    CascadeMux I__13277 (
            .O(N__64756),
            .I(N__64752));
    InMux I__13276 (
            .O(N__64755),
            .I(N__64747));
    InMux I__13275 (
            .O(N__64752),
            .I(N__64747));
    LocalMux I__13274 (
            .O(N__64747),
            .I(N__64744));
    Span4Mux_v I__13273 (
            .O(N__64744),
            .I(N__64740));
    InMux I__13272 (
            .O(N__64743),
            .I(N__64737));
    Span4Mux_h I__13271 (
            .O(N__64740),
            .I(N__64734));
    LocalMux I__13270 (
            .O(N__64737),
            .I(\pid_side.pid_preregZ0Z_15 ));
    Odrv4 I__13269 (
            .O(N__64734),
            .I(\pid_side.pid_preregZ0Z_15 ));
    InMux I__13268 (
            .O(N__64729),
            .I(bfn_16_6_0_));
    CascadeMux I__13267 (
            .O(N__64726),
            .I(N__64723));
    InMux I__13266 (
            .O(N__64723),
            .I(N__64720));
    LocalMux I__13265 (
            .O(N__64720),
            .I(\pid_side.error_d_reg_prev_esr_RNI2SL2GZ0Z_12 ));
    InMux I__13264 (
            .O(N__64717),
            .I(N__64714));
    LocalMux I__13263 (
            .O(N__64714),
            .I(\pid_side.pid_preregZ0Z_16 ));
    InMux I__13262 (
            .O(N__64711),
            .I(\pid_side.un1_pid_prereg_0_cry_15 ));
    InMux I__13261 (
            .O(N__64708),
            .I(N__64705));
    LocalMux I__13260 (
            .O(N__64705),
            .I(\pid_side.error_d_reg_prev_esr_RNISHTJ9Z0Z_14 ));
    CascadeMux I__13259 (
            .O(N__64702),
            .I(N__64699));
    InMux I__13258 (
            .O(N__64699),
            .I(N__64696));
    LocalMux I__13257 (
            .O(N__64696),
            .I(\pid_side.error_d_reg_prev_esr_RNIMFTP4Z0Z_14 ));
    InMux I__13256 (
            .O(N__64693),
            .I(N__64690));
    LocalMux I__13255 (
            .O(N__64690),
            .I(\pid_side.pid_preregZ0Z_17 ));
    InMux I__13254 (
            .O(N__64687),
            .I(\pid_side.un1_pid_prereg_0_cry_16 ));
    InMux I__13253 (
            .O(N__64684),
            .I(N__64681));
    LocalMux I__13252 (
            .O(N__64681),
            .I(\pid_side.error_d_reg_prev_esr_RNISM2K9Z0Z_15 ));
    CascadeMux I__13251 (
            .O(N__64678),
            .I(N__64675));
    InMux I__13250 (
            .O(N__64675),
            .I(N__64672));
    LocalMux I__13249 (
            .O(N__64672),
            .I(\pid_side.error_d_reg_prev_esr_RNI620Q4Z0Z_15 ));
    InMux I__13248 (
            .O(N__64669),
            .I(N__64666));
    LocalMux I__13247 (
            .O(N__64666),
            .I(\pid_side.pid_preregZ0Z_18 ));
    InMux I__13246 (
            .O(N__64663),
            .I(\pid_side.un1_pid_prereg_0_cry_17 ));
    InMux I__13245 (
            .O(N__64660),
            .I(N__64653));
    InMux I__13244 (
            .O(N__64659),
            .I(N__64653));
    CascadeMux I__13243 (
            .O(N__64658),
            .I(N__64650));
    LocalMux I__13242 (
            .O(N__64653),
            .I(N__64647));
    InMux I__13241 (
            .O(N__64650),
            .I(N__64644));
    Odrv4 I__13240 (
            .O(N__64647),
            .I(\pid_side.pid_preregZ0Z_3 ));
    LocalMux I__13239 (
            .O(N__64644),
            .I(\pid_side.pid_preregZ0Z_3 ));
    InMux I__13238 (
            .O(N__64639),
            .I(\pid_side.un1_pid_prereg_0_cry_2 ));
    InMux I__13237 (
            .O(N__64636),
            .I(N__64629));
    InMux I__13236 (
            .O(N__64635),
            .I(N__64629));
    InMux I__13235 (
            .O(N__64634),
            .I(N__64625));
    LocalMux I__13234 (
            .O(N__64629),
            .I(N__64622));
    InMux I__13233 (
            .O(N__64628),
            .I(N__64619));
    LocalMux I__13232 (
            .O(N__64625),
            .I(N__64616));
    Span4Mux_v I__13231 (
            .O(N__64622),
            .I(N__64611));
    LocalMux I__13230 (
            .O(N__64619),
            .I(N__64611));
    Span4Mux_h I__13229 (
            .O(N__64616),
            .I(N__64608));
    Odrv4 I__13228 (
            .O(N__64611),
            .I(\pid_side.pid_preregZ0Z_4 ));
    Odrv4 I__13227 (
            .O(N__64608),
            .I(\pid_side.pid_preregZ0Z_4 ));
    InMux I__13226 (
            .O(N__64603),
            .I(\pid_side.un1_pid_prereg_0_cry_3 ));
    InMux I__13225 (
            .O(N__64600),
            .I(N__64593));
    InMux I__13224 (
            .O(N__64599),
            .I(N__64593));
    InMux I__13223 (
            .O(N__64598),
            .I(N__64589));
    LocalMux I__13222 (
            .O(N__64593),
            .I(N__64586));
    InMux I__13221 (
            .O(N__64592),
            .I(N__64583));
    LocalMux I__13220 (
            .O(N__64589),
            .I(N__64580));
    Span4Mux_v I__13219 (
            .O(N__64586),
            .I(N__64575));
    LocalMux I__13218 (
            .O(N__64583),
            .I(N__64575));
    Span4Mux_h I__13217 (
            .O(N__64580),
            .I(N__64572));
    Odrv4 I__13216 (
            .O(N__64575),
            .I(\pid_side.pid_preregZ0Z_5 ));
    Odrv4 I__13215 (
            .O(N__64572),
            .I(\pid_side.pid_preregZ0Z_5 ));
    InMux I__13214 (
            .O(N__64567),
            .I(\pid_side.un1_pid_prereg_0_cry_4 ));
    CascadeMux I__13213 (
            .O(N__64564),
            .I(N__64560));
    InMux I__13212 (
            .O(N__64563),
            .I(N__64556));
    InMux I__13211 (
            .O(N__64560),
            .I(N__64553));
    InMux I__13210 (
            .O(N__64559),
            .I(N__64550));
    LocalMux I__13209 (
            .O(N__64556),
            .I(N__64547));
    LocalMux I__13208 (
            .O(N__64553),
            .I(N__64544));
    LocalMux I__13207 (
            .O(N__64550),
            .I(N__64541));
    Span4Mux_h I__13206 (
            .O(N__64547),
            .I(N__64538));
    Span4Mux_h I__13205 (
            .O(N__64544),
            .I(N__64533));
    Span4Mux_h I__13204 (
            .O(N__64541),
            .I(N__64533));
    Odrv4 I__13203 (
            .O(N__64538),
            .I(\pid_side.pid_preregZ0Z_6 ));
    Odrv4 I__13202 (
            .O(N__64533),
            .I(\pid_side.pid_preregZ0Z_6 ));
    InMux I__13201 (
            .O(N__64528),
            .I(\pid_side.un1_pid_prereg_0_cry_5 ));
    CascadeMux I__13200 (
            .O(N__64525),
            .I(N__64520));
    CascadeMux I__13199 (
            .O(N__64524),
            .I(N__64517));
    InMux I__13198 (
            .O(N__64523),
            .I(N__64514));
    InMux I__13197 (
            .O(N__64520),
            .I(N__64511));
    InMux I__13196 (
            .O(N__64517),
            .I(N__64508));
    LocalMux I__13195 (
            .O(N__64514),
            .I(N__64505));
    LocalMux I__13194 (
            .O(N__64511),
            .I(N__64502));
    LocalMux I__13193 (
            .O(N__64508),
            .I(N__64499));
    Span4Mux_h I__13192 (
            .O(N__64505),
            .I(N__64494));
    Span4Mux_h I__13191 (
            .O(N__64502),
            .I(N__64494));
    Odrv4 I__13190 (
            .O(N__64499),
            .I(\pid_side.pid_preregZ0Z_7 ));
    Odrv4 I__13189 (
            .O(N__64494),
            .I(\pid_side.pid_preregZ0Z_7 ));
    InMux I__13188 (
            .O(N__64489),
            .I(bfn_16_5_0_));
    CascadeMux I__13187 (
            .O(N__64486),
            .I(N__64483));
    InMux I__13186 (
            .O(N__64483),
            .I(N__64480));
    LocalMux I__13185 (
            .O(N__64480),
            .I(N__64475));
    InMux I__13184 (
            .O(N__64479),
            .I(N__64470));
    InMux I__13183 (
            .O(N__64478),
            .I(N__64470));
    Span4Mux_h I__13182 (
            .O(N__64475),
            .I(N__64467));
    LocalMux I__13181 (
            .O(N__64470),
            .I(N__64464));
    Odrv4 I__13180 (
            .O(N__64467),
            .I(\pid_side.pid_preregZ0Z_8 ));
    Odrv4 I__13179 (
            .O(N__64464),
            .I(\pid_side.pid_preregZ0Z_8 ));
    InMux I__13178 (
            .O(N__64459),
            .I(\pid_side.un1_pid_prereg_0_cry_7 ));
    InMux I__13177 (
            .O(N__64456),
            .I(N__64453));
    LocalMux I__13176 (
            .O(N__64453),
            .I(N__64448));
    InMux I__13175 (
            .O(N__64452),
            .I(N__64443));
    InMux I__13174 (
            .O(N__64451),
            .I(N__64443));
    Span4Mux_v I__13173 (
            .O(N__64448),
            .I(N__64438));
    LocalMux I__13172 (
            .O(N__64443),
            .I(N__64438));
    Odrv4 I__13171 (
            .O(N__64438),
            .I(\pid_side.pid_preregZ0Z_9 ));
    InMux I__13170 (
            .O(N__64435),
            .I(\pid_side.un1_pid_prereg_0_cry_8 ));
    CascadeMux I__13169 (
            .O(N__64432),
            .I(N__64429));
    InMux I__13168 (
            .O(N__64429),
            .I(N__64426));
    LocalMux I__13167 (
            .O(N__64426),
            .I(N__64421));
    InMux I__13166 (
            .O(N__64425),
            .I(N__64416));
    InMux I__13165 (
            .O(N__64424),
            .I(N__64416));
    Span4Mux_v I__13164 (
            .O(N__64421),
            .I(N__64411));
    LocalMux I__13163 (
            .O(N__64416),
            .I(N__64411));
    Odrv4 I__13162 (
            .O(N__64411),
            .I(\pid_side.pid_preregZ0Z_10 ));
    InMux I__13161 (
            .O(N__64408),
            .I(\pid_side.un1_pid_prereg_0_cry_9 ));
    InMux I__13160 (
            .O(N__64405),
            .I(N__64401));
    InMux I__13159 (
            .O(N__64404),
            .I(N__64398));
    LocalMux I__13158 (
            .O(N__64401),
            .I(N__64393));
    LocalMux I__13157 (
            .O(N__64398),
            .I(N__64390));
    InMux I__13156 (
            .O(N__64397),
            .I(N__64385));
    InMux I__13155 (
            .O(N__64396),
            .I(N__64385));
    Sp12to4 I__13154 (
            .O(N__64393),
            .I(N__64382));
    Span4Mux_s3_v I__13153 (
            .O(N__64390),
            .I(N__64377));
    LocalMux I__13152 (
            .O(N__64385),
            .I(N__64377));
    Span12Mux_s10_v I__13151 (
            .O(N__64382),
            .I(N__64374));
    Span4Mux_v I__13150 (
            .O(N__64377),
            .I(N__64371));
    Odrv12 I__13149 (
            .O(N__64374),
            .I(\pid_front.error_i_reg_esr_RNI29BUZ0Z_13 ));
    Odrv4 I__13148 (
            .O(N__64371),
            .I(\pid_front.error_i_reg_esr_RNI29BUZ0Z_13 ));
    CascadeMux I__13147 (
            .O(N__64366),
            .I(\pid_front.g1_3_cascade_ ));
    InMux I__13146 (
            .O(N__64363),
            .I(N__64357));
    InMux I__13145 (
            .O(N__64362),
            .I(N__64357));
    LocalMux I__13144 (
            .O(N__64357),
            .I(N__64354));
    Span4Mux_v I__13143 (
            .O(N__64354),
            .I(N__64349));
    InMux I__13142 (
            .O(N__64353),
            .I(N__64343));
    InMux I__13141 (
            .O(N__64352),
            .I(N__64340));
    Span4Mux_v I__13140 (
            .O(N__64349),
            .I(N__64337));
    InMux I__13139 (
            .O(N__64348),
            .I(N__64330));
    InMux I__13138 (
            .O(N__64347),
            .I(N__64330));
    InMux I__13137 (
            .O(N__64346),
            .I(N__64330));
    LocalMux I__13136 (
            .O(N__64343),
            .I(\pid_front.error_d_regZ0Z_13 ));
    LocalMux I__13135 (
            .O(N__64340),
            .I(\pid_front.error_d_regZ0Z_13 ));
    Odrv4 I__13134 (
            .O(N__64337),
            .I(\pid_front.error_d_regZ0Z_13 ));
    LocalMux I__13133 (
            .O(N__64330),
            .I(\pid_front.error_d_regZ0Z_13 ));
    CascadeMux I__13132 (
            .O(N__64321),
            .I(\pid_front.N_2401_0_cascade_ ));
    InMux I__13131 (
            .O(N__64318),
            .I(N__64315));
    LocalMux I__13130 (
            .O(N__64315),
            .I(N__64312));
    Odrv4 I__13129 (
            .O(N__64312),
            .I(\pid_front.g0_2 ));
    InMux I__13128 (
            .O(N__64309),
            .I(N__64306));
    LocalMux I__13127 (
            .O(N__64306),
            .I(N__64303));
    Odrv4 I__13126 (
            .O(N__64303),
            .I(\pid_side.source_pid10lt4_0 ));
    InMux I__13125 (
            .O(N__64300),
            .I(N__64297));
    LocalMux I__13124 (
            .O(N__64297),
            .I(N__64293));
    InMux I__13123 (
            .O(N__64296),
            .I(N__64290));
    Span4Mux_v I__13122 (
            .O(N__64293),
            .I(N__64284));
    LocalMux I__13121 (
            .O(N__64290),
            .I(N__64284));
    InMux I__13120 (
            .O(N__64289),
            .I(N__64281));
    Odrv4 I__13119 (
            .O(N__64284),
            .I(\pid_side.pid_preregZ0Z_0 ));
    LocalMux I__13118 (
            .O(N__64281),
            .I(\pid_side.pid_preregZ0Z_0 ));
    InMux I__13117 (
            .O(N__64276),
            .I(\pid_side.un1_pid_prereg_0_cry_0_c_THRU_CO ));
    InMux I__13116 (
            .O(N__64273),
            .I(N__64267));
    InMux I__13115 (
            .O(N__64272),
            .I(N__64267));
    LocalMux I__13114 (
            .O(N__64267),
            .I(N__64263));
    InMux I__13113 (
            .O(N__64266),
            .I(N__64260));
    Odrv4 I__13112 (
            .O(N__64263),
            .I(\pid_side.pid_preregZ0Z_1 ));
    LocalMux I__13111 (
            .O(N__64260),
            .I(\pid_side.pid_preregZ0Z_1 ));
    InMux I__13110 (
            .O(N__64255),
            .I(\pid_side.un1_pid_prereg_0_cry_0 ));
    InMux I__13109 (
            .O(N__64252),
            .I(N__64246));
    InMux I__13108 (
            .O(N__64251),
            .I(N__64246));
    LocalMux I__13107 (
            .O(N__64246),
            .I(N__64242));
    InMux I__13106 (
            .O(N__64245),
            .I(N__64239));
    Odrv4 I__13105 (
            .O(N__64242),
            .I(\pid_side.pid_preregZ0Z_2 ));
    LocalMux I__13104 (
            .O(N__64239),
            .I(\pid_side.pid_preregZ0Z_2 ));
    InMux I__13103 (
            .O(N__64234),
            .I(\pid_side.un1_pid_prereg_0_cry_1 ));
    InMux I__13102 (
            .O(N__64231),
            .I(N__64225));
    InMux I__13101 (
            .O(N__64230),
            .I(N__64225));
    LocalMux I__13100 (
            .O(N__64225),
            .I(N__64222));
    Span4Mux_h I__13099 (
            .O(N__64222),
            .I(N__64219));
    Span4Mux_h I__13098 (
            .O(N__64219),
            .I(N__64216));
    Span4Mux_h I__13097 (
            .O(N__64216),
            .I(N__64213));
    Odrv4 I__13096 (
            .O(N__64213),
            .I(\pid_front.O_16 ));
    InMux I__13095 (
            .O(N__64210),
            .I(N__64207));
    LocalMux I__13094 (
            .O(N__64207),
            .I(N__64204));
    Span4Mux_h I__13093 (
            .O(N__64204),
            .I(N__64201));
    Sp12to4 I__13092 (
            .O(N__64201),
            .I(N__64198));
    Span12Mux_s4_v I__13091 (
            .O(N__64198),
            .I(N__64195));
    Span12Mux_h I__13090 (
            .O(N__64195),
            .I(N__64192));
    Odrv12 I__13089 (
            .O(N__64192),
            .I(\pid_front.O_0_17 ));
    InMux I__13088 (
            .O(N__64189),
            .I(N__64183));
    InMux I__13087 (
            .O(N__64188),
            .I(N__64183));
    LocalMux I__13086 (
            .O(N__64183),
            .I(N__64180));
    Span4Mux_h I__13085 (
            .O(N__64180),
            .I(N__64177));
    Odrv4 I__13084 (
            .O(N__64177),
            .I(\pid_front.error_d_reg_prev_esr_RNI8QE61_0Z0Z_20 ));
    InMux I__13083 (
            .O(N__64174),
            .I(N__64170));
    InMux I__13082 (
            .O(N__64173),
            .I(N__64167));
    LocalMux I__13081 (
            .O(N__64170),
            .I(N__64164));
    LocalMux I__13080 (
            .O(N__64167),
            .I(N__64161));
    Span4Mux_v I__13079 (
            .O(N__64164),
            .I(N__64158));
    Span4Mux_h I__13078 (
            .O(N__64161),
            .I(N__64155));
    Odrv4 I__13077 (
            .O(N__64158),
            .I(\pid_front.error_d_reg_prev_esr_RNI8QE61Z0Z_20 ));
    Odrv4 I__13076 (
            .O(N__64155),
            .I(\pid_front.error_d_reg_prev_esr_RNI8QE61Z0Z_20 ));
    InMux I__13075 (
            .O(N__64150),
            .I(N__64147));
    LocalMux I__13074 (
            .O(N__64147),
            .I(N__64144));
    Span4Mux_v I__13073 (
            .O(N__64144),
            .I(N__64141));
    Span4Mux_h I__13072 (
            .O(N__64141),
            .I(N__64138));
    Sp12to4 I__13071 (
            .O(N__64138),
            .I(N__64135));
    Span12Mux_h I__13070 (
            .O(N__64135),
            .I(N__64132));
    Odrv12 I__13069 (
            .O(N__64132),
            .I(\pid_front.O_0_24 ));
    CascadeMux I__13068 (
            .O(N__64129),
            .I(\pid_front.error_d_reg_fast_esr_RNISQ181Z0Z_12_cascade_ ));
    InMux I__13067 (
            .O(N__64126),
            .I(N__64123));
    LocalMux I__13066 (
            .O(N__64123),
            .I(\pid_front.error_d_reg_esr_RNIETB61_3Z0Z_13 ));
    InMux I__13065 (
            .O(N__64120),
            .I(N__64117));
    LocalMux I__13064 (
            .O(N__64117),
            .I(N__64114));
    Span4Mux_v I__13063 (
            .O(N__64114),
            .I(N__64111));
    Odrv4 I__13062 (
            .O(N__64111),
            .I(\pid_front.g1_2_1 ));
    CascadeMux I__13061 (
            .O(N__64108),
            .I(\pid_front.g0_3_2_cascade_ ));
    InMux I__13060 (
            .O(N__64105),
            .I(N__64099));
    InMux I__13059 (
            .O(N__64104),
            .I(N__64099));
    LocalMux I__13058 (
            .O(N__64099),
            .I(\pid_front.error_i_acumm_preregZ0Z_13 ));
    InMux I__13057 (
            .O(N__64096),
            .I(N__64090));
    InMux I__13056 (
            .O(N__64095),
            .I(N__64090));
    LocalMux I__13055 (
            .O(N__64090),
            .I(\pid_front.error_i_acumm_preregZ0Z_18 ));
    InMux I__13054 (
            .O(N__64087),
            .I(N__64082));
    InMux I__13053 (
            .O(N__64086),
            .I(N__64079));
    InMux I__13052 (
            .O(N__64085),
            .I(N__64076));
    LocalMux I__13051 (
            .O(N__64082),
            .I(N__64069));
    LocalMux I__13050 (
            .O(N__64079),
            .I(N__64069));
    LocalMux I__13049 (
            .O(N__64076),
            .I(N__64069));
    Span4Mux_v I__13048 (
            .O(N__64069),
            .I(N__64066));
    Odrv4 I__13047 (
            .O(N__64066),
            .I(\pid_front.error_i_reg_esr_RNI8KHVZ0Z_25 ));
    InMux I__13046 (
            .O(N__64063),
            .I(N__64057));
    InMux I__13045 (
            .O(N__64062),
            .I(N__64057));
    LocalMux I__13044 (
            .O(N__64057),
            .I(\pid_front.error_i_acumm_preregZ0Z_25 ));
    InMux I__13043 (
            .O(N__64054),
            .I(N__64049));
    InMux I__13042 (
            .O(N__64053),
            .I(N__64046));
    InMux I__13041 (
            .O(N__64052),
            .I(N__64043));
    LocalMux I__13040 (
            .O(N__64049),
            .I(N__64036));
    LocalMux I__13039 (
            .O(N__64046),
            .I(N__64036));
    LocalMux I__13038 (
            .O(N__64043),
            .I(N__64036));
    Span4Mux_v I__13037 (
            .O(N__64036),
            .I(N__64033));
    Odrv4 I__13036 (
            .O(N__64033),
            .I(\pid_front.error_i_reg_esr_RNIANIVZ0Z_26 ));
    CascadeMux I__13035 (
            .O(N__64030),
            .I(N__64026));
    CascadeMux I__13034 (
            .O(N__64029),
            .I(N__64023));
    InMux I__13033 (
            .O(N__64026),
            .I(N__64018));
    InMux I__13032 (
            .O(N__64023),
            .I(N__64018));
    LocalMux I__13031 (
            .O(N__64018),
            .I(\pid_front.error_i_acumm_preregZ0Z_26 ));
    InMux I__13030 (
            .O(N__64015),
            .I(N__64011));
    InMux I__13029 (
            .O(N__64014),
            .I(N__64008));
    LocalMux I__13028 (
            .O(N__64011),
            .I(N__64005));
    LocalMux I__13027 (
            .O(N__64008),
            .I(N__64002));
    Span4Mux_h I__13026 (
            .O(N__64005),
            .I(N__63999));
    Odrv4 I__13025 (
            .O(N__64002),
            .I(\pid_front.error_d_reg_prev_esr_RNIL8SR5Z0Z_12 ));
    Odrv4 I__13024 (
            .O(N__63999),
            .I(\pid_front.error_d_reg_prev_esr_RNIL8SR5Z0Z_12 ));
    InMux I__13023 (
            .O(N__63994),
            .I(N__63990));
    InMux I__13022 (
            .O(N__63993),
            .I(N__63987));
    LocalMux I__13021 (
            .O(N__63990),
            .I(N__63984));
    LocalMux I__13020 (
            .O(N__63987),
            .I(N__63981));
    Odrv12 I__13019 (
            .O(N__63984),
            .I(\pid_front.error_p_reg_esr_RNITCC61_0Z0Z_18 ));
    Odrv4 I__13018 (
            .O(N__63981),
            .I(\pid_front.error_p_reg_esr_RNITCC61_0Z0Z_18 ));
    InMux I__13017 (
            .O(N__63976),
            .I(N__63972));
    InMux I__13016 (
            .O(N__63975),
            .I(N__63969));
    LocalMux I__13015 (
            .O(N__63972),
            .I(N__63964));
    LocalMux I__13014 (
            .O(N__63969),
            .I(N__63964));
    Odrv4 I__13013 (
            .O(N__63964),
            .I(\pid_front.error_p_reg_esr_RNIQ9C61Z0Z_17 ));
    InMux I__13012 (
            .O(N__63961),
            .I(N__63956));
    InMux I__13011 (
            .O(N__63960),
            .I(N__63951));
    InMux I__13010 (
            .O(N__63959),
            .I(N__63951));
    LocalMux I__13009 (
            .O(N__63956),
            .I(N__63946));
    LocalMux I__13008 (
            .O(N__63951),
            .I(N__63946));
    Odrv12 I__13007 (
            .O(N__63946),
            .I(\pid_front.error_i_reg_esr_RNICOGUZ0Z_18 ));
    InMux I__13006 (
            .O(N__63943),
            .I(N__63934));
    InMux I__13005 (
            .O(N__63942),
            .I(N__63934));
    InMux I__13004 (
            .O(N__63941),
            .I(N__63934));
    LocalMux I__13003 (
            .O(N__63934),
            .I(\pid_front.un1_pid_prereg_0_5 ));
    CascadeMux I__13002 (
            .O(N__63931),
            .I(\pid_front.error_d_reg_prev_esr_RNI5JRF4Z0Z_10_cascade_ ));
    CascadeMux I__13001 (
            .O(N__63928),
            .I(N__63925));
    InMux I__13000 (
            .O(N__63925),
            .I(N__63922));
    LocalMux I__12999 (
            .O(N__63922),
            .I(N__63919));
    Odrv4 I__12998 (
            .O(N__63919),
            .I(\pid_front.error_p_reg_esr_RNIEU1SDZ0Z_12 ));
    CascadeMux I__12997 (
            .O(N__63916),
            .I(N__63913));
    InMux I__12996 (
            .O(N__63913),
            .I(N__63910));
    LocalMux I__12995 (
            .O(N__63910),
            .I(N__63907));
    Span4Mux_h I__12994 (
            .O(N__63907),
            .I(N__63904));
    Odrv4 I__12993 (
            .O(N__63904),
            .I(\pid_front.error_p_reg_esr_RNIUKHM6Z0Z_16 ));
    CascadeMux I__12992 (
            .O(N__63901),
            .I(\pid_front.un1_pid_prereg_0_6_cascade_ ));
    InMux I__12991 (
            .O(N__63898),
            .I(N__63895));
    LocalMux I__12990 (
            .O(N__63895),
            .I(N__63892));
    Odrv12 I__12989 (
            .O(N__63892),
            .I(\pid_front.error_p_reg_esr_RNICS5DDZ0Z_16 ));
    InMux I__12988 (
            .O(N__63889),
            .I(N__63886));
    LocalMux I__12987 (
            .O(N__63886),
            .I(N__63883));
    Span4Mux_v I__12986 (
            .O(N__63883),
            .I(N__63879));
    InMux I__12985 (
            .O(N__63882),
            .I(N__63876));
    Odrv4 I__12984 (
            .O(N__63879),
            .I(\pid_front.error_p_reg_esr_RNIQ9C61_0Z0Z_17 ));
    LocalMux I__12983 (
            .O(N__63876),
            .I(\pid_front.error_p_reg_esr_RNIQ9C61_0Z0Z_17 ));
    InMux I__12982 (
            .O(N__63871),
            .I(N__63867));
    InMux I__12981 (
            .O(N__63870),
            .I(N__63864));
    LocalMux I__12980 (
            .O(N__63867),
            .I(\pid_front.error_p_reg_esr_RNIN6C61Z0Z_16 ));
    LocalMux I__12979 (
            .O(N__63864),
            .I(\pid_front.error_p_reg_esr_RNIN6C61Z0Z_16 ));
    InMux I__12978 (
            .O(N__63859),
            .I(N__63853));
    InMux I__12977 (
            .O(N__63858),
            .I(N__63853));
    LocalMux I__12976 (
            .O(N__63853),
            .I(\pid_front.un1_pid_prereg_0_4 ));
    InMux I__12975 (
            .O(N__63850),
            .I(N__63846));
    InMux I__12974 (
            .O(N__63849),
            .I(N__63843));
    LocalMux I__12973 (
            .O(N__63846),
            .I(\pid_front.un1_pid_prereg_0_2 ));
    LocalMux I__12972 (
            .O(N__63843),
            .I(\pid_front.un1_pid_prereg_0_2 ));
    InMux I__12971 (
            .O(N__63838),
            .I(N__63833));
    InMux I__12970 (
            .O(N__63837),
            .I(N__63830));
    InMux I__12969 (
            .O(N__63836),
            .I(N__63827));
    LocalMux I__12968 (
            .O(N__63833),
            .I(\pid_front.un1_pid_prereg_0_3 ));
    LocalMux I__12967 (
            .O(N__63830),
            .I(\pid_front.un1_pid_prereg_0_3 ));
    LocalMux I__12966 (
            .O(N__63827),
            .I(\pid_front.un1_pid_prereg_0_3 ));
    CascadeMux I__12965 (
            .O(N__63820),
            .I(\pid_front.un1_pid_prereg_0_4_cascade_ ));
    InMux I__12964 (
            .O(N__63817),
            .I(N__63814));
    LocalMux I__12963 (
            .O(N__63814),
            .I(N__63811));
    Odrv4 I__12962 (
            .O(N__63811),
            .I(\pid_front.error_p_reg_esr_RNICN0DDZ0Z_15 ));
    InMux I__12961 (
            .O(N__63808),
            .I(N__63802));
    InMux I__12960 (
            .O(N__63807),
            .I(N__63802));
    LocalMux I__12959 (
            .O(N__63802),
            .I(N__63799));
    Sp12to4 I__12958 (
            .O(N__63799),
            .I(N__63796));
    Span12Mux_s7_v I__12957 (
            .O(N__63796),
            .I(N__63793));
    Odrv12 I__12956 (
            .O(N__63793),
            .I(\pid_front.error_p_regZ0Z_16 ));
    InMux I__12955 (
            .O(N__63790),
            .I(N__63784));
    InMux I__12954 (
            .O(N__63789),
            .I(N__63784));
    LocalMux I__12953 (
            .O(N__63784),
            .I(N__63781));
    Odrv4 I__12952 (
            .O(N__63781),
            .I(\pid_front.error_p_reg_esr_RNIN6C61_0Z0Z_16 ));
    InMux I__12951 (
            .O(N__63778),
            .I(N__63772));
    InMux I__12950 (
            .O(N__63777),
            .I(N__63772));
    LocalMux I__12949 (
            .O(N__63772),
            .I(\pid_front.error_d_reg_prevZ0Z_16 ));
    CascadeMux I__12948 (
            .O(N__63769),
            .I(\pid_front.error_p_reg_esr_RNIKG5U_0Z0Z_10_cascade_ ));
    CascadeMux I__12947 (
            .O(N__63766),
            .I(\pid_front.error_d_reg_prev_esr_RNI379B2Z0Z_10_cascade_ ));
    InMux I__12946 (
            .O(N__63763),
            .I(N__63758));
    InMux I__12945 (
            .O(N__63762),
            .I(N__63753));
    InMux I__12944 (
            .O(N__63761),
            .I(N__63753));
    LocalMux I__12943 (
            .O(N__63758),
            .I(\pid_front.error_d_reg_prev_esr_RNI5JRF4_0Z0Z_10 ));
    LocalMux I__12942 (
            .O(N__63753),
            .I(\pid_front.error_d_reg_prev_esr_RNI5JRF4_0Z0Z_10 ));
    InMux I__12941 (
            .O(N__63748),
            .I(N__63745));
    LocalMux I__12940 (
            .O(N__63745),
            .I(\pid_front.error_p_reg_esr_RNIKG5UZ0Z_10 ));
    InMux I__12939 (
            .O(N__63742),
            .I(N__63739));
    LocalMux I__12938 (
            .O(N__63739),
            .I(\pid_front.un1_pid_prereg_153_0 ));
    InMux I__12937 (
            .O(N__63736),
            .I(N__63727));
    InMux I__12936 (
            .O(N__63735),
            .I(N__63727));
    InMux I__12935 (
            .O(N__63734),
            .I(N__63727));
    LocalMux I__12934 (
            .O(N__63727),
            .I(\pid_front.un1_pid_prereg_0_16 ));
    InMux I__12933 (
            .O(N__63724),
            .I(N__63721));
    LocalMux I__12932 (
            .O(N__63721),
            .I(\pid_front.error_d_reg_prev_esr_RNI379B2Z0Z_10 ));
    InMux I__12931 (
            .O(N__63718),
            .I(N__63715));
    LocalMux I__12930 (
            .O(N__63715),
            .I(\pid_front.error_d_reg_prev_esr_RNI5JRF4Z0Z_10 ));
    InMux I__12929 (
            .O(N__63712),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_26 ));
    CascadeMux I__12928 (
            .O(N__63709),
            .I(N__63699));
    CascadeMux I__12927 (
            .O(N__63708),
            .I(N__63695));
    CascadeMux I__12926 (
            .O(N__63707),
            .I(N__63691));
    CascadeMux I__12925 (
            .O(N__63706),
            .I(N__63687));
    CascadeMux I__12924 (
            .O(N__63705),
            .I(N__63683));
    CascadeMux I__12923 (
            .O(N__63704),
            .I(N__63679));
    CascadeMux I__12922 (
            .O(N__63703),
            .I(N__63674));
    InMux I__12921 (
            .O(N__63702),
            .I(N__63662));
    InMux I__12920 (
            .O(N__63699),
            .I(N__63662));
    InMux I__12919 (
            .O(N__63698),
            .I(N__63662));
    InMux I__12918 (
            .O(N__63695),
            .I(N__63662));
    InMux I__12917 (
            .O(N__63694),
            .I(N__63662));
    InMux I__12916 (
            .O(N__63691),
            .I(N__63645));
    InMux I__12915 (
            .O(N__63690),
            .I(N__63645));
    InMux I__12914 (
            .O(N__63687),
            .I(N__63645));
    InMux I__12913 (
            .O(N__63686),
            .I(N__63645));
    InMux I__12912 (
            .O(N__63683),
            .I(N__63645));
    InMux I__12911 (
            .O(N__63682),
            .I(N__63645));
    InMux I__12910 (
            .O(N__63679),
            .I(N__63645));
    InMux I__12909 (
            .O(N__63678),
            .I(N__63645));
    InMux I__12908 (
            .O(N__63677),
            .I(N__63638));
    InMux I__12907 (
            .O(N__63674),
            .I(N__63638));
    InMux I__12906 (
            .O(N__63673),
            .I(N__63638));
    LocalMux I__12905 (
            .O(N__63662),
            .I(N__63635));
    LocalMux I__12904 (
            .O(N__63645),
            .I(N__63632));
    LocalMux I__12903 (
            .O(N__63638),
            .I(N__63629));
    Span4Mux_v I__12902 (
            .O(N__63635),
            .I(N__63622));
    Span4Mux_h I__12901 (
            .O(N__63632),
            .I(N__63622));
    Span4Mux_v I__12900 (
            .O(N__63629),
            .I(N__63622));
    Odrv4 I__12899 (
            .O(N__63622),
            .I(\pid_front.error_i_acummZ0Z_13 ));
    InMux I__12898 (
            .O(N__63619),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_27 ));
    InMux I__12897 (
            .O(N__63616),
            .I(N__63612));
    CascadeMux I__12896 (
            .O(N__63615),
            .I(N__63609));
    LocalMux I__12895 (
            .O(N__63612),
            .I(N__63606));
    InMux I__12894 (
            .O(N__63609),
            .I(N__63603));
    Span4Mux_v I__12893 (
            .O(N__63606),
            .I(N__63600));
    LocalMux I__12892 (
            .O(N__63603),
            .I(\pid_front.error_p_reg_esr_RNIO4E8_0Z0Z_2 ));
    Odrv4 I__12891 (
            .O(N__63600),
            .I(\pid_front.error_p_reg_esr_RNIO4E8_0Z0Z_2 ));
    InMux I__12890 (
            .O(N__63595),
            .I(N__63589));
    InMux I__12889 (
            .O(N__63594),
            .I(N__63589));
    LocalMux I__12888 (
            .O(N__63589),
            .I(N__63586));
    Odrv12 I__12887 (
            .O(N__63586),
            .I(\pid_front.error_p_regZ0Z_2 ));
    InMux I__12886 (
            .O(N__63583),
            .I(N__63577));
    InMux I__12885 (
            .O(N__63582),
            .I(N__63577));
    LocalMux I__12884 (
            .O(N__63577),
            .I(\pid_front.error_d_reg_prevZ0Z_2 ));
    InMux I__12883 (
            .O(N__63574),
            .I(N__63568));
    InMux I__12882 (
            .O(N__63573),
            .I(N__63568));
    LocalMux I__12881 (
            .O(N__63568),
            .I(\pid_front.error_p_reg_esr_RNIO4E8Z0Z_2 ));
    InMux I__12880 (
            .O(N__63565),
            .I(N__63559));
    InMux I__12879 (
            .O(N__63564),
            .I(N__63559));
    LocalMux I__12878 (
            .O(N__63559),
            .I(N__63556));
    Span4Mux_v I__12877 (
            .O(N__63556),
            .I(N__63553));
    Sp12to4 I__12876 (
            .O(N__63553),
            .I(N__63550));
    Span12Mux_h I__12875 (
            .O(N__63550),
            .I(N__63547));
    Odrv12 I__12874 (
            .O(N__63547),
            .I(\pid_front.error_p_regZ0Z_17 ));
    InMux I__12873 (
            .O(N__63544),
            .I(N__63538));
    InMux I__12872 (
            .O(N__63543),
            .I(N__63538));
    LocalMux I__12871 (
            .O(N__63538),
            .I(\pid_front.error_d_reg_prevZ0Z_17 ));
    CascadeMux I__12870 (
            .O(N__63535),
            .I(N__63532));
    InMux I__12869 (
            .O(N__63532),
            .I(N__63529));
    LocalMux I__12868 (
            .O(N__63529),
            .I(\pid_front.error_i_regZ0Z_18 ));
    InMux I__12867 (
            .O(N__63526),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_17 ));
    InMux I__12866 (
            .O(N__63523),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_18 ));
    InMux I__12865 (
            .O(N__63520),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_19 ));
    InMux I__12864 (
            .O(N__63517),
            .I(N__63514));
    LocalMux I__12863 (
            .O(N__63514),
            .I(N__63511));
    Span4Mux_v I__12862 (
            .O(N__63511),
            .I(N__63508));
    Odrv4 I__12861 (
            .O(N__63508),
            .I(\pid_front.error_i_regZ0Z_21 ));
    InMux I__12860 (
            .O(N__63505),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_20 ));
    CascadeMux I__12859 (
            .O(N__63502),
            .I(N__63499));
    InMux I__12858 (
            .O(N__63499),
            .I(N__63496));
    LocalMux I__12857 (
            .O(N__63496),
            .I(N__63493));
    Span4Mux_v I__12856 (
            .O(N__63493),
            .I(N__63490));
    Odrv4 I__12855 (
            .O(N__63490),
            .I(\pid_front.error_i_regZ0Z_22 ));
    InMux I__12854 (
            .O(N__63487),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_21 ));
    InMux I__12853 (
            .O(N__63484),
            .I(N__63481));
    LocalMux I__12852 (
            .O(N__63481),
            .I(N__63478));
    Odrv4 I__12851 (
            .O(N__63478),
            .I(\pid_front.error_i_regZ0Z_23 ));
    InMux I__12850 (
            .O(N__63475),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_22 ));
    CascadeMux I__12849 (
            .O(N__63472),
            .I(N__63469));
    InMux I__12848 (
            .O(N__63469),
            .I(N__63466));
    LocalMux I__12847 (
            .O(N__63466),
            .I(N__63463));
    Span4Mux_v I__12846 (
            .O(N__63463),
            .I(N__63460));
    Odrv4 I__12845 (
            .O(N__63460),
            .I(\pid_front.error_i_regZ0Z_24 ));
    InMux I__12844 (
            .O(N__63457),
            .I(bfn_15_22_0_));
    InMux I__12843 (
            .O(N__63454),
            .I(N__63451));
    LocalMux I__12842 (
            .O(N__63451),
            .I(N__63448));
    Span4Mux_v I__12841 (
            .O(N__63448),
            .I(N__63445));
    Odrv4 I__12840 (
            .O(N__63445),
            .I(\pid_front.error_i_regZ0Z_25 ));
    InMux I__12839 (
            .O(N__63442),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_24 ));
    CascadeMux I__12838 (
            .O(N__63439),
            .I(N__63436));
    InMux I__12837 (
            .O(N__63436),
            .I(N__63433));
    LocalMux I__12836 (
            .O(N__63433),
            .I(N__63430));
    Span4Mux_v I__12835 (
            .O(N__63430),
            .I(N__63427));
    Odrv4 I__12834 (
            .O(N__63427),
            .I(\pid_front.error_i_regZ0Z_26 ));
    InMux I__12833 (
            .O(N__63424),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_25 ));
    CascadeMux I__12832 (
            .O(N__63421),
            .I(N__63418));
    InMux I__12831 (
            .O(N__63418),
            .I(N__63415));
    LocalMux I__12830 (
            .O(N__63415),
            .I(N__63412));
    Odrv4 I__12829 (
            .O(N__63412),
            .I(\pid_front.error_i_regZ0Z_9 ));
    InMux I__12828 (
            .O(N__63409),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_8 ));
    CascadeMux I__12827 (
            .O(N__63406),
            .I(N__63403));
    InMux I__12826 (
            .O(N__63403),
            .I(N__63400));
    LocalMux I__12825 (
            .O(N__63400),
            .I(N__63397));
    Span4Mux_v I__12824 (
            .O(N__63397),
            .I(N__63394));
    Odrv4 I__12823 (
            .O(N__63394),
            .I(\pid_front.error_i_regZ0Z_10 ));
    InMux I__12822 (
            .O(N__63391),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_9 ));
    CascadeMux I__12821 (
            .O(N__63388),
            .I(N__63385));
    InMux I__12820 (
            .O(N__63385),
            .I(N__63382));
    LocalMux I__12819 (
            .O(N__63382),
            .I(N__63379));
    Span4Mux_v I__12818 (
            .O(N__63379),
            .I(N__63376));
    Odrv4 I__12817 (
            .O(N__63376),
            .I(\pid_front.error_i_regZ0Z_11 ));
    InMux I__12816 (
            .O(N__63373),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_10 ));
    InMux I__12815 (
            .O(N__63370),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_11 ));
    InMux I__12814 (
            .O(N__63367),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_12 ));
    InMux I__12813 (
            .O(N__63364),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_13 ));
    InMux I__12812 (
            .O(N__63361),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_14 ));
    InMux I__12811 (
            .O(N__63358),
            .I(bfn_15_21_0_));
    InMux I__12810 (
            .O(N__63355),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_16 ));
    InMux I__12809 (
            .O(N__63352),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_0 ));
    InMux I__12808 (
            .O(N__63349),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_1 ));
    InMux I__12807 (
            .O(N__63346),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_2 ));
    InMux I__12806 (
            .O(N__63343),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_3 ));
    CascadeMux I__12805 (
            .O(N__63340),
            .I(N__63336));
    InMux I__12804 (
            .O(N__63339),
            .I(N__63333));
    InMux I__12803 (
            .O(N__63336),
            .I(N__63330));
    LocalMux I__12802 (
            .O(N__63333),
            .I(N__63325));
    LocalMux I__12801 (
            .O(N__63330),
            .I(N__63325));
    Odrv4 I__12800 (
            .O(N__63325),
            .I(\pid_front.error_i_regZ0Z_5 ));
    InMux I__12799 (
            .O(N__63322),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_4 ));
    InMux I__12798 (
            .O(N__63319),
            .I(N__63316));
    LocalMux I__12797 (
            .O(N__63316),
            .I(N__63313));
    Odrv4 I__12796 (
            .O(N__63313),
            .I(\pid_front.error_i_regZ0Z_6 ));
    InMux I__12795 (
            .O(N__63310),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_5 ));
    CascadeMux I__12794 (
            .O(N__63307),
            .I(N__63303));
    InMux I__12793 (
            .O(N__63306),
            .I(N__63300));
    InMux I__12792 (
            .O(N__63303),
            .I(N__63297));
    LocalMux I__12791 (
            .O(N__63300),
            .I(\pid_front.error_i_regZ0Z_7 ));
    LocalMux I__12790 (
            .O(N__63297),
            .I(\pid_front.error_i_regZ0Z_7 ));
    InMux I__12789 (
            .O(N__63292),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_6 ));
    CascadeMux I__12788 (
            .O(N__63289),
            .I(N__63286));
    InMux I__12787 (
            .O(N__63286),
            .I(N__63283));
    LocalMux I__12786 (
            .O(N__63283),
            .I(N__63280));
    Odrv4 I__12785 (
            .O(N__63280),
            .I(\pid_front.error_i_regZ0Z_8 ));
    InMux I__12784 (
            .O(N__63277),
            .I(bfn_15_20_0_));
    CascadeMux I__12783 (
            .O(N__63274),
            .I(\pid_front.m13_2_03_4_i_0_o2_2_cascade_ ));
    CascadeMux I__12782 (
            .O(N__63271),
            .I(\pid_front.error_i_reg_esr_RNO_0Z0Z_9_cascade_ ));
    InMux I__12781 (
            .O(N__63268),
            .I(N__63264));
    InMux I__12780 (
            .O(N__63267),
            .I(N__63261));
    LocalMux I__12779 (
            .O(N__63264),
            .I(\pid_front.m13_2_03_4_i_0_o2_1 ));
    LocalMux I__12778 (
            .O(N__63261),
            .I(\pid_front.m13_2_03_4_i_0_o2_1 ));
    CascadeMux I__12777 (
            .O(N__63256),
            .I(\pid_front.N_184_cascade_ ));
    InMux I__12776 (
            .O(N__63253),
            .I(N__63250));
    LocalMux I__12775 (
            .O(N__63250),
            .I(N__63247));
    Odrv4 I__12774 (
            .O(N__63247),
            .I(\pid_front.N_576 ));
    CascadeMux I__12773 (
            .O(N__63244),
            .I(\pid_front.N_575_cascade_ ));
    InMux I__12772 (
            .O(N__63241),
            .I(N__63238));
    LocalMux I__12771 (
            .O(N__63238),
            .I(N__63234));
    InMux I__12770 (
            .O(N__63237),
            .I(N__63231));
    Odrv4 I__12769 (
            .O(N__63234),
            .I(\pid_front.N_229 ));
    LocalMux I__12768 (
            .O(N__63231),
            .I(\pid_front.N_229 ));
    InMux I__12767 (
            .O(N__63226),
            .I(N__63223));
    LocalMux I__12766 (
            .O(N__63223),
            .I(\pid_front.m11_2_03_3_i_3 ));
    CascadeMux I__12765 (
            .O(N__63220),
            .I(\pid_front.m11_2_03_3_i_3_cascade_ ));
    InMux I__12764 (
            .O(N__63217),
            .I(N__63214));
    LocalMux I__12763 (
            .O(N__63214),
            .I(N__63210));
    CascadeMux I__12762 (
            .O(N__63213),
            .I(N__63207));
    Span4Mux_s3_v I__12761 (
            .O(N__63210),
            .I(N__63204));
    InMux I__12760 (
            .O(N__63207),
            .I(N__63201));
    Span4Mux_v I__12759 (
            .O(N__63204),
            .I(N__63196));
    LocalMux I__12758 (
            .O(N__63201),
            .I(N__63196));
    Span4Mux_v I__12757 (
            .O(N__63196),
            .I(N__63193));
    Odrv4 I__12756 (
            .O(N__63193),
            .I(\pid_front.un1_pid_prereg_0 ));
    CascadeMux I__12755 (
            .O(N__63190),
            .I(\pid_front.error_i_reg_esr_RNO_0Z0Z_6_cascade_ ));
    InMux I__12754 (
            .O(N__63187),
            .I(N__63184));
    LocalMux I__12753 (
            .O(N__63184),
            .I(N__63181));
    Span4Mux_h I__12752 (
            .O(N__63181),
            .I(N__63178));
    Span4Mux_v I__12751 (
            .O(N__63178),
            .I(N__63174));
    InMux I__12750 (
            .O(N__63177),
            .I(N__63171));
    Odrv4 I__12749 (
            .O(N__63174),
            .I(\pid_front.N_232 ));
    LocalMux I__12748 (
            .O(N__63171),
            .I(\pid_front.N_232 ));
    InMux I__12747 (
            .O(N__63166),
            .I(N__63163));
    LocalMux I__12746 (
            .O(N__63163),
            .I(\pid_front.m10_2_03_3_i_0_o2_0 ));
    InMux I__12745 (
            .O(N__63160),
            .I(N__63157));
    LocalMux I__12744 (
            .O(N__63157),
            .I(N__63151));
    InMux I__12743 (
            .O(N__63156),
            .I(N__63146));
    InMux I__12742 (
            .O(N__63155),
            .I(N__63146));
    InMux I__12741 (
            .O(N__63154),
            .I(N__63143));
    Span4Mux_v I__12740 (
            .O(N__63151),
            .I(N__63138));
    LocalMux I__12739 (
            .O(N__63146),
            .I(N__63138));
    LocalMux I__12738 (
            .O(N__63143),
            .I(N__63133));
    Span4Mux_h I__12737 (
            .O(N__63138),
            .I(N__63133));
    Odrv4 I__12736 (
            .O(N__63133),
            .I(\pid_front.N_207 ));
    CascadeMux I__12735 (
            .O(N__63130),
            .I(N__63127));
    InMux I__12734 (
            .O(N__63127),
            .I(N__63121));
    InMux I__12733 (
            .O(N__63126),
            .I(N__63121));
    LocalMux I__12732 (
            .O(N__63121),
            .I(\pid_front.N_556 ));
    CascadeMux I__12731 (
            .O(N__63118),
            .I(\pid_front.m10_2_03_3_i_0_o2_0_cascade_ ));
    CascadeMux I__12730 (
            .O(N__63115),
            .I(\pid_front.m10_2_03_3_i_3_cascade_ ));
    InMux I__12729 (
            .O(N__63112),
            .I(N__63109));
    LocalMux I__12728 (
            .O(N__63109),
            .I(N__63106));
    Odrv4 I__12727 (
            .O(N__63106),
            .I(\pid_front.N_301 ));
    InMux I__12726 (
            .O(N__63103),
            .I(N__63100));
    LocalMux I__12725 (
            .O(N__63100),
            .I(N__63097));
    Span4Mux_h I__12724 (
            .O(N__63097),
            .I(N__63094));
    Odrv4 I__12723 (
            .O(N__63094),
            .I(\pid_front.N_510 ));
    CascadeMux I__12722 (
            .O(N__63091),
            .I(\pid_front.N_554_cascade_ ));
    InMux I__12721 (
            .O(N__63088),
            .I(N__63085));
    LocalMux I__12720 (
            .O(N__63085),
            .I(\pid_front.N_543 ));
    CascadeMux I__12719 (
            .O(N__63082),
            .I(N__63079));
    InMux I__12718 (
            .O(N__63079),
            .I(N__63076));
    LocalMux I__12717 (
            .O(N__63076),
            .I(N__63073));
    Span4Mux_v I__12716 (
            .O(N__63073),
            .I(N__63070));
    Odrv4 I__12715 (
            .O(N__63070),
            .I(pid_side_m13_2_03_4_i_0_a2_3_0));
    InMux I__12714 (
            .O(N__63067),
            .I(N__63064));
    LocalMux I__12713 (
            .O(N__63064),
            .I(\pid_front.m13_2_03_4_i_0_o2_2 ));
    InMux I__12712 (
            .O(N__63061),
            .I(N__63058));
    LocalMux I__12711 (
            .O(N__63058),
            .I(N__63055));
    Odrv4 I__12710 (
            .O(N__63055),
            .I(\pid_side.N_111 ));
    CascadeMux I__12709 (
            .O(N__63052),
            .I(\pid_front.N_161_cascade_ ));
    InMux I__12708 (
            .O(N__63049),
            .I(N__63046));
    LocalMux I__12707 (
            .O(N__63046),
            .I(\pid_front.N_398 ));
    InMux I__12706 (
            .O(N__63043),
            .I(N__63040));
    LocalMux I__12705 (
            .O(N__63040),
            .I(\pid_front.m78_0_0 ));
    CascadeMux I__12704 (
            .O(N__63037),
            .I(\pid_front.m78_0_1_cascade_ ));
    CascadeMux I__12703 (
            .O(N__63034),
            .I(N__63031));
    InMux I__12702 (
            .O(N__63031),
            .I(N__63028));
    LocalMux I__12701 (
            .O(N__63028),
            .I(\pid_front.N_626 ));
    CascadeMux I__12700 (
            .O(N__63025),
            .I(\pid_front.N_626_cascade_ ));
    CascadeMux I__12699 (
            .O(N__63022),
            .I(pid_side_N_495_cascade_));
    CascadeMux I__12698 (
            .O(N__63019),
            .I(\pid_side.m4_2_01_cascade_ ));
    InMux I__12697 (
            .O(N__63016),
            .I(N__63012));
    CascadeMux I__12696 (
            .O(N__63015),
            .I(N__63009));
    LocalMux I__12695 (
            .O(N__63012),
            .I(N__63006));
    InMux I__12694 (
            .O(N__63009),
            .I(N__63002));
    Span4Mux_h I__12693 (
            .O(N__63006),
            .I(N__62999));
    InMux I__12692 (
            .O(N__63005),
            .I(N__62996));
    LocalMux I__12691 (
            .O(N__63002),
            .I(N__62993));
    Odrv4 I__12690 (
            .O(N__62999),
            .I(\pid_side.error_i_regZ0Z_0 ));
    LocalMux I__12689 (
            .O(N__62996),
            .I(\pid_side.error_i_regZ0Z_0 ));
    Odrv12 I__12688 (
            .O(N__62993),
            .I(\pid_side.error_i_regZ0Z_0 ));
    InMux I__12687 (
            .O(N__62986),
            .I(N__62983));
    LocalMux I__12686 (
            .O(N__62983),
            .I(\pid_side.m4_2_01_1 ));
    CascadeMux I__12685 (
            .O(N__62980),
            .I(\pid_side.m64_i_o2_0_cascade_ ));
    CascadeMux I__12684 (
            .O(N__62977),
            .I(\pid_side.error_cry_1_c_RNI6K4BZ0Z1_cascade_ ));
    CascadeMux I__12683 (
            .O(N__62974),
            .I(\pid_side.error_i_reg_9_rn_0_27_cascade_ ));
    InMux I__12682 (
            .O(N__62971),
            .I(N__62968));
    LocalMux I__12681 (
            .O(N__62968),
            .I(\pid_side.N_42_i_i_0 ));
    InMux I__12680 (
            .O(N__62965),
            .I(N__62959));
    InMux I__12679 (
            .O(N__62964),
            .I(N__62959));
    LocalMux I__12678 (
            .O(N__62959),
            .I(\pid_side.error_i_regZ0Z_27 ));
    InMux I__12677 (
            .O(N__62956),
            .I(N__62953));
    LocalMux I__12676 (
            .O(N__62953),
            .I(N__62950));
    Odrv12 I__12675 (
            .O(N__62950),
            .I(\pid_side.error_i_regZ0Z_14 ));
    InMux I__12674 (
            .O(N__62947),
            .I(N__62944));
    LocalMux I__12673 (
            .O(N__62944),
            .I(N__62941));
    Span4Mux_v I__12672 (
            .O(N__62941),
            .I(N__62938));
    Odrv4 I__12671 (
            .O(N__62938),
            .I(\pid_front.error_i_reg_esr_RNO_5Z0Z_21 ));
    CascadeMux I__12670 (
            .O(N__62935),
            .I(pid_side_N_174_cascade_));
    InMux I__12669 (
            .O(N__62932),
            .I(N__62929));
    LocalMux I__12668 (
            .O(N__62929),
            .I(N__62926));
    Span4Mux_v I__12667 (
            .O(N__62926),
            .I(N__62923));
    Odrv4 I__12666 (
            .O(N__62923),
            .I(\pid_front.error_i_reg_esr_RNO_4Z0Z_21 ));
    InMux I__12665 (
            .O(N__62920),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_24 ));
    InMux I__12664 (
            .O(N__62917),
            .I(N__62912));
    InMux I__12663 (
            .O(N__62916),
            .I(N__62907));
    InMux I__12662 (
            .O(N__62915),
            .I(N__62907));
    LocalMux I__12661 (
            .O(N__62912),
            .I(\pid_side.error_i_reg_esr_RNIUHTSZ0Z_26 ));
    LocalMux I__12660 (
            .O(N__62907),
            .I(\pid_side.error_i_reg_esr_RNIUHTSZ0Z_26 ));
    InMux I__12659 (
            .O(N__62902),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_25 ));
    InMux I__12658 (
            .O(N__62899),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_26 ));
    CascadeMux I__12657 (
            .O(N__62896),
            .I(N__62890));
    CascadeMux I__12656 (
            .O(N__62895),
            .I(N__62886));
    CascadeMux I__12655 (
            .O(N__62894),
            .I(N__62877));
    InMux I__12654 (
            .O(N__62893),
            .I(N__62865));
    InMux I__12653 (
            .O(N__62890),
            .I(N__62865));
    InMux I__12652 (
            .O(N__62889),
            .I(N__62865));
    InMux I__12651 (
            .O(N__62886),
            .I(N__62865));
    InMux I__12650 (
            .O(N__62885),
            .I(N__62865));
    CascadeMux I__12649 (
            .O(N__62884),
            .I(N__62862));
    CascadeMux I__12648 (
            .O(N__62883),
            .I(N__62858));
    CascadeMux I__12647 (
            .O(N__62882),
            .I(N__62854));
    CascadeMux I__12646 (
            .O(N__62881),
            .I(N__62850));
    InMux I__12645 (
            .O(N__62880),
            .I(N__62842));
    InMux I__12644 (
            .O(N__62877),
            .I(N__62842));
    InMux I__12643 (
            .O(N__62876),
            .I(N__62842));
    LocalMux I__12642 (
            .O(N__62865),
            .I(N__62839));
    InMux I__12641 (
            .O(N__62862),
            .I(N__62822));
    InMux I__12640 (
            .O(N__62861),
            .I(N__62822));
    InMux I__12639 (
            .O(N__62858),
            .I(N__62822));
    InMux I__12638 (
            .O(N__62857),
            .I(N__62822));
    InMux I__12637 (
            .O(N__62854),
            .I(N__62822));
    InMux I__12636 (
            .O(N__62853),
            .I(N__62822));
    InMux I__12635 (
            .O(N__62850),
            .I(N__62822));
    InMux I__12634 (
            .O(N__62849),
            .I(N__62822));
    LocalMux I__12633 (
            .O(N__62842),
            .I(N__62819));
    Span4Mux_v I__12632 (
            .O(N__62839),
            .I(N__62812));
    LocalMux I__12631 (
            .O(N__62822),
            .I(N__62812));
    Span4Mux_v I__12630 (
            .O(N__62819),
            .I(N__62812));
    Span4Mux_h I__12629 (
            .O(N__62812),
            .I(N__62809));
    Span4Mux_v I__12628 (
            .O(N__62809),
            .I(N__62806));
    Span4Mux_v I__12627 (
            .O(N__62806),
            .I(N__62803));
    Odrv4 I__12626 (
            .O(N__62803),
            .I(\pid_side.error_i_acummZ0Z_13 ));
    InMux I__12625 (
            .O(N__62800),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_27 ));
    InMux I__12624 (
            .O(N__62797),
            .I(N__62794));
    LocalMux I__12623 (
            .O(N__62794),
            .I(N__62784));
    CascadeMux I__12622 (
            .O(N__62793),
            .I(N__62780));
    InMux I__12621 (
            .O(N__62792),
            .I(N__62777));
    CascadeMux I__12620 (
            .O(N__62791),
            .I(N__62773));
    InMux I__12619 (
            .O(N__62790),
            .I(N__62759));
    InMux I__12618 (
            .O(N__62789),
            .I(N__62759));
    InMux I__12617 (
            .O(N__62788),
            .I(N__62759));
    InMux I__12616 (
            .O(N__62787),
            .I(N__62759));
    Span4Mux_h I__12615 (
            .O(N__62784),
            .I(N__62756));
    InMux I__12614 (
            .O(N__62783),
            .I(N__62751));
    InMux I__12613 (
            .O(N__62780),
            .I(N__62751));
    LocalMux I__12612 (
            .O(N__62777),
            .I(N__62748));
    InMux I__12611 (
            .O(N__62776),
            .I(N__62743));
    InMux I__12610 (
            .O(N__62773),
            .I(N__62743));
    CascadeMux I__12609 (
            .O(N__62772),
            .I(N__62739));
    CascadeMux I__12608 (
            .O(N__62771),
            .I(N__62736));
    InMux I__12607 (
            .O(N__62770),
            .I(N__62733));
    InMux I__12606 (
            .O(N__62769),
            .I(N__62730));
    InMux I__12605 (
            .O(N__62768),
            .I(N__62727));
    LocalMux I__12604 (
            .O(N__62759),
            .I(N__62724));
    Span4Mux_v I__12603 (
            .O(N__62756),
            .I(N__62721));
    LocalMux I__12602 (
            .O(N__62751),
            .I(N__62714));
    Span4Mux_h I__12601 (
            .O(N__62748),
            .I(N__62714));
    LocalMux I__12600 (
            .O(N__62743),
            .I(N__62714));
    InMux I__12599 (
            .O(N__62742),
            .I(N__62707));
    InMux I__12598 (
            .O(N__62739),
            .I(N__62707));
    InMux I__12597 (
            .O(N__62736),
            .I(N__62707));
    LocalMux I__12596 (
            .O(N__62733),
            .I(N__62704));
    LocalMux I__12595 (
            .O(N__62730),
            .I(N__62699));
    LocalMux I__12594 (
            .O(N__62727),
            .I(N__62699));
    Span4Mux_v I__12593 (
            .O(N__62724),
            .I(N__62696));
    Span4Mux_h I__12592 (
            .O(N__62721),
            .I(N__62691));
    Span4Mux_v I__12591 (
            .O(N__62714),
            .I(N__62691));
    LocalMux I__12590 (
            .O(N__62707),
            .I(N__62684));
    Span4Mux_h I__12589 (
            .O(N__62704),
            .I(N__62684));
    Span4Mux_h I__12588 (
            .O(N__62699),
            .I(N__62684));
    Odrv4 I__12587 (
            .O(N__62696),
            .I(\pid_side.error_i_acumm_preregZ0Z_28 ));
    Odrv4 I__12586 (
            .O(N__62691),
            .I(\pid_side.error_i_acumm_preregZ0Z_28 ));
    Odrv4 I__12585 (
            .O(N__62684),
            .I(\pid_side.error_i_acumm_preregZ0Z_28 ));
    CascadeMux I__12584 (
            .O(N__62677),
            .I(N__62673));
    CascadeMux I__12583 (
            .O(N__62676),
            .I(N__62670));
    InMux I__12582 (
            .O(N__62673),
            .I(N__62667));
    InMux I__12581 (
            .O(N__62670),
            .I(N__62664));
    LocalMux I__12580 (
            .O(N__62667),
            .I(N__62659));
    LocalMux I__12579 (
            .O(N__62664),
            .I(N__62659));
    Span12Mux_s4_v I__12578 (
            .O(N__62659),
            .I(N__62656));
    Odrv12 I__12577 (
            .O(N__62656),
            .I(\pid_side.error_i_acumm_preregZ0Z_24 ));
    CascadeMux I__12576 (
            .O(N__62653),
            .I(N__62650));
    InMux I__12575 (
            .O(N__62650),
            .I(N__62647));
    LocalMux I__12574 (
            .O(N__62647),
            .I(N__62644));
    Odrv12 I__12573 (
            .O(N__62644),
            .I(\pid_side.error_i_regZ0Z_1 ));
    CascadeMux I__12572 (
            .O(N__62641),
            .I(\pid_side.N_302_cascade_ ));
    InMux I__12571 (
            .O(N__62638),
            .I(N__62635));
    LocalMux I__12570 (
            .O(N__62635),
            .I(\pid_side.error_i_regZ0Z_25 ));
    InMux I__12569 (
            .O(N__62632),
            .I(N__62627));
    InMux I__12568 (
            .O(N__62631),
            .I(N__62622));
    InMux I__12567 (
            .O(N__62630),
            .I(N__62622));
    LocalMux I__12566 (
            .O(N__62627),
            .I(N__62617));
    LocalMux I__12565 (
            .O(N__62622),
            .I(N__62617));
    Odrv12 I__12564 (
            .O(N__62617),
            .I(\pid_side.error_i_reg_esr_RNISCPRZ0Z_16 ));
    InMux I__12563 (
            .O(N__62614),
            .I(bfn_15_10_0_));
    InMux I__12562 (
            .O(N__62611),
            .I(N__62608));
    LocalMux I__12561 (
            .O(N__62608),
            .I(N__62603));
    InMux I__12560 (
            .O(N__62607),
            .I(N__62600));
    InMux I__12559 (
            .O(N__62606),
            .I(N__62597));
    Span4Mux_h I__12558 (
            .O(N__62603),
            .I(N__62592));
    LocalMux I__12557 (
            .O(N__62600),
            .I(N__62592));
    LocalMux I__12556 (
            .O(N__62597),
            .I(N__62589));
    Odrv4 I__12555 (
            .O(N__62592),
            .I(\pid_side.error_i_reg_esr_RNIUFQRZ0Z_17 ));
    Odrv12 I__12554 (
            .O(N__62589),
            .I(\pid_side.error_i_reg_esr_RNIUFQRZ0Z_17 ));
    InMux I__12553 (
            .O(N__62584),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_16 ));
    InMux I__12552 (
            .O(N__62581),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_17 ));
    InMux I__12551 (
            .O(N__62578),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_18 ));
    InMux I__12550 (
            .O(N__62575),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_19 ));
    InMux I__12549 (
            .O(N__62572),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_20 ));
    InMux I__12548 (
            .O(N__62569),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_21 ));
    InMux I__12547 (
            .O(N__62566),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_22 ));
    InMux I__12546 (
            .O(N__62563),
            .I(bfn_15_11_0_));
    CascadeMux I__12545 (
            .O(N__62560),
            .I(N__62557));
    InMux I__12544 (
            .O(N__62557),
            .I(N__62554));
    LocalMux I__12543 (
            .O(N__62554),
            .I(\pid_side.error_i_acummZ0Z_7 ));
    InMux I__12542 (
            .O(N__62551),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_6 ));
    InMux I__12541 (
            .O(N__62548),
            .I(N__62545));
    LocalMux I__12540 (
            .O(N__62545),
            .I(N__62542));
    Odrv4 I__12539 (
            .O(N__62542),
            .I(\pid_side.error_i_acummZ0Z_8 ));
    InMux I__12538 (
            .O(N__62539),
            .I(bfn_15_9_0_));
    InMux I__12537 (
            .O(N__62536),
            .I(N__62533));
    LocalMux I__12536 (
            .O(N__62533),
            .I(N__62530));
    Odrv4 I__12535 (
            .O(N__62530),
            .I(\pid_side.error_i_acummZ0Z_9 ));
    InMux I__12534 (
            .O(N__62527),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_8 ));
    InMux I__12533 (
            .O(N__62524),
            .I(N__62521));
    LocalMux I__12532 (
            .O(N__62521),
            .I(\pid_side.error_i_acummZ0Z_10 ));
    InMux I__12531 (
            .O(N__62518),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_9 ));
    InMux I__12530 (
            .O(N__62515),
            .I(N__62512));
    LocalMux I__12529 (
            .O(N__62512),
            .I(\pid_side.error_i_acummZ0Z_11 ));
    InMux I__12528 (
            .O(N__62509),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_10 ));
    InMux I__12527 (
            .O(N__62506),
            .I(N__62503));
    LocalMux I__12526 (
            .O(N__62503),
            .I(\pid_side.error_i_acummZ0Z_12 ));
    InMux I__12525 (
            .O(N__62500),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_11 ));
    InMux I__12524 (
            .O(N__62497),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_12 ));
    InMux I__12523 (
            .O(N__62494),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_13 ));
    InMux I__12522 (
            .O(N__62491),
            .I(N__62488));
    LocalMux I__12521 (
            .O(N__62488),
            .I(N__62484));
    InMux I__12520 (
            .O(N__62487),
            .I(N__62481));
    Span12Mux_s3_v I__12519 (
            .O(N__62484),
            .I(N__62475));
    LocalMux I__12518 (
            .O(N__62481),
            .I(N__62475));
    InMux I__12517 (
            .O(N__62480),
            .I(N__62472));
    Odrv12 I__12516 (
            .O(N__62475),
            .I(\pid_side.error_i_reg_esr_RNIQ9ORZ0Z_15 ));
    LocalMux I__12515 (
            .O(N__62472),
            .I(\pid_side.error_i_reg_esr_RNIQ9ORZ0Z_15 ));
    InMux I__12514 (
            .O(N__62467),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_14 ));
    CascadeMux I__12513 (
            .O(N__62464),
            .I(\pid_side.un1_pid_prereg_0_5_cascade_ ));
    InMux I__12512 (
            .O(N__62461),
            .I(N__62458));
    LocalMux I__12511 (
            .O(N__62458),
            .I(N__62455));
    Span4Mux_v I__12510 (
            .O(N__62455),
            .I(N__62452));
    Span4Mux_v I__12509 (
            .O(N__62452),
            .I(N__62448));
    InMux I__12508 (
            .O(N__62451),
            .I(N__62445));
    Odrv4 I__12507 (
            .O(N__62448),
            .I(\pid_side.error_i_acummZ0Z_0 ));
    LocalMux I__12506 (
            .O(N__62445),
            .I(\pid_side.error_i_acummZ0Z_0 ));
    InMux I__12505 (
            .O(N__62440),
            .I(N__62437));
    LocalMux I__12504 (
            .O(N__62437),
            .I(\pid_side.error_i_acummZ0Z_1 ));
    InMux I__12503 (
            .O(N__62434),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_0 ));
    InMux I__12502 (
            .O(N__62431),
            .I(N__62428));
    LocalMux I__12501 (
            .O(N__62428),
            .I(\pid_side.error_i_acummZ0Z_2 ));
    InMux I__12500 (
            .O(N__62425),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_1 ));
    CascadeMux I__12499 (
            .O(N__62422),
            .I(N__62418));
    InMux I__12498 (
            .O(N__62421),
            .I(N__62415));
    InMux I__12497 (
            .O(N__62418),
            .I(N__62412));
    LocalMux I__12496 (
            .O(N__62415),
            .I(N__62409));
    LocalMux I__12495 (
            .O(N__62412),
            .I(N__62404));
    Span4Mux_h I__12494 (
            .O(N__62409),
            .I(N__62404));
    Odrv4 I__12493 (
            .O(N__62404),
            .I(\pid_side.error_i_regZ0Z_3 ));
    CascadeMux I__12492 (
            .O(N__62401),
            .I(N__62398));
    InMux I__12491 (
            .O(N__62398),
            .I(N__62395));
    LocalMux I__12490 (
            .O(N__62395),
            .I(N__62392));
    Odrv4 I__12489 (
            .O(N__62392),
            .I(\pid_side.error_i_acummZ0Z_3 ));
    InMux I__12488 (
            .O(N__62389),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_2 ));
    InMux I__12487 (
            .O(N__62386),
            .I(N__62383));
    LocalMux I__12486 (
            .O(N__62383),
            .I(N__62380));
    Odrv12 I__12485 (
            .O(N__62380),
            .I(\pid_side.error_i_acummZ0Z_4 ));
    InMux I__12484 (
            .O(N__62377),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_3 ));
    InMux I__12483 (
            .O(N__62374),
            .I(N__62371));
    LocalMux I__12482 (
            .O(N__62371),
            .I(\pid_side.error_i_acummZ0Z_5 ));
    InMux I__12481 (
            .O(N__62368),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_4 ));
    InMux I__12480 (
            .O(N__62365),
            .I(N__62362));
    LocalMux I__12479 (
            .O(N__62362),
            .I(\pid_side.error_i_acummZ0Z_6 ));
    InMux I__12478 (
            .O(N__62359),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_5 ));
    InMux I__12477 (
            .O(N__62356),
            .I(N__62353));
    LocalMux I__12476 (
            .O(N__62353),
            .I(N__62350));
    Span4Mux_v I__12475 (
            .O(N__62350),
            .I(N__62347));
    Odrv4 I__12474 (
            .O(N__62347),
            .I(\pid_side.error_d_reg_prev_esr_RNI5RIOZ0Z_14 ));
    InMux I__12473 (
            .O(N__62344),
            .I(N__62340));
    InMux I__12472 (
            .O(N__62343),
            .I(N__62337));
    LocalMux I__12471 (
            .O(N__62340),
            .I(\pid_side.un1_pid_prereg_0_0 ));
    LocalMux I__12470 (
            .O(N__62337),
            .I(\pid_side.un1_pid_prereg_0_0 ));
    CascadeMux I__12469 (
            .O(N__62332),
            .I(\pid_side.un1_pid_prereg_0_0_cascade_ ));
    InMux I__12468 (
            .O(N__62329),
            .I(N__62323));
    InMux I__12467 (
            .O(N__62328),
            .I(N__62323));
    LocalMux I__12466 (
            .O(N__62323),
            .I(\pid_side.un1_pid_prereg_0_1 ));
    InMux I__12465 (
            .O(N__62320),
            .I(N__62317));
    LocalMux I__12464 (
            .O(N__62317),
            .I(N__62314));
    Odrv4 I__12463 (
            .O(N__62314),
            .I(\pid_side.error_d_reg_prev_esr_RNIB1JOZ0Z_16 ));
    CascadeMux I__12462 (
            .O(N__62311),
            .I(\pid_side.error_d_reg_prev_esr_RNIB1JOZ0Z_16_cascade_ ));
    InMux I__12461 (
            .O(N__62308),
            .I(N__62304));
    InMux I__12460 (
            .O(N__62307),
            .I(N__62301));
    LocalMux I__12459 (
            .O(N__62304),
            .I(\pid_side.un1_pid_prereg_0_2 ));
    LocalMux I__12458 (
            .O(N__62301),
            .I(\pid_side.un1_pid_prereg_0_2 ));
    InMux I__12457 (
            .O(N__62296),
            .I(N__62292));
    InMux I__12456 (
            .O(N__62295),
            .I(N__62289));
    LocalMux I__12455 (
            .O(N__62292),
            .I(\pid_side.un1_pid_prereg_0_3 ));
    LocalMux I__12454 (
            .O(N__62289),
            .I(\pid_side.un1_pid_prereg_0_3 ));
    CascadeMux I__12453 (
            .O(N__62284),
            .I(\pid_side.un1_pid_prereg_0_4_cascade_ ));
    InMux I__12452 (
            .O(N__62281),
            .I(N__62275));
    InMux I__12451 (
            .O(N__62280),
            .I(N__62275));
    LocalMux I__12450 (
            .O(N__62275),
            .I(\pid_side.error_d_reg_prevZ0Z_16 ));
    InMux I__12449 (
            .O(N__62272),
            .I(N__62266));
    InMux I__12448 (
            .O(N__62271),
            .I(N__62266));
    LocalMux I__12447 (
            .O(N__62266),
            .I(N__62263));
    Odrv4 I__12446 (
            .O(N__62263),
            .I(\pid_side.error_d_reg_prev_esr_RNIB1JO_0Z0Z_16 ));
    InMux I__12445 (
            .O(N__62260),
            .I(N__62256));
    InMux I__12444 (
            .O(N__62259),
            .I(N__62253));
    LocalMux I__12443 (
            .O(N__62256),
            .I(\pid_side.error_d_reg_prev_esr_RNIE4JO_0Z0Z_17 ));
    LocalMux I__12442 (
            .O(N__62253),
            .I(\pid_side.error_d_reg_prev_esr_RNIE4JO_0Z0Z_17 ));
    InMux I__12441 (
            .O(N__62248),
            .I(N__62245));
    LocalMux I__12440 (
            .O(N__62245),
            .I(N__62241));
    InMux I__12439 (
            .O(N__62244),
            .I(N__62238));
    Odrv4 I__12438 (
            .O(N__62241),
            .I(\pid_side.un11lto30_i_a2_6_and ));
    LocalMux I__12437 (
            .O(N__62238),
            .I(\pid_side.un11lto30_i_a2_6_and ));
    InMux I__12436 (
            .O(N__62233),
            .I(N__62229));
    InMux I__12435 (
            .O(N__62232),
            .I(N__62226));
    LocalMux I__12434 (
            .O(N__62229),
            .I(N__62223));
    LocalMux I__12433 (
            .O(N__62226),
            .I(\pid_side.un11lto30_i_a2_3_and ));
    Odrv4 I__12432 (
            .O(N__62223),
            .I(\pid_side.un11lto30_i_a2_3_and ));
    InMux I__12431 (
            .O(N__62218),
            .I(N__62214));
    InMux I__12430 (
            .O(N__62217),
            .I(N__62211));
    LocalMux I__12429 (
            .O(N__62214),
            .I(N__62208));
    LocalMux I__12428 (
            .O(N__62211),
            .I(\pid_side.un11lto30_i_a2_4_and ));
    Odrv4 I__12427 (
            .O(N__62208),
            .I(\pid_side.un11lto30_i_a2_4_and ));
    CascadeMux I__12426 (
            .O(N__62203),
            .I(\pid_side.un1_pid_prereg_0_1_cascade_ ));
    CascadeMux I__12425 (
            .O(N__62200),
            .I(\pid_side.un1_pid_prereg_0_2_cascade_ ));
    CascadeMux I__12424 (
            .O(N__62197),
            .I(\pid_side.un1_pid_prereg_0_3_cascade_ ));
    InMux I__12423 (
            .O(N__62194),
            .I(N__62190));
    InMux I__12422 (
            .O(N__62193),
            .I(N__62187));
    LocalMux I__12421 (
            .O(N__62190),
            .I(\pid_side.error_i_acumm_preregZ0Z_20 ));
    LocalMux I__12420 (
            .O(N__62187),
            .I(\pid_side.error_i_acumm_preregZ0Z_20 ));
    InMux I__12419 (
            .O(N__62182),
            .I(N__62178));
    InMux I__12418 (
            .O(N__62181),
            .I(N__62175));
    LocalMux I__12417 (
            .O(N__62178),
            .I(\pid_side.error_i_acumm_preregZ0Z_21 ));
    LocalMux I__12416 (
            .O(N__62175),
            .I(\pid_side.error_i_acumm_preregZ0Z_21 ));
    CascadeMux I__12415 (
            .O(N__62170),
            .I(N__62166));
    CascadeMux I__12414 (
            .O(N__62169),
            .I(N__62163));
    InMux I__12413 (
            .O(N__62166),
            .I(N__62160));
    InMux I__12412 (
            .O(N__62163),
            .I(N__62157));
    LocalMux I__12411 (
            .O(N__62160),
            .I(\pid_side.error_i_acumm_preregZ0Z_23 ));
    LocalMux I__12410 (
            .O(N__62157),
            .I(\pid_side.error_i_acumm_preregZ0Z_23 ));
    InMux I__12409 (
            .O(N__62152),
            .I(N__62148));
    InMux I__12408 (
            .O(N__62151),
            .I(N__62145));
    LocalMux I__12407 (
            .O(N__62148),
            .I(N__62142));
    LocalMux I__12406 (
            .O(N__62145),
            .I(N__62139));
    Span4Mux_h I__12405 (
            .O(N__62142),
            .I(N__62136));
    Odrv4 I__12404 (
            .O(N__62139),
            .I(\pid_side.error_i_acumm_preregZ0Z_17 ));
    Odrv4 I__12403 (
            .O(N__62136),
            .I(\pid_side.error_i_acumm_preregZ0Z_17 ));
    InMux I__12402 (
            .O(N__62131),
            .I(N__62128));
    LocalMux I__12401 (
            .O(N__62128),
            .I(N__62125));
    Span4Mux_h I__12400 (
            .O(N__62125),
            .I(N__62122));
    Odrv4 I__12399 (
            .O(N__62122),
            .I(\pid_side.error_i_acumm_13_i_o2_0_9_3 ));
    InMux I__12398 (
            .O(N__62119),
            .I(N__62115));
    InMux I__12397 (
            .O(N__62118),
            .I(N__62112));
    LocalMux I__12396 (
            .O(N__62115),
            .I(\pid_side.error_i_acumm_preregZ0Z_15 ));
    LocalMux I__12395 (
            .O(N__62112),
            .I(\pid_side.error_i_acumm_preregZ0Z_15 ));
    InMux I__12394 (
            .O(N__62107),
            .I(N__62103));
    InMux I__12393 (
            .O(N__62106),
            .I(N__62100));
    LocalMux I__12392 (
            .O(N__62103),
            .I(\pid_side.error_i_acumm_preregZ0Z_16 ));
    LocalMux I__12391 (
            .O(N__62100),
            .I(\pid_side.error_i_acumm_preregZ0Z_16 ));
    InMux I__12390 (
            .O(N__62095),
            .I(N__62092));
    LocalMux I__12389 (
            .O(N__62092),
            .I(N__62089));
    Odrv4 I__12388 (
            .O(N__62089),
            .I(\pid_side.un11lto30_i_a2_5_and ));
    CascadeMux I__12387 (
            .O(N__62086),
            .I(\pid_side.un11lto30_i_a2_5_and_cascade_ ));
    InMux I__12386 (
            .O(N__62083),
            .I(N__62080));
    LocalMux I__12385 (
            .O(N__62080),
            .I(N__62076));
    InMux I__12384 (
            .O(N__62079),
            .I(N__62073));
    Odrv12 I__12383 (
            .O(N__62076),
            .I(\pid_side.N_175 ));
    LocalMux I__12382 (
            .O(N__62073),
            .I(\pid_side.N_175 ));
    CascadeMux I__12381 (
            .O(N__62068),
            .I(\pid_side.N_175_cascade_ ));
    InMux I__12380 (
            .O(N__62065),
            .I(N__62061));
    InMux I__12379 (
            .O(N__62064),
            .I(N__62058));
    LocalMux I__12378 (
            .O(N__62061),
            .I(N__62051));
    LocalMux I__12377 (
            .O(N__62058),
            .I(N__62051));
    InMux I__12376 (
            .O(N__62057),
            .I(N__62046));
    InMux I__12375 (
            .O(N__62056),
            .I(N__62046));
    Odrv4 I__12374 (
            .O(N__62051),
            .I(\pid_side.pid_preregZ0Z_14 ));
    LocalMux I__12373 (
            .O(N__62046),
            .I(\pid_side.pid_preregZ0Z_14 ));
    InMux I__12372 (
            .O(N__62041),
            .I(N__62036));
    InMux I__12371 (
            .O(N__62040),
            .I(N__62031));
    InMux I__12370 (
            .O(N__62039),
            .I(N__62031));
    LocalMux I__12369 (
            .O(N__62036),
            .I(N__62028));
    LocalMux I__12368 (
            .O(N__62031),
            .I(N__62025));
    Span4Mux_h I__12367 (
            .O(N__62028),
            .I(N__62022));
    Odrv4 I__12366 (
            .O(N__62025),
            .I(\pid_side.N_277 ));
    Odrv4 I__12365 (
            .O(N__62022),
            .I(\pid_side.N_277 ));
    InMux I__12364 (
            .O(N__62017),
            .I(N__62014));
    LocalMux I__12363 (
            .O(N__62014),
            .I(N__62010));
    InMux I__12362 (
            .O(N__62013),
            .I(N__62007));
    Odrv4 I__12361 (
            .O(N__62010),
            .I(\pid_side.error_i_acumm_preregZ0Z_14 ));
    LocalMux I__12360 (
            .O(N__62007),
            .I(\pid_side.error_i_acumm_preregZ0Z_14 ));
    InMux I__12359 (
            .O(N__62002),
            .I(N__61999));
    LocalMux I__12358 (
            .O(N__61999),
            .I(N__61996));
    Span4Mux_v I__12357 (
            .O(N__61996),
            .I(N__61993));
    Span4Mux_v I__12356 (
            .O(N__61993),
            .I(N__61990));
    Odrv4 I__12355 (
            .O(N__61990),
            .I(\pid_side.error_i_acumm_13_i_o2_0_10_12 ));
    InMux I__12354 (
            .O(N__61987),
            .I(N__61984));
    LocalMux I__12353 (
            .O(N__61984),
            .I(\pid_side.error_i_acumm_13_i_o2_0_8_12 ));
    CascadeMux I__12352 (
            .O(N__61981),
            .I(\pid_side.error_i_acumm_13_i_o2_0_9_12_cascade_ ));
    InMux I__12351 (
            .O(N__61978),
            .I(N__61975));
    LocalMux I__12350 (
            .O(N__61975),
            .I(\pid_side.error_i_acumm_13_i_o2_0_7_12 ));
    InMux I__12349 (
            .O(N__61972),
            .I(N__61969));
    LocalMux I__12348 (
            .O(N__61969),
            .I(N__61963));
    InMux I__12347 (
            .O(N__61968),
            .I(N__61958));
    InMux I__12346 (
            .O(N__61967),
            .I(N__61958));
    InMux I__12345 (
            .O(N__61966),
            .I(N__61955));
    Span4Mux_v I__12344 (
            .O(N__61963),
            .I(N__61952));
    LocalMux I__12343 (
            .O(N__61958),
            .I(N__61949));
    LocalMux I__12342 (
            .O(N__61955),
            .I(N__61944));
    Span4Mux_s2_v I__12341 (
            .O(N__61952),
            .I(N__61944));
    Span4Mux_v I__12340 (
            .O(N__61949),
            .I(N__61941));
    Odrv4 I__12339 (
            .O(N__61944),
            .I(\pid_side.N_203 ));
    Odrv4 I__12338 (
            .O(N__61941),
            .I(\pid_side.N_203 ));
    InMux I__12337 (
            .O(N__61936),
            .I(N__61933));
    LocalMux I__12336 (
            .O(N__61933),
            .I(N__61929));
    InMux I__12335 (
            .O(N__61932),
            .I(N__61926));
    Odrv4 I__12334 (
            .O(N__61929),
            .I(\pid_side.error_i_acumm_preregZ0Z_22 ));
    LocalMux I__12333 (
            .O(N__61926),
            .I(\pid_side.error_i_acumm_preregZ0Z_22 ));
    InMux I__12332 (
            .O(N__61921),
            .I(N__61918));
    LocalMux I__12331 (
            .O(N__61918),
            .I(N__61914));
    InMux I__12330 (
            .O(N__61917),
            .I(N__61911));
    Odrv4 I__12329 (
            .O(N__61914),
            .I(\pid_side.error_i_acumm_preregZ0Z_27 ));
    LocalMux I__12328 (
            .O(N__61911),
            .I(\pid_side.error_i_acumm_preregZ0Z_27 ));
    InMux I__12327 (
            .O(N__61906),
            .I(N__61903));
    LocalMux I__12326 (
            .O(N__61903),
            .I(N__61900));
    Span4Mux_s3_v I__12325 (
            .O(N__61900),
            .I(N__61897));
    Odrv4 I__12324 (
            .O(N__61897),
            .I(\pid_side.error_i_acumm_13_i_o2_0_8_3 ));
    InMux I__12323 (
            .O(N__61894),
            .I(N__61890));
    InMux I__12322 (
            .O(N__61893),
            .I(N__61887));
    LocalMux I__12321 (
            .O(N__61890),
            .I(\pid_side.error_i_acumm_preregZ0Z_19 ));
    LocalMux I__12320 (
            .O(N__61887),
            .I(\pid_side.error_i_acumm_preregZ0Z_19 ));
    CascadeMux I__12319 (
            .O(N__61882),
            .I(\pid_front.un1_pid_prereg_0_20_cascade_ ));
    CascadeMux I__12318 (
            .O(N__61879),
            .I(N__61876));
    InMux I__12317 (
            .O(N__61876),
            .I(N__61873));
    LocalMux I__12316 (
            .O(N__61873),
            .I(\pid_front.error_d_reg_prev_esr_RNI642C4Z0Z_21 ));
    CascadeMux I__12315 (
            .O(N__61870),
            .I(\pid_front.un1_pid_prereg_0_22_cascade_ ));
    InMux I__12314 (
            .O(N__61867),
            .I(N__61864));
    LocalMux I__12313 (
            .O(N__61864),
            .I(\pid_front.error_d_reg_prev_esr_RNIGE6O8Z0Z_21 ));
    InMux I__12312 (
            .O(N__61861),
            .I(N__61858));
    LocalMux I__12311 (
            .O(N__61858),
            .I(N__61855));
    Span4Mux_v I__12310 (
            .O(N__61855),
            .I(N__61851));
    InMux I__12309 (
            .O(N__61854),
            .I(N__61848));
    Odrv4 I__12308 (
            .O(N__61851),
            .I(\pid_front.un1_pid_prereg_0_18 ));
    LocalMux I__12307 (
            .O(N__61848),
            .I(\pid_front.un1_pid_prereg_0_18 ));
    CascadeMux I__12306 (
            .O(N__61843),
            .I(N__61840));
    InMux I__12305 (
            .O(N__61840),
            .I(N__61837));
    LocalMux I__12304 (
            .O(N__61837),
            .I(N__61833));
    InMux I__12303 (
            .O(N__61836),
            .I(N__61830));
    Odrv4 I__12302 (
            .O(N__61833),
            .I(\pid_front.un1_pid_prereg_0_19 ));
    LocalMux I__12301 (
            .O(N__61830),
            .I(\pid_front.un1_pid_prereg_0_19 ));
    InMux I__12300 (
            .O(N__61825),
            .I(N__61821));
    InMux I__12299 (
            .O(N__61824),
            .I(N__61818));
    LocalMux I__12298 (
            .O(N__61821),
            .I(\pid_front.un1_pid_prereg_0_20 ));
    LocalMux I__12297 (
            .O(N__61818),
            .I(\pid_front.un1_pid_prereg_0_20 ));
    InMux I__12296 (
            .O(N__61813),
            .I(N__61810));
    LocalMux I__12295 (
            .O(N__61810),
            .I(\pid_front.error_d_reg_prev_esr_RNI822O8Z0Z_21 ));
    CascadeMux I__12294 (
            .O(N__61807),
            .I(\pid_front.un1_pid_prereg_0_23_cascade_ ));
    CascadeMux I__12293 (
            .O(N__61804),
            .I(N__61801));
    InMux I__12292 (
            .O(N__61801),
            .I(N__61798));
    LocalMux I__12291 (
            .O(N__61798),
            .I(\pid_front.error_d_reg_prev_esr_RNIAA4C4Z0Z_21 ));
    InMux I__12290 (
            .O(N__61795),
            .I(N__61786));
    InMux I__12289 (
            .O(N__61794),
            .I(N__61786));
    InMux I__12288 (
            .O(N__61793),
            .I(N__61786));
    LocalMux I__12287 (
            .O(N__61786),
            .I(\pid_front.un1_pid_prereg_0_21 ));
    InMux I__12286 (
            .O(N__61783),
            .I(N__61779));
    CascadeMux I__12285 (
            .O(N__61782),
            .I(N__61775));
    LocalMux I__12284 (
            .O(N__61779),
            .I(N__61772));
    InMux I__12283 (
            .O(N__61778),
            .I(N__61767));
    InMux I__12282 (
            .O(N__61775),
            .I(N__61767));
    Span4Mux_h I__12281 (
            .O(N__61772),
            .I(N__61764));
    LocalMux I__12280 (
            .O(N__61767),
            .I(\pid_front.error_p_regZ0Z_6 ));
    Odrv4 I__12279 (
            .O(N__61764),
            .I(\pid_front.error_p_regZ0Z_6 ));
    InMux I__12278 (
            .O(N__61759),
            .I(N__61756));
    LocalMux I__12277 (
            .O(N__61756),
            .I(\pid_front.error_p_reg_esr_RNIMVC9_0Z0Z_6 ));
    CascadeMux I__12276 (
            .O(N__61753),
            .I(N__61750));
    InMux I__12275 (
            .O(N__61750),
            .I(N__61747));
    LocalMux I__12274 (
            .O(N__61747),
            .I(N__61744));
    Odrv4 I__12273 (
            .O(N__61744),
            .I(\pid_front.error_p_reg_esr_RNIJ26O1Z0Z_5 ));
    CascadeMux I__12272 (
            .O(N__61741),
            .I(N__61738));
    InMux I__12271 (
            .O(N__61738),
            .I(N__61732));
    InMux I__12270 (
            .O(N__61737),
            .I(N__61732));
    LocalMux I__12269 (
            .O(N__61732),
            .I(\pid_front.error_d_reg_prev_esr_RNISAJOZ0Z_6 ));
    CascadeMux I__12268 (
            .O(N__61729),
            .I(\pid_front.un1_pid_prereg_66_0_cascade_ ));
    InMux I__12267 (
            .O(N__61726),
            .I(N__61723));
    LocalMux I__12266 (
            .O(N__61723),
            .I(N__61720));
    Odrv4 I__12265 (
            .O(N__61720),
            .I(\pid_front.error_p_reg_esr_RNIUBTV2Z0Z_5 ));
    InMux I__12264 (
            .O(N__61717),
            .I(N__61711));
    InMux I__12263 (
            .O(N__61716),
            .I(N__61711));
    LocalMux I__12262 (
            .O(N__61711),
            .I(\pid_front.error_p_reg_esr_RNIVOSGZ0Z_5 ));
    InMux I__12261 (
            .O(N__61708),
            .I(N__61701));
    InMux I__12260 (
            .O(N__61707),
            .I(N__61698));
    InMux I__12259 (
            .O(N__61706),
            .I(N__61691));
    InMux I__12258 (
            .O(N__61705),
            .I(N__61691));
    InMux I__12257 (
            .O(N__61704),
            .I(N__61691));
    LocalMux I__12256 (
            .O(N__61701),
            .I(\pid_front.error_d_reg_prevZ0Z_5 ));
    LocalMux I__12255 (
            .O(N__61698),
            .I(\pid_front.error_d_reg_prevZ0Z_5 ));
    LocalMux I__12254 (
            .O(N__61691),
            .I(\pid_front.error_d_reg_prevZ0Z_5 ));
    CascadeMux I__12253 (
            .O(N__61684),
            .I(N__61681));
    InMux I__12252 (
            .O(N__61681),
            .I(N__61675));
    InMux I__12251 (
            .O(N__61680),
            .I(N__61675));
    LocalMux I__12250 (
            .O(N__61675),
            .I(N__61672));
    Odrv12 I__12249 (
            .O(N__61672),
            .I(\pid_front.error_p_reg_esr_RNIUAE8Z0Z_4 ));
    CascadeMux I__12248 (
            .O(N__61669),
            .I(N__61665));
    InMux I__12247 (
            .O(N__61668),
            .I(N__61660));
    InMux I__12246 (
            .O(N__61665),
            .I(N__61660));
    LocalMux I__12245 (
            .O(N__61660),
            .I(N__61657));
    Span12Mux_h I__12244 (
            .O(N__61657),
            .I(N__61654));
    Odrv12 I__12243 (
            .O(N__61654),
            .I(\pid_front.error_p_regZ0Z_5 ));
    InMux I__12242 (
            .O(N__61651),
            .I(N__61647));
    InMux I__12241 (
            .O(N__61650),
            .I(N__61644));
    LocalMux I__12240 (
            .O(N__61647),
            .I(N__61641));
    LocalMux I__12239 (
            .O(N__61644),
            .I(\pid_front.error_p_reg_esr_RNIVOSG_0Z0Z_5 ));
    Odrv12 I__12238 (
            .O(N__61641),
            .I(\pid_front.error_p_reg_esr_RNIVOSG_0Z0Z_5 ));
    CascadeMux I__12237 (
            .O(N__61636),
            .I(\pid_front.error_p_reg_esr_RNIVOSG_0Z0Z_5_cascade_ ));
    InMux I__12236 (
            .O(N__61633),
            .I(N__61629));
    InMux I__12235 (
            .O(N__61632),
            .I(N__61626));
    LocalMux I__12234 (
            .O(N__61629),
            .I(N__61623));
    LocalMux I__12233 (
            .O(N__61626),
            .I(N__61620));
    Span4Mux_h I__12232 (
            .O(N__61623),
            .I(N__61617));
    Odrv12 I__12231 (
            .O(N__61620),
            .I(\pid_front.error_p_reg_esr_RNIB9N71_0Z0Z_5 ));
    Odrv4 I__12230 (
            .O(N__61617),
            .I(\pid_front.error_p_reg_esr_RNIB9N71_0Z0Z_5 ));
    InMux I__12229 (
            .O(N__61612),
            .I(N__61609));
    LocalMux I__12228 (
            .O(N__61609),
            .I(\pid_front.error_d_reg_prev_esr_RNIQ9AEDZ0Z_10 ));
    CascadeMux I__12227 (
            .O(N__61606),
            .I(\pid_front.un1_pid_prereg_0_17_cascade_ ));
    CascadeMux I__12226 (
            .O(N__61603),
            .I(N__61600));
    InMux I__12225 (
            .O(N__61600),
            .I(N__61597));
    LocalMux I__12224 (
            .O(N__61597),
            .I(\pid_front.error_d_reg_prev_esr_RNIUNTB4Z0Z_21 ));
    CascadeMux I__12223 (
            .O(N__61594),
            .I(\pid_front.un1_pid_prereg_0_18_cascade_ ));
    InMux I__12222 (
            .O(N__61591),
            .I(N__61588));
    LocalMux I__12221 (
            .O(N__61588),
            .I(\pid_front.error_d_reg_prev_esr_RNI0MTN8Z0Z_21 ));
    InMux I__12220 (
            .O(N__61585),
            .I(N__61582));
    LocalMux I__12219 (
            .O(N__61582),
            .I(N__61579));
    Span4Mux_v I__12218 (
            .O(N__61579),
            .I(N__61575));
    InMux I__12217 (
            .O(N__61578),
            .I(N__61572));
    Odrv4 I__12216 (
            .O(N__61575),
            .I(\pid_front.un1_pid_prereg_0_14 ));
    LocalMux I__12215 (
            .O(N__61572),
            .I(\pid_front.un1_pid_prereg_0_14 ));
    CascadeMux I__12214 (
            .O(N__61567),
            .I(N__61564));
    InMux I__12213 (
            .O(N__61564),
            .I(N__61561));
    LocalMux I__12212 (
            .O(N__61561),
            .I(N__61558));
    Span4Mux_v I__12211 (
            .O(N__61558),
            .I(N__61554));
    InMux I__12210 (
            .O(N__61557),
            .I(N__61551));
    Odrv4 I__12209 (
            .O(N__61554),
            .I(\pid_front.un1_pid_prereg_0_15 ));
    LocalMux I__12208 (
            .O(N__61551),
            .I(\pid_front.un1_pid_prereg_0_15 ));
    InMux I__12207 (
            .O(N__61546),
            .I(N__61542));
    InMux I__12206 (
            .O(N__61545),
            .I(N__61539));
    LocalMux I__12205 (
            .O(N__61542),
            .I(\pid_front.un1_pid_prereg_0_17 ));
    LocalMux I__12204 (
            .O(N__61539),
            .I(\pid_front.un1_pid_prereg_0_17 ));
    InMux I__12203 (
            .O(N__61534),
            .I(N__61531));
    LocalMux I__12202 (
            .O(N__61531),
            .I(\pid_front.error_d_reg_prev_esr_RNIO9PN8Z0Z_21 ));
    CascadeMux I__12201 (
            .O(N__61528),
            .I(N__61525));
    InMux I__12200 (
            .O(N__61525),
            .I(N__61522));
    LocalMux I__12199 (
            .O(N__61522),
            .I(\pid_front.error_p_reg_esr_RNIE2FM6Z0Z_15 ));
    CascadeMux I__12198 (
            .O(N__61519),
            .I(\pid_front.un1_pid_prereg_0_19_cascade_ ));
    CascadeMux I__12197 (
            .O(N__61516),
            .I(N__61513));
    InMux I__12196 (
            .O(N__61513),
            .I(N__61510));
    LocalMux I__12195 (
            .O(N__61510),
            .I(\pid_front.error_d_reg_prev_esr_RNI2UVB4Z0Z_21 ));
    CascadeMux I__12194 (
            .O(N__61507),
            .I(N__61504));
    InMux I__12193 (
            .O(N__61504),
            .I(N__61501));
    LocalMux I__12192 (
            .O(N__61501),
            .I(\pid_front.error_p_reg_esr_RNIB9N71Z0Z_5 ));
    CascadeMux I__12191 (
            .O(N__61498),
            .I(\pid_front.un1_pid_prereg_0_1_cascade_ ));
    CascadeMux I__12190 (
            .O(N__61495),
            .I(N__61492));
    InMux I__12189 (
            .O(N__61492),
            .I(N__61489));
    LocalMux I__12188 (
            .O(N__61489),
            .I(\pid_front.error_p_reg_esr_RNIUFCM6Z0Z_14 ));
    CascadeMux I__12187 (
            .O(N__61486),
            .I(\pid_front.un1_pid_prereg_0_2_cascade_ ));
    InMux I__12186 (
            .O(N__61483),
            .I(N__61480));
    LocalMux I__12185 (
            .O(N__61480),
            .I(\pid_front.error_p_reg_esr_RNICIRCDZ0Z_14 ));
    InMux I__12184 (
            .O(N__61477),
            .I(N__61471));
    InMux I__12183 (
            .O(N__61476),
            .I(N__61471));
    LocalMux I__12182 (
            .O(N__61471),
            .I(\pid_front.un1_pid_prereg_0_0 ));
    InMux I__12181 (
            .O(N__61468),
            .I(N__61462));
    InMux I__12180 (
            .O(N__61467),
            .I(N__61462));
    LocalMux I__12179 (
            .O(N__61462),
            .I(\pid_front.un1_pid_prereg_0_1 ));
    CascadeMux I__12178 (
            .O(N__61459),
            .I(\pid_front.un1_pid_prereg_0_0_cascade_ ));
    CascadeMux I__12177 (
            .O(N__61456),
            .I(N__61453));
    InMux I__12176 (
            .O(N__61453),
            .I(N__61450));
    LocalMux I__12175 (
            .O(N__61450),
            .I(N__61447));
    Odrv4 I__12174 (
            .O(N__61447),
            .I(\pid_front.error_p_reg_esr_RNIA6C3NZ0Z_14 ));
    CascadeMux I__12173 (
            .O(N__61444),
            .I(N__61440));
    InMux I__12172 (
            .O(N__61443),
            .I(N__61437));
    InMux I__12171 (
            .O(N__61440),
            .I(N__61434));
    LocalMux I__12170 (
            .O(N__61437),
            .I(\pid_front.error_p_reg_esr_RNIPKK71Z0Z_2 ));
    LocalMux I__12169 (
            .O(N__61434),
            .I(\pid_front.error_p_reg_esr_RNIPKK71Z0Z_2 ));
    InMux I__12168 (
            .O(N__61429),
            .I(N__61423));
    InMux I__12167 (
            .O(N__61428),
            .I(N__61423));
    LocalMux I__12166 (
            .O(N__61423),
            .I(N__61420));
    Span4Mux_v I__12165 (
            .O(N__61420),
            .I(N__61417));
    Span4Mux_h I__12164 (
            .O(N__61417),
            .I(N__61414));
    Span4Mux_h I__12163 (
            .O(N__61414),
            .I(N__61411));
    Odrv4 I__12162 (
            .O(N__61411),
            .I(\pid_front.error_p_regZ0Z_3 ));
    CascadeMux I__12161 (
            .O(N__61408),
            .I(N__61405));
    InMux I__12160 (
            .O(N__61405),
            .I(N__61399));
    InMux I__12159 (
            .O(N__61404),
            .I(N__61399));
    LocalMux I__12158 (
            .O(N__61399),
            .I(\pid_front.error_d_reg_prevZ0Z_3 ));
    InMux I__12157 (
            .O(N__61396),
            .I(N__61393));
    LocalMux I__12156 (
            .O(N__61393),
            .I(\pid_front.error_p_reg_esr_RNIR7E8_0Z0Z_3 ));
    CascadeMux I__12155 (
            .O(N__61390),
            .I(\pid_front.error_p_reg_esr_RNIR7E8_0Z0Z_3_cascade_ ));
    CascadeMux I__12154 (
            .O(N__61387),
            .I(N__61384));
    InMux I__12153 (
            .O(N__61384),
            .I(N__61381));
    LocalMux I__12152 (
            .O(N__61381),
            .I(\pid_front.error_p_reg_esr_RNIQ7CF2Z0Z_2 ));
    InMux I__12151 (
            .O(N__61378),
            .I(N__61375));
    LocalMux I__12150 (
            .O(N__61375),
            .I(N__61372));
    Span4Mux_h I__12149 (
            .O(N__61372),
            .I(N__61368));
    InMux I__12148 (
            .O(N__61371),
            .I(N__61365));
    Span4Mux_v I__12147 (
            .O(N__61368),
            .I(N__61360));
    LocalMux I__12146 (
            .O(N__61365),
            .I(N__61357));
    InMux I__12145 (
            .O(N__61364),
            .I(N__61352));
    InMux I__12144 (
            .O(N__61363),
            .I(N__61352));
    Odrv4 I__12143 (
            .O(N__61360),
            .I(\pid_front.error_d_reg_prevZ0Z_1 ));
    Odrv4 I__12142 (
            .O(N__61357),
            .I(\pid_front.error_d_reg_prevZ0Z_1 ));
    LocalMux I__12141 (
            .O(N__61352),
            .I(\pid_front.error_d_reg_prevZ0Z_1 ));
    InMux I__12140 (
            .O(N__61345),
            .I(N__61342));
    LocalMux I__12139 (
            .O(N__61342),
            .I(N__61339));
    Span4Mux_v I__12138 (
            .O(N__61339),
            .I(N__61331));
    InMux I__12137 (
            .O(N__61338),
            .I(N__61328));
    InMux I__12136 (
            .O(N__61337),
            .I(N__61319));
    InMux I__12135 (
            .O(N__61336),
            .I(N__61319));
    InMux I__12134 (
            .O(N__61335),
            .I(N__61319));
    InMux I__12133 (
            .O(N__61334),
            .I(N__61319));
    Odrv4 I__12132 (
            .O(N__61331),
            .I(\pid_front.error_d_regZ0Z_1 ));
    LocalMux I__12131 (
            .O(N__61328),
            .I(\pid_front.error_d_regZ0Z_1 ));
    LocalMux I__12130 (
            .O(N__61319),
            .I(\pid_front.error_d_regZ0Z_1 ));
    InMux I__12129 (
            .O(N__61312),
            .I(N__61309));
    LocalMux I__12128 (
            .O(N__61309),
            .I(N__61306));
    Span4Mux_h I__12127 (
            .O(N__61306),
            .I(N__61303));
    Span4Mux_v I__12126 (
            .O(N__61303),
            .I(N__61299));
    InMux I__12125 (
            .O(N__61302),
            .I(N__61296));
    Odrv4 I__12124 (
            .O(N__61299),
            .I(\pid_front.error_d_reg_prev_esr_RNIFSHOZ0Z_1 ));
    LocalMux I__12123 (
            .O(N__61296),
            .I(\pid_front.error_d_reg_prev_esr_RNIFSHOZ0Z_1 ));
    InMux I__12122 (
            .O(N__61291),
            .I(N__61287));
    InMux I__12121 (
            .O(N__61290),
            .I(N__61284));
    LocalMux I__12120 (
            .O(N__61287),
            .I(\pid_front.error_d_reg_prev_esr_RNI1JN71Z0Z_1 ));
    LocalMux I__12119 (
            .O(N__61284),
            .I(\pid_front.error_d_reg_prev_esr_RNI1JN71Z0Z_1 ));
    IoInMux I__12118 (
            .O(N__61279),
            .I(N__61276));
    LocalMux I__12117 (
            .O(N__61276),
            .I(N__61273));
    Span4Mux_s3_v I__12116 (
            .O(N__61273),
            .I(N__61270));
    Span4Mux_v I__12115 (
            .O(N__61270),
            .I(N__61267));
    Odrv4 I__12114 (
            .O(N__61267),
            .I(\pid_alt.state_0_0 ));
    CascadeMux I__12113 (
            .O(N__61264),
            .I(N__61261));
    InMux I__12112 (
            .O(N__61261),
            .I(N__61258));
    LocalMux I__12111 (
            .O(N__61258),
            .I(\pid_front.error_d_reg_prev_esr_RNI1K4E5Z0Z_10 ));
    InMux I__12110 (
            .O(N__61255),
            .I(N__61249));
    InMux I__12109 (
            .O(N__61254),
            .I(N__61249));
    LocalMux I__12108 (
            .O(N__61249),
            .I(N__61246));
    Odrv4 I__12107 (
            .O(N__61246),
            .I(\pid_front.N_2370_i ));
    InMux I__12106 (
            .O(N__61243),
            .I(N__61237));
    InMux I__12105 (
            .O(N__61242),
            .I(N__61237));
    LocalMux I__12104 (
            .O(N__61237),
            .I(\pid_front.un1_pid_prereg_0_12 ));
    CascadeMux I__12103 (
            .O(N__61234),
            .I(\pid_front.un1_pid_prereg_0_14_cascade_ ));
    CascadeMux I__12102 (
            .O(N__61231),
            .I(N__61228));
    InMux I__12101 (
            .O(N__61228),
            .I(N__61225));
    LocalMux I__12100 (
            .O(N__61225),
            .I(N__61222));
    Span4Mux_v I__12099 (
            .O(N__61222),
            .I(N__61219));
    Odrv4 I__12098 (
            .O(N__61219),
            .I(\pid_front.error_d_reg_prev_esr_RNION3U9Z0Z_21 ));
    InMux I__12097 (
            .O(N__61216),
            .I(N__61207));
    InMux I__12096 (
            .O(N__61215),
            .I(N__61207));
    InMux I__12095 (
            .O(N__61214),
            .I(N__61207));
    LocalMux I__12094 (
            .O(N__61207),
            .I(\pid_front.un1_pid_prereg_0_13 ));
    CascadeMux I__12093 (
            .O(N__61204),
            .I(\pid_front.un1_pid_prereg_0_15_cascade_ ));
    CascadeMux I__12092 (
            .O(N__61201),
            .I(N__61198));
    InMux I__12091 (
            .O(N__61198),
            .I(N__61195));
    LocalMux I__12090 (
            .O(N__61195),
            .I(N__61192));
    Span4Mux_v I__12089 (
            .O(N__61192),
            .I(N__61189));
    Odrv4 I__12088 (
            .O(N__61189),
            .I(\pid_front.error_d_reg_prev_esr_RNIQHRB4Z0Z_21 ));
    CascadeMux I__12087 (
            .O(N__61186),
            .I(N__61183));
    InMux I__12086 (
            .O(N__61183),
            .I(N__61180));
    LocalMux I__12085 (
            .O(N__61180),
            .I(\pid_front.error_p_reg_esr_RNID8DF2Z0Z_3 ));
    CascadeMux I__12084 (
            .O(N__61177),
            .I(N__61174));
    InMux I__12083 (
            .O(N__61174),
            .I(N__61171));
    LocalMux I__12082 (
            .O(N__61171),
            .I(\pid_front.error_p_reg_esr_RNIR7E8Z0Z_3 ));
    CascadeMux I__12081 (
            .O(N__61168),
            .I(\pid_front.error_p_reg_esr_RNIR7E8Z0Z_3_cascade_ ));
    InMux I__12080 (
            .O(N__61165),
            .I(N__61162));
    LocalMux I__12079 (
            .O(N__61162),
            .I(\pid_front.error_p_reg_esr_RNIRJAF2Z0Z_3 ));
    InMux I__12078 (
            .O(N__61159),
            .I(N__61156));
    LocalMux I__12077 (
            .O(N__61156),
            .I(N__61153));
    Span4Mux_v I__12076 (
            .O(N__61153),
            .I(N__61149));
    InMux I__12075 (
            .O(N__61152),
            .I(N__61146));
    Odrv4 I__12074 (
            .O(N__61149),
            .I(\pid_front.error_p_regZ0Z_4 ));
    LocalMux I__12073 (
            .O(N__61146),
            .I(\pid_front.error_p_regZ0Z_4 ));
    InMux I__12072 (
            .O(N__61141),
            .I(N__61135));
    InMux I__12071 (
            .O(N__61140),
            .I(N__61135));
    LocalMux I__12070 (
            .O(N__61135),
            .I(\pid_front.error_p_reg_esr_RNIUAE8_0Z0Z_4 ));
    CascadeMux I__12069 (
            .O(N__61132),
            .I(\pid_front.N_45_i_i_0_cascade_ ));
    CascadeMux I__12068 (
            .O(N__61129),
            .I(\pid_front.error_cry_1_0_c_RNINF5AZ0Z3_cascade_ ));
    CascadeMux I__12067 (
            .O(N__61126),
            .I(\pid_front.un4_error_i_reg_28_ns_1_1_cascade_ ));
    InMux I__12066 (
            .O(N__61123),
            .I(N__61120));
    LocalMux I__12065 (
            .O(N__61120),
            .I(N__61117));
    Span4Mux_h I__12064 (
            .O(N__61117),
            .I(N__61114));
    Odrv4 I__12063 (
            .O(N__61114),
            .I(\pid_front.error_i_reg_9_1_18 ));
    CascadeMux I__12062 (
            .O(N__61111),
            .I(\pid_front.un4_error_i_reg_28_ns_1_cascade_ ));
    InMux I__12061 (
            .O(N__61108),
            .I(N__61105));
    LocalMux I__12060 (
            .O(N__61105),
            .I(\pid_front.m6_2_01 ));
    InMux I__12059 (
            .O(N__61102),
            .I(N__61099));
    LocalMux I__12058 (
            .O(N__61099),
            .I(N__61096));
    Span4Mux_h I__12057 (
            .O(N__61096),
            .I(N__61093));
    Span4Mux_v I__12056 (
            .O(N__61093),
            .I(N__61088));
    InMux I__12055 (
            .O(N__61092),
            .I(N__61083));
    InMux I__12054 (
            .O(N__61091),
            .I(N__61083));
    Odrv4 I__12053 (
            .O(N__61088),
            .I(\pid_front.un1_pid_prereg_0_11 ));
    LocalMux I__12052 (
            .O(N__61083),
            .I(\pid_front.un1_pid_prereg_0_11 ));
    CascadeMux I__12051 (
            .O(N__61078),
            .I(\pid_front.un1_pid_prereg_0_12_cascade_ ));
    InMux I__12050 (
            .O(N__61075),
            .I(N__61072));
    LocalMux I__12049 (
            .O(N__61072),
            .I(N__61069));
    Span4Mux_h I__12048 (
            .O(N__61069),
            .I(N__61066));
    Span4Mux_h I__12047 (
            .O(N__61066),
            .I(N__61062));
    InMux I__12046 (
            .O(N__61065),
            .I(N__61059));
    Odrv4 I__12045 (
            .O(N__61062),
            .I(\pid_front.un1_pid_prereg_0_10 ));
    LocalMux I__12044 (
            .O(N__61059),
            .I(\pid_front.un1_pid_prereg_0_10 ));
    InMux I__12043 (
            .O(N__61054),
            .I(N__61051));
    LocalMux I__12042 (
            .O(N__61051),
            .I(N__61048));
    Span4Mux_v I__12041 (
            .O(N__61048),
            .I(N__61045));
    Odrv4 I__12040 (
            .O(N__61045),
            .I(\pid_front.error_d_reg_prev_esr_RNIV42ACZ0Z_21 ));
    InMux I__12039 (
            .O(N__61042),
            .I(N__61039));
    LocalMux I__12038 (
            .O(N__61039),
            .I(N__61036));
    Span4Mux_v I__12037 (
            .O(N__61036),
            .I(N__61033));
    Odrv4 I__12036 (
            .O(N__61033),
            .I(\pid_front.error_d_reg_prev_esr_RNIU58I5Z0Z_21 ));
    InMux I__12035 (
            .O(N__61030),
            .I(N__61027));
    LocalMux I__12034 (
            .O(N__61027),
            .I(N__61024));
    Span4Mux_v I__12033 (
            .O(N__61024),
            .I(N__61021));
    Odrv4 I__12032 (
            .O(N__61021),
            .I(\pid_front.m27_2_03_0 ));
    InMux I__12031 (
            .O(N__61018),
            .I(N__61015));
    LocalMux I__12030 (
            .O(N__61015),
            .I(N__61011));
    InMux I__12029 (
            .O(N__61014),
            .I(N__61008));
    Odrv12 I__12028 (
            .O(N__61011),
            .I(\pid_front.N_154 ));
    LocalMux I__12027 (
            .O(N__61008),
            .I(\pid_front.N_154 ));
    CascadeMux I__12026 (
            .O(N__61003),
            .I(\pid_front.N_225_cascade_ ));
    CascadeMux I__12025 (
            .O(N__61000),
            .I(\pid_front.N_478_cascade_ ));
    CascadeMux I__12024 (
            .O(N__60997),
            .I(\pid_front.error_i_reg_9_N_5L8_0_1_cascade_ ));
    InMux I__12023 (
            .O(N__60994),
            .I(N__60991));
    LocalMux I__12022 (
            .O(N__60991),
            .I(\pid_front.error_i_reg_esr_RNO_0Z0Z_21 ));
    CascadeMux I__12021 (
            .O(N__60988),
            .I(\pid_front.N_583_cascade_ ));
    InMux I__12020 (
            .O(N__60985),
            .I(N__60982));
    LocalMux I__12019 (
            .O(N__60982),
            .I(\pid_front.N_597 ));
    CascadeMux I__12018 (
            .O(N__60979),
            .I(\pid_front.error_i_reg_esr_RNO_0Z0Z_8_cascade_ ));
    InMux I__12017 (
            .O(N__60976),
            .I(N__60970));
    InMux I__12016 (
            .O(N__60975),
            .I(N__60970));
    LocalMux I__12015 (
            .O(N__60970),
            .I(\pid_front.N_598 ));
    InMux I__12014 (
            .O(N__60967),
            .I(N__60964));
    LocalMux I__12013 (
            .O(N__60964),
            .I(\pid_front.m28_2_03_0 ));
    InMux I__12012 (
            .O(N__60961),
            .I(N__60958));
    LocalMux I__12011 (
            .O(N__60958),
            .I(\pid_front.m28_2_03_0_0 ));
    CascadeMux I__12010 (
            .O(N__60955),
            .I(\pid_front.N_302_cascade_ ));
    CascadeMux I__12009 (
            .O(N__60952),
            .I(\pid_front.error_i_reg_9_rn_2_25_cascade_ ));
    InMux I__12008 (
            .O(N__60949),
            .I(N__60946));
    LocalMux I__12007 (
            .O(N__60946),
            .I(\pid_front.error_i_reg_9_sn_25 ));
    CascadeMux I__12006 (
            .O(N__60943),
            .I(N__60940));
    InMux I__12005 (
            .O(N__60940),
            .I(N__60937));
    LocalMux I__12004 (
            .O(N__60937),
            .I(\pid_front.m9_2_03_3_i_3 ));
    CascadeMux I__12003 (
            .O(N__60934),
            .I(\pid_front.error_cry_1_0_c_RNII2EF1Z0Z_0_cascade_ ));
    InMux I__12002 (
            .O(N__60931),
            .I(N__60928));
    LocalMux I__12001 (
            .O(N__60928),
            .I(\pid_front.N_228 ));
    CascadeMux I__12000 (
            .O(N__60925),
            .I(\pid_front.N_228_cascade_ ));
    InMux I__11999 (
            .O(N__60922),
            .I(N__60919));
    LocalMux I__11998 (
            .O(N__60919),
            .I(\pid_front.error_i_reg_9_sn_26 ));
    InMux I__11997 (
            .O(N__60916),
            .I(N__60913));
    LocalMux I__11996 (
            .O(N__60913),
            .I(\pid_front.error_cry_1_0_c_RNII2EFZ0Z1 ));
    CascadeMux I__11995 (
            .O(N__60910),
            .I(\pid_front.N_182_cascade_ ));
    CascadeMux I__11994 (
            .O(N__60907),
            .I(\pid_front.N_597_cascade_ ));
    CascadeMux I__11993 (
            .O(N__60904),
            .I(\pid_front.m12_2_03_4_i_0_cascade_ ));
    InMux I__11992 (
            .O(N__60901),
            .I(N__60898));
    LocalMux I__11991 (
            .O(N__60898),
            .I(\pid_front.N_583 ));
    InMux I__11990 (
            .O(N__60895),
            .I(N__60892));
    LocalMux I__11989 (
            .O(N__60892),
            .I(N__60889));
    Span4Mux_v I__11988 (
            .O(N__60889),
            .I(N__60886));
    Span4Mux_h I__11987 (
            .O(N__60886),
            .I(N__60883));
    Span4Mux_h I__11986 (
            .O(N__60883),
            .I(N__60880));
    Span4Mux_h I__11985 (
            .O(N__60880),
            .I(N__60877));
    Odrv4 I__11984 (
            .O(N__60877),
            .I(\pid_front.O_0_8 ));
    InMux I__11983 (
            .O(N__60874),
            .I(N__60871));
    LocalMux I__11982 (
            .O(N__60871),
            .I(N__60868));
    Span12Mux_v I__11981 (
            .O(N__60868),
            .I(N__60865));
    Odrv12 I__11980 (
            .O(N__60865),
            .I(\pid_front.O_7 ));
    InMux I__11979 (
            .O(N__60862),
            .I(N__60856));
    InMux I__11978 (
            .O(N__60861),
            .I(N__60856));
    LocalMux I__11977 (
            .O(N__60856),
            .I(N__60853));
    Span4Mux_v I__11976 (
            .O(N__60853),
            .I(N__60850));
    Odrv4 I__11975 (
            .O(N__60850),
            .I(drone_H_disp_side_11));
    CascadeMux I__11974 (
            .O(N__60847),
            .I(\pid_front.N_581_cascade_ ));
    CascadeMux I__11973 (
            .O(N__60844),
            .I(\pid_front.error_i_reg_esr_RNO_0Z0Z_10_cascade_ ));
    InMux I__11972 (
            .O(N__60841),
            .I(N__60838));
    LocalMux I__11971 (
            .O(N__60838),
            .I(\pid_front.N_581 ));
    CascadeMux I__11970 (
            .O(N__60835),
            .I(\pid_side.state_RNIL5IFZ0Z_0_cascade_ ));
    IoInMux I__11969 (
            .O(N__60832),
            .I(N__60829));
    LocalMux I__11968 (
            .O(N__60829),
            .I(N__60826));
    Span4Mux_s1_v I__11967 (
            .O(N__60826),
            .I(N__60823));
    Span4Mux_v I__11966 (
            .O(N__60823),
            .I(N__60820));
    Span4Mux_v I__11965 (
            .O(N__60820),
            .I(N__60817));
    Span4Mux_v I__11964 (
            .O(N__60817),
            .I(N__60814));
    Span4Mux_v I__11963 (
            .O(N__60814),
            .I(N__60811));
    Odrv4 I__11962 (
            .O(N__60811),
            .I(\pid_side.state_RNIIIOOZ0Z_0 ));
    CascadeMux I__11961 (
            .O(N__60808),
            .I(N__60805));
    InMux I__11960 (
            .O(N__60805),
            .I(N__60799));
    InMux I__11959 (
            .O(N__60804),
            .I(N__60799));
    LocalMux I__11958 (
            .O(N__60799),
            .I(N__60795));
    InMux I__11957 (
            .O(N__60798),
            .I(N__60792));
    Span4Mux_h I__11956 (
            .O(N__60795),
            .I(N__60786));
    LocalMux I__11955 (
            .O(N__60792),
            .I(N__60780));
    InMux I__11954 (
            .O(N__60791),
            .I(N__60773));
    InMux I__11953 (
            .O(N__60790),
            .I(N__60773));
    InMux I__11952 (
            .O(N__60789),
            .I(N__60773));
    Span4Mux_v I__11951 (
            .O(N__60786),
            .I(N__60770));
    InMux I__11950 (
            .O(N__60785),
            .I(N__60763));
    InMux I__11949 (
            .O(N__60784),
            .I(N__60763));
    InMux I__11948 (
            .O(N__60783),
            .I(N__60763));
    Odrv4 I__11947 (
            .O(N__60780),
            .I(\pid_side.stateZ0Z_0 ));
    LocalMux I__11946 (
            .O(N__60773),
            .I(\pid_side.stateZ0Z_0 ));
    Odrv4 I__11945 (
            .O(N__60770),
            .I(\pid_side.stateZ0Z_0 ));
    LocalMux I__11944 (
            .O(N__60763),
            .I(\pid_side.stateZ0Z_0 ));
    CascadeMux I__11943 (
            .O(N__60754),
            .I(N__60749));
    CascadeMux I__11942 (
            .O(N__60753),
            .I(N__60740));
    CascadeMux I__11941 (
            .O(N__60752),
            .I(N__60737));
    InMux I__11940 (
            .O(N__60749),
            .I(N__60724));
    InMux I__11939 (
            .O(N__60748),
            .I(N__60724));
    InMux I__11938 (
            .O(N__60747),
            .I(N__60724));
    InMux I__11937 (
            .O(N__60746),
            .I(N__60724));
    InMux I__11936 (
            .O(N__60745),
            .I(N__60724));
    InMux I__11935 (
            .O(N__60744),
            .I(N__60724));
    InMux I__11934 (
            .O(N__60743),
            .I(N__60719));
    InMux I__11933 (
            .O(N__60740),
            .I(N__60719));
    InMux I__11932 (
            .O(N__60737),
            .I(N__60716));
    LocalMux I__11931 (
            .O(N__60724),
            .I(N__60712));
    LocalMux I__11930 (
            .O(N__60719),
            .I(N__60706));
    LocalMux I__11929 (
            .O(N__60716),
            .I(N__60706));
    InMux I__11928 (
            .O(N__60715),
            .I(N__60703));
    Span4Mux_h I__11927 (
            .O(N__60712),
            .I(N__60700));
    InMux I__11926 (
            .O(N__60711),
            .I(N__60695));
    Span4Mux_v I__11925 (
            .O(N__60706),
            .I(N__60692));
    LocalMux I__11924 (
            .O(N__60703),
            .I(N__60688));
    Span4Mux_v I__11923 (
            .O(N__60700),
            .I(N__60685));
    InMux I__11922 (
            .O(N__60699),
            .I(N__60680));
    InMux I__11921 (
            .O(N__60698),
            .I(N__60680));
    LocalMux I__11920 (
            .O(N__60695),
            .I(N__60677));
    Span4Mux_v I__11919 (
            .O(N__60692),
            .I(N__60674));
    InMux I__11918 (
            .O(N__60691),
            .I(N__60671));
    Span4Mux_h I__11917 (
            .O(N__60688),
            .I(N__60668));
    Odrv4 I__11916 (
            .O(N__60685),
            .I(\pid_side.stateZ0Z_1 ));
    LocalMux I__11915 (
            .O(N__60680),
            .I(\pid_side.stateZ0Z_1 ));
    Odrv12 I__11914 (
            .O(N__60677),
            .I(\pid_side.stateZ0Z_1 ));
    Odrv4 I__11913 (
            .O(N__60674),
            .I(\pid_side.stateZ0Z_1 ));
    LocalMux I__11912 (
            .O(N__60671),
            .I(\pid_side.stateZ0Z_1 ));
    Odrv4 I__11911 (
            .O(N__60668),
            .I(\pid_side.stateZ0Z_1 ));
    CascadeMux I__11910 (
            .O(N__60655),
            .I(\pid_front.state_ns_0_cascade_ ));
    InMux I__11909 (
            .O(N__60652),
            .I(N__60649));
    LocalMux I__11908 (
            .O(N__60649),
            .I(N__60646));
    Span4Mux_h I__11907 (
            .O(N__60646),
            .I(N__60643));
    Odrv4 I__11906 (
            .O(N__60643),
            .I(\pid_front.N_536_1 ));
    InMux I__11905 (
            .O(N__60640),
            .I(N__60637));
    LocalMux I__11904 (
            .O(N__60637),
            .I(\pid_front.N_297 ));
    InMux I__11903 (
            .O(N__60634),
            .I(N__60631));
    LocalMux I__11902 (
            .O(N__60631),
            .I(N__60628));
    Span12Mux_v I__11901 (
            .O(N__60628),
            .I(N__60625));
    Span12Mux_h I__11900 (
            .O(N__60625),
            .I(N__60622));
    Odrv12 I__11899 (
            .O(N__60622),
            .I(\pid_front.O_0_22 ));
    InMux I__11898 (
            .O(N__60619),
            .I(N__60613));
    InMux I__11897 (
            .O(N__60618),
            .I(N__60613));
    LocalMux I__11896 (
            .O(N__60613),
            .I(\pid_side.error_i_acumm_preregZ0Z_13 ));
    InMux I__11895 (
            .O(N__60610),
            .I(N__60607));
    LocalMux I__11894 (
            .O(N__60607),
            .I(N__60604));
    Span4Mux_s3_v I__11893 (
            .O(N__60604),
            .I(N__60601));
    Span4Mux_v I__11892 (
            .O(N__60601),
            .I(N__60598));
    Odrv4 I__11891 (
            .O(N__60598),
            .I(\pid_side.error_i_acumm_13_i_o2_0_10_3 ));
    InMux I__11890 (
            .O(N__60595),
            .I(N__60589));
    InMux I__11889 (
            .O(N__60594),
            .I(N__60589));
    LocalMux I__11888 (
            .O(N__60589),
            .I(\pid_side.error_i_acumm_preregZ0Z_18 ));
    InMux I__11887 (
            .O(N__60586),
            .I(N__60580));
    InMux I__11886 (
            .O(N__60585),
            .I(N__60580));
    LocalMux I__11885 (
            .O(N__60580),
            .I(\pid_side.error_i_acumm_preregZ0Z_25 ));
    CascadeMux I__11884 (
            .O(N__60577),
            .I(N__60573));
    CascadeMux I__11883 (
            .O(N__60576),
            .I(N__60570));
    InMux I__11882 (
            .O(N__60573),
            .I(N__60565));
    InMux I__11881 (
            .O(N__60570),
            .I(N__60565));
    LocalMux I__11880 (
            .O(N__60565),
            .I(\pid_side.error_i_acumm_preregZ0Z_26 ));
    InMux I__11879 (
            .O(N__60562),
            .I(N__60559));
    LocalMux I__11878 (
            .O(N__60559),
            .I(\pid_side.N_338 ));
    CascadeMux I__11877 (
            .O(N__60556),
            .I(pid_side_N_382_4_cascade_));
    CascadeMux I__11876 (
            .O(N__60553),
            .I(\pid_side.N_382_cascade_ ));
    CEMux I__11875 (
            .O(N__60550),
            .I(N__60545));
    CEMux I__11874 (
            .O(N__60549),
            .I(N__60542));
    CEMux I__11873 (
            .O(N__60548),
            .I(N__60538));
    LocalMux I__11872 (
            .O(N__60545),
            .I(N__60533));
    LocalMux I__11871 (
            .O(N__60542),
            .I(N__60530));
    CEMux I__11870 (
            .O(N__60541),
            .I(N__60527));
    LocalMux I__11869 (
            .O(N__60538),
            .I(N__60524));
    CEMux I__11868 (
            .O(N__60537),
            .I(N__60521));
    CEMux I__11867 (
            .O(N__60536),
            .I(N__60518));
    Span4Mux_v I__11866 (
            .O(N__60533),
            .I(N__60511));
    Span4Mux_h I__11865 (
            .O(N__60530),
            .I(N__60511));
    LocalMux I__11864 (
            .O(N__60527),
            .I(N__60511));
    Span4Mux_v I__11863 (
            .O(N__60524),
            .I(N__60508));
    LocalMux I__11862 (
            .O(N__60521),
            .I(N__60503));
    LocalMux I__11861 (
            .O(N__60518),
            .I(N__60503));
    Span4Mux_h I__11860 (
            .O(N__60511),
            .I(N__60500));
    Span4Mux_h I__11859 (
            .O(N__60508),
            .I(N__60497));
    Sp12to4 I__11858 (
            .O(N__60503),
            .I(N__60494));
    Span4Mux_h I__11857 (
            .O(N__60500),
            .I(N__60491));
    Odrv4 I__11856 (
            .O(N__60497),
            .I(\pid_side.N_64 ));
    Odrv12 I__11855 (
            .O(N__60494),
            .I(\pid_side.N_64 ));
    Odrv4 I__11854 (
            .O(N__60491),
            .I(\pid_side.N_64 ));
    CascadeMux I__11853 (
            .O(N__60484),
            .I(\pid_side.un1_pid_prereg_0_20_cascade_ ));
    CascadeMux I__11852 (
            .O(N__60481),
            .I(\pid_side.un1_pid_prereg_0_22_cascade_ ));
    InMux I__11851 (
            .O(N__60478),
            .I(N__60472));
    InMux I__11850 (
            .O(N__60477),
            .I(N__60472));
    LocalMux I__11849 (
            .O(N__60472),
            .I(\pid_side.un1_pid_prereg_0_20 ));
    InMux I__11848 (
            .O(N__60469),
            .I(N__60464));
    InMux I__11847 (
            .O(N__60468),
            .I(N__60459));
    InMux I__11846 (
            .O(N__60467),
            .I(N__60459));
    LocalMux I__11845 (
            .O(N__60464),
            .I(\pid_side.un1_pid_prereg_0_21 ));
    LocalMux I__11844 (
            .O(N__60459),
            .I(\pid_side.un1_pid_prereg_0_21 ));
    InMux I__11843 (
            .O(N__60454),
            .I(N__60446));
    InMux I__11842 (
            .O(N__60453),
            .I(N__60439));
    InMux I__11841 (
            .O(N__60452),
            .I(N__60434));
    InMux I__11840 (
            .O(N__60451),
            .I(N__60434));
    InMux I__11839 (
            .O(N__60450),
            .I(N__60431));
    InMux I__11838 (
            .O(N__60449),
            .I(N__60427));
    LocalMux I__11837 (
            .O(N__60446),
            .I(N__60424));
    InMux I__11836 (
            .O(N__60445),
            .I(N__60421));
    InMux I__11835 (
            .O(N__60444),
            .I(N__60416));
    InMux I__11834 (
            .O(N__60443),
            .I(N__60416));
    InMux I__11833 (
            .O(N__60442),
            .I(N__60413));
    LocalMux I__11832 (
            .O(N__60439),
            .I(N__60406));
    LocalMux I__11831 (
            .O(N__60434),
            .I(N__60406));
    LocalMux I__11830 (
            .O(N__60431),
            .I(N__60406));
    InMux I__11829 (
            .O(N__60430),
            .I(N__60403));
    LocalMux I__11828 (
            .O(N__60427),
            .I(N__60400));
    Span4Mux_v I__11827 (
            .O(N__60424),
            .I(N__60397));
    LocalMux I__11826 (
            .O(N__60421),
            .I(N__60394));
    LocalMux I__11825 (
            .O(N__60416),
            .I(N__60391));
    LocalMux I__11824 (
            .O(N__60413),
            .I(N__60388));
    Span4Mux_h I__11823 (
            .O(N__60406),
            .I(N__60385));
    LocalMux I__11822 (
            .O(N__60403),
            .I(N__60380));
    Span4Mux_h I__11821 (
            .O(N__60400),
            .I(N__60380));
    Span4Mux_h I__11820 (
            .O(N__60397),
            .I(N__60377));
    Span4Mux_v I__11819 (
            .O(N__60394),
            .I(N__60374));
    Span4Mux_v I__11818 (
            .O(N__60391),
            .I(N__60367));
    Span4Mux_v I__11817 (
            .O(N__60388),
            .I(N__60367));
    Span4Mux_v I__11816 (
            .O(N__60385),
            .I(N__60367));
    Span4Mux_v I__11815 (
            .O(N__60380),
            .I(N__60364));
    Odrv4 I__11814 (
            .O(N__60377),
            .I(\pid_side.N_205 ));
    Odrv4 I__11813 (
            .O(N__60374),
            .I(\pid_side.N_205 ));
    Odrv4 I__11812 (
            .O(N__60367),
            .I(\pid_side.N_205 ));
    Odrv4 I__11811 (
            .O(N__60364),
            .I(\pid_side.N_205 ));
    InMux I__11810 (
            .O(N__60355),
            .I(N__60346));
    InMux I__11809 (
            .O(N__60354),
            .I(N__60346));
    InMux I__11808 (
            .O(N__60353),
            .I(N__60346));
    LocalMux I__11807 (
            .O(N__60346),
            .I(N__60343));
    Span4Mux_v I__11806 (
            .O(N__60343),
            .I(N__60340));
    Odrv4 I__11805 (
            .O(N__60340),
            .I(\pid_side.N_285 ));
    CascadeMux I__11804 (
            .O(N__60337),
            .I(\pid_side.N_353_cascade_ ));
    InMux I__11803 (
            .O(N__60334),
            .I(N__60327));
    InMux I__11802 (
            .O(N__60333),
            .I(N__60327));
    CascadeMux I__11801 (
            .O(N__60332),
            .I(N__60323));
    LocalMux I__11800 (
            .O(N__60327),
            .I(N__60318));
    InMux I__11799 (
            .O(N__60326),
            .I(N__60315));
    InMux I__11798 (
            .O(N__60323),
            .I(N__60310));
    InMux I__11797 (
            .O(N__60322),
            .I(N__60310));
    InMux I__11796 (
            .O(N__60321),
            .I(N__60307));
    Odrv4 I__11795 (
            .O(N__60318),
            .I(\pid_side.error_i_acumm_preregZ0Z_11 ));
    LocalMux I__11794 (
            .O(N__60315),
            .I(\pid_side.error_i_acumm_preregZ0Z_11 ));
    LocalMux I__11793 (
            .O(N__60310),
            .I(\pid_side.error_i_acumm_preregZ0Z_11 ));
    LocalMux I__11792 (
            .O(N__60307),
            .I(\pid_side.error_i_acumm_preregZ0Z_11 ));
    InMux I__11791 (
            .O(N__60298),
            .I(N__60295));
    LocalMux I__11790 (
            .O(N__60295),
            .I(N__60292));
    Span4Mux_v I__11789 (
            .O(N__60292),
            .I(N__60289));
    Span4Mux_v I__11788 (
            .O(N__60289),
            .I(N__60286));
    Span4Mux_v I__11787 (
            .O(N__60286),
            .I(N__60281));
    InMux I__11786 (
            .O(N__60285),
            .I(N__60276));
    InMux I__11785 (
            .O(N__60284),
            .I(N__60276));
    Odrv4 I__11784 (
            .O(N__60281),
            .I(\pid_front.pid_preregZ0Z_0 ));
    LocalMux I__11783 (
            .O(N__60276),
            .I(\pid_front.pid_preregZ0Z_0 ));
    InMux I__11782 (
            .O(N__60271),
            .I(N__60268));
    LocalMux I__11781 (
            .O(N__60268),
            .I(N__60264));
    InMux I__11780 (
            .O(N__60267),
            .I(N__60261));
    Span4Mux_v I__11779 (
            .O(N__60264),
            .I(N__60256));
    LocalMux I__11778 (
            .O(N__60261),
            .I(N__60256));
    Span4Mux_h I__11777 (
            .O(N__60256),
            .I(N__60253));
    Odrv4 I__11776 (
            .O(N__60253),
            .I(front_order_0));
    InMux I__11775 (
            .O(N__60250),
            .I(N__60247));
    LocalMux I__11774 (
            .O(N__60247),
            .I(N__60244));
    Span12Mux_h I__11773 (
            .O(N__60244),
            .I(N__60241));
    Span12Mux_v I__11772 (
            .O(N__60241),
            .I(N__60236));
    InMux I__11771 (
            .O(N__60240),
            .I(N__60231));
    InMux I__11770 (
            .O(N__60239),
            .I(N__60231));
    Odrv12 I__11769 (
            .O(N__60236),
            .I(\pid_front.pid_preregZ0Z_2 ));
    LocalMux I__11768 (
            .O(N__60231),
            .I(\pid_front.pid_preregZ0Z_2 ));
    InMux I__11767 (
            .O(N__60226),
            .I(N__60223));
    LocalMux I__11766 (
            .O(N__60223),
            .I(N__60220));
    Span4Mux_v I__11765 (
            .O(N__60220),
            .I(N__60216));
    InMux I__11764 (
            .O(N__60219),
            .I(N__60213));
    Span4Mux_h I__11763 (
            .O(N__60216),
            .I(N__60210));
    LocalMux I__11762 (
            .O(N__60213),
            .I(N__60207));
    Span4Mux_h I__11761 (
            .O(N__60210),
            .I(N__60204));
    Span4Mux_h I__11760 (
            .O(N__60207),
            .I(N__60201));
    Odrv4 I__11759 (
            .O(N__60204),
            .I(front_order_2));
    Odrv4 I__11758 (
            .O(N__60201),
            .I(front_order_2));
    InMux I__11757 (
            .O(N__60196),
            .I(N__60187));
    InMux I__11756 (
            .O(N__60195),
            .I(N__60187));
    InMux I__11755 (
            .O(N__60194),
            .I(N__60187));
    LocalMux I__11754 (
            .O(N__60187),
            .I(N__60176));
    InMux I__11753 (
            .O(N__60186),
            .I(N__60163));
    InMux I__11752 (
            .O(N__60185),
            .I(N__60163));
    InMux I__11751 (
            .O(N__60184),
            .I(N__60163));
    InMux I__11750 (
            .O(N__60183),
            .I(N__60163));
    InMux I__11749 (
            .O(N__60182),
            .I(N__60163));
    InMux I__11748 (
            .O(N__60181),
            .I(N__60163));
    InMux I__11747 (
            .O(N__60180),
            .I(N__60158));
    InMux I__11746 (
            .O(N__60179),
            .I(N__60158));
    Span12Mux_s11_v I__11745 (
            .O(N__60176),
            .I(N__60155));
    LocalMux I__11744 (
            .O(N__60163),
            .I(N__60150));
    LocalMux I__11743 (
            .O(N__60158),
            .I(N__60150));
    Span12Mux_v I__11742 (
            .O(N__60155),
            .I(N__60146));
    Span12Mux_v I__11741 (
            .O(N__60150),
            .I(N__60143));
    InMux I__11740 (
            .O(N__60149),
            .I(N__60140));
    Odrv12 I__11739 (
            .O(N__60146),
            .I(\pid_front.N_386 ));
    Odrv12 I__11738 (
            .O(N__60143),
            .I(\pid_front.N_386 ));
    LocalMux I__11737 (
            .O(N__60140),
            .I(\pid_front.N_386 ));
    InMux I__11736 (
            .O(N__60133),
            .I(N__60124));
    InMux I__11735 (
            .O(N__60132),
            .I(N__60124));
    InMux I__11734 (
            .O(N__60131),
            .I(N__60124));
    LocalMux I__11733 (
            .O(N__60124),
            .I(N__60119));
    InMux I__11732 (
            .O(N__60123),
            .I(N__60114));
    InMux I__11731 (
            .O(N__60122),
            .I(N__60114));
    Span4Mux_v I__11730 (
            .O(N__60119),
            .I(N__60109));
    LocalMux I__11729 (
            .O(N__60114),
            .I(N__60109));
    Span4Mux_h I__11728 (
            .O(N__60109),
            .I(N__60105));
    InMux I__11727 (
            .O(N__60108),
            .I(N__60102));
    Sp12to4 I__11726 (
            .O(N__60105),
            .I(N__60099));
    LocalMux I__11725 (
            .O(N__60102),
            .I(N__60096));
    Odrv12 I__11724 (
            .O(N__60099),
            .I(\pid_front.N_631 ));
    Odrv4 I__11723 (
            .O(N__60096),
            .I(\pid_front.N_631 ));
    InMux I__11722 (
            .O(N__60091),
            .I(N__60088));
    LocalMux I__11721 (
            .O(N__60088),
            .I(N__60085));
    Span4Mux_v I__11720 (
            .O(N__60085),
            .I(N__60082));
    Span4Mux_v I__11719 (
            .O(N__60082),
            .I(N__60078));
    CascadeMux I__11718 (
            .O(N__60081),
            .I(N__60074));
    Span4Mux_v I__11717 (
            .O(N__60078),
            .I(N__60071));
    InMux I__11716 (
            .O(N__60077),
            .I(N__60066));
    InMux I__11715 (
            .O(N__60074),
            .I(N__60066));
    Odrv4 I__11714 (
            .O(N__60071),
            .I(\pid_front.pid_preregZ0Z_3 ));
    LocalMux I__11713 (
            .O(N__60066),
            .I(\pid_front.pid_preregZ0Z_3 ));
    InMux I__11712 (
            .O(N__60061),
            .I(N__60058));
    LocalMux I__11711 (
            .O(N__60058),
            .I(N__60054));
    InMux I__11710 (
            .O(N__60057),
            .I(N__60051));
    Span4Mux_h I__11709 (
            .O(N__60054),
            .I(N__60046));
    LocalMux I__11708 (
            .O(N__60051),
            .I(N__60046));
    Span4Mux_h I__11707 (
            .O(N__60046),
            .I(N__60043));
    Odrv4 I__11706 (
            .O(N__60043),
            .I(front_order_3));
    CEMux I__11705 (
            .O(N__60040),
            .I(N__60037));
    LocalMux I__11704 (
            .O(N__60037),
            .I(N__60033));
    CEMux I__11703 (
            .O(N__60036),
            .I(N__60030));
    Span4Mux_h I__11702 (
            .O(N__60033),
            .I(N__60024));
    LocalMux I__11701 (
            .O(N__60030),
            .I(N__60024));
    CEMux I__11700 (
            .O(N__60029),
            .I(N__60021));
    Span4Mux_v I__11699 (
            .O(N__60024),
            .I(N__60017));
    LocalMux I__11698 (
            .O(N__60021),
            .I(N__60014));
    CEMux I__11697 (
            .O(N__60020),
            .I(N__60011));
    Span4Mux_v I__11696 (
            .O(N__60017),
            .I(N__60008));
    Span4Mux_h I__11695 (
            .O(N__60014),
            .I(N__60005));
    LocalMux I__11694 (
            .O(N__60011),
            .I(N__60002));
    Odrv4 I__11693 (
            .O(N__60008),
            .I(\pid_front.state_0_1 ));
    Odrv4 I__11692 (
            .O(N__60005),
            .I(\pid_front.state_0_1 ));
    Odrv4 I__11691 (
            .O(N__60002),
            .I(\pid_front.state_0_1 ));
    SRMux I__11690 (
            .O(N__59995),
            .I(N__59992));
    LocalMux I__11689 (
            .O(N__59992),
            .I(N__59987));
    SRMux I__11688 (
            .O(N__59991),
            .I(N__59984));
    SRMux I__11687 (
            .O(N__59990),
            .I(N__59981));
    Span4Mux_h I__11686 (
            .O(N__59987),
            .I(N__59978));
    LocalMux I__11685 (
            .O(N__59984),
            .I(N__59975));
    LocalMux I__11684 (
            .O(N__59981),
            .I(N__59972));
    Span4Mux_v I__11683 (
            .O(N__59978),
            .I(N__59968));
    Span4Mux_v I__11682 (
            .O(N__59975),
            .I(N__59963));
    Span4Mux_v I__11681 (
            .O(N__59972),
            .I(N__59963));
    SRMux I__11680 (
            .O(N__59971),
            .I(N__59960));
    Span4Mux_v I__11679 (
            .O(N__59968),
            .I(N__59957));
    Span4Mux_v I__11678 (
            .O(N__59963),
            .I(N__59954));
    LocalMux I__11677 (
            .O(N__59960),
            .I(N__59951));
    Span4Mux_h I__11676 (
            .O(N__59957),
            .I(N__59947));
    Span4Mux_v I__11675 (
            .O(N__59954),
            .I(N__59942));
    Span4Mux_h I__11674 (
            .O(N__59951),
            .I(N__59942));
    SRMux I__11673 (
            .O(N__59950),
            .I(N__59939));
    Odrv4 I__11672 (
            .O(N__59947),
            .I(\pid_front.un1_reset_0_i_3 ));
    Odrv4 I__11671 (
            .O(N__59942),
            .I(\pid_front.un1_reset_0_i_3 ));
    LocalMux I__11670 (
            .O(N__59939),
            .I(\pid_front.un1_reset_0_i_3 ));
    CascadeMux I__11669 (
            .O(N__59932),
            .I(\pid_side.error_d_reg_prev_esr_RNI5RIOZ0Z_14_cascade_ ));
    CascadeMux I__11668 (
            .O(N__59929),
            .I(\pid_side.N_488_cascade_ ));
    CascadeMux I__11667 (
            .O(N__59926),
            .I(N__59923));
    InMux I__11666 (
            .O(N__59923),
            .I(N__59917));
    InMux I__11665 (
            .O(N__59922),
            .I(N__59917));
    LocalMux I__11664 (
            .O(N__59917),
            .I(N__59912));
    InMux I__11663 (
            .O(N__59916),
            .I(N__59907));
    InMux I__11662 (
            .O(N__59915),
            .I(N__59907));
    Odrv4 I__11661 (
            .O(N__59912),
            .I(\pid_side.N_601 ));
    LocalMux I__11660 (
            .O(N__59907),
            .I(\pid_side.N_601 ));
    CascadeMux I__11659 (
            .O(N__59902),
            .I(\pid_side.N_601_cascade_ ));
    InMux I__11658 (
            .O(N__59899),
            .I(N__59896));
    LocalMux I__11657 (
            .O(N__59896),
            .I(N__59893));
    Span4Mux_h I__11656 (
            .O(N__59893),
            .I(N__59890));
    Span4Mux_h I__11655 (
            .O(N__59890),
            .I(N__59887));
    Span4Mux_v I__11654 (
            .O(N__59887),
            .I(N__59884));
    Odrv4 I__11653 (
            .O(N__59884),
            .I(\pid_side.error_i_acumm_preregZ0Z_0 ));
    CascadeMux I__11652 (
            .O(N__59881),
            .I(\pid_side.N_484_cascade_ ));
    InMux I__11651 (
            .O(N__59878),
            .I(N__59872));
    InMux I__11650 (
            .O(N__59877),
            .I(N__59872));
    LocalMux I__11649 (
            .O(N__59872),
            .I(\pid_side.N_484 ));
    InMux I__11648 (
            .O(N__59869),
            .I(N__59866));
    LocalMux I__11647 (
            .O(N__59866),
            .I(N__59863));
    Odrv12 I__11646 (
            .O(N__59863),
            .I(\pid_side.error_i_acumm_preregZ0Z_2 ));
    CascadeMux I__11645 (
            .O(N__59860),
            .I(N__59857));
    InMux I__11644 (
            .O(N__59857),
            .I(N__59848));
    InMux I__11643 (
            .O(N__59856),
            .I(N__59848));
    InMux I__11642 (
            .O(N__59855),
            .I(N__59848));
    LocalMux I__11641 (
            .O(N__59848),
            .I(\pid_side.error_i_acumm_13_0_tz_0_0 ));
    InMux I__11640 (
            .O(N__59845),
            .I(N__59838));
    InMux I__11639 (
            .O(N__59844),
            .I(N__59838));
    InMux I__11638 (
            .O(N__59843),
            .I(N__59835));
    LocalMux I__11637 (
            .O(N__59838),
            .I(N__59830));
    LocalMux I__11636 (
            .O(N__59835),
            .I(N__59830));
    Span4Mux_h I__11635 (
            .O(N__59830),
            .I(N__59827));
    Odrv4 I__11634 (
            .O(N__59827),
            .I(\pid_side.N_634 ));
    InMux I__11633 (
            .O(N__59824),
            .I(N__59818));
    InMux I__11632 (
            .O(N__59823),
            .I(N__59818));
    LocalMux I__11631 (
            .O(N__59818),
            .I(N__59811));
    InMux I__11630 (
            .O(N__59817),
            .I(N__59808));
    InMux I__11629 (
            .O(N__59816),
            .I(N__59803));
    InMux I__11628 (
            .O(N__59815),
            .I(N__59803));
    InMux I__11627 (
            .O(N__59814),
            .I(N__59800));
    Odrv4 I__11626 (
            .O(N__59811),
            .I(\pid_side.error_i_acumm_preregZ0Z_10 ));
    LocalMux I__11625 (
            .O(N__59808),
            .I(\pid_side.error_i_acumm_preregZ0Z_10 ));
    LocalMux I__11624 (
            .O(N__59803),
            .I(\pid_side.error_i_acumm_preregZ0Z_10 ));
    LocalMux I__11623 (
            .O(N__59800),
            .I(\pid_side.error_i_acumm_preregZ0Z_10 ));
    CascadeMux I__11622 (
            .O(N__59791),
            .I(\pid_side.N_355_cascade_ ));
    CascadeMux I__11621 (
            .O(N__59788),
            .I(\pid_side.N_242_cascade_ ));
    InMux I__11620 (
            .O(N__59785),
            .I(N__59778));
    InMux I__11619 (
            .O(N__59784),
            .I(N__59773));
    InMux I__11618 (
            .O(N__59783),
            .I(N__59773));
    InMux I__11617 (
            .O(N__59782),
            .I(N__59770));
    CascadeMux I__11616 (
            .O(N__59781),
            .I(N__59764));
    LocalMux I__11615 (
            .O(N__59778),
            .I(N__59759));
    LocalMux I__11614 (
            .O(N__59773),
            .I(N__59759));
    LocalMux I__11613 (
            .O(N__59770),
            .I(N__59756));
    InMux I__11612 (
            .O(N__59769),
            .I(N__59753));
    CascadeMux I__11611 (
            .O(N__59768),
            .I(N__59749));
    InMux I__11610 (
            .O(N__59767),
            .I(N__59746));
    InMux I__11609 (
            .O(N__59764),
            .I(N__59743));
    Span4Mux_v I__11608 (
            .O(N__59759),
            .I(N__59736));
    Span4Mux_s3_v I__11607 (
            .O(N__59756),
            .I(N__59736));
    LocalMux I__11606 (
            .O(N__59753),
            .I(N__59736));
    InMux I__11605 (
            .O(N__59752),
            .I(N__59733));
    InMux I__11604 (
            .O(N__59749),
            .I(N__59730));
    LocalMux I__11603 (
            .O(N__59746),
            .I(\pid_side.un10lto12 ));
    LocalMux I__11602 (
            .O(N__59743),
            .I(\pid_side.un10lto12 ));
    Odrv4 I__11601 (
            .O(N__59736),
            .I(\pid_side.un10lto12 ));
    LocalMux I__11600 (
            .O(N__59733),
            .I(\pid_side.un10lto12 ));
    LocalMux I__11599 (
            .O(N__59730),
            .I(\pid_side.un10lto12 ));
    InMux I__11598 (
            .O(N__59719),
            .I(N__59708));
    InMux I__11597 (
            .O(N__59718),
            .I(N__59708));
    InMux I__11596 (
            .O(N__59717),
            .I(N__59708));
    InMux I__11595 (
            .O(N__59716),
            .I(N__59705));
    InMux I__11594 (
            .O(N__59715),
            .I(N__59702));
    LocalMux I__11593 (
            .O(N__59708),
            .I(N__59694));
    LocalMux I__11592 (
            .O(N__59705),
            .I(N__59694));
    LocalMux I__11591 (
            .O(N__59702),
            .I(N__59691));
    InMux I__11590 (
            .O(N__59701),
            .I(N__59688));
    InMux I__11589 (
            .O(N__59700),
            .I(N__59683));
    InMux I__11588 (
            .O(N__59699),
            .I(N__59683));
    Span4Mux_v I__11587 (
            .O(N__59694),
            .I(N__59680));
    Sp12to4 I__11586 (
            .O(N__59691),
            .I(N__59673));
    LocalMux I__11585 (
            .O(N__59688),
            .I(N__59673));
    LocalMux I__11584 (
            .O(N__59683),
            .I(N__59673));
    Odrv4 I__11583 (
            .O(N__59680),
            .I(\pid_side.N_227 ));
    Odrv12 I__11582 (
            .O(N__59673),
            .I(\pid_side.N_227 ));
    InMux I__11581 (
            .O(N__59668),
            .I(N__59661));
    InMux I__11580 (
            .O(N__59667),
            .I(N__59661));
    InMux I__11579 (
            .O(N__59666),
            .I(N__59658));
    LocalMux I__11578 (
            .O(N__59661),
            .I(N__59655));
    LocalMux I__11577 (
            .O(N__59658),
            .I(N__59652));
    Span4Mux_v I__11576 (
            .O(N__59655),
            .I(N__59646));
    Span4Mux_h I__11575 (
            .O(N__59652),
            .I(N__59646));
    InMux I__11574 (
            .O(N__59651),
            .I(N__59643));
    Odrv4 I__11573 (
            .O(N__59646),
            .I(\pid_side.error_i_acumm16lto3 ));
    LocalMux I__11572 (
            .O(N__59643),
            .I(\pid_side.error_i_acumm16lto3 ));
    InMux I__11571 (
            .O(N__59638),
            .I(N__59633));
    InMux I__11570 (
            .O(N__59637),
            .I(N__59630));
    InMux I__11569 (
            .O(N__59636),
            .I(N__59627));
    LocalMux I__11568 (
            .O(N__59633),
            .I(\pid_side.error_i_acumm_preregZ0Z_5 ));
    LocalMux I__11567 (
            .O(N__59630),
            .I(\pid_side.error_i_acumm_preregZ0Z_5 ));
    LocalMux I__11566 (
            .O(N__59627),
            .I(\pid_side.error_i_acumm_preregZ0Z_5 ));
    CascadeMux I__11565 (
            .O(N__59620),
            .I(N__59615));
    InMux I__11564 (
            .O(N__59619),
            .I(N__59612));
    InMux I__11563 (
            .O(N__59618),
            .I(N__59607));
    InMux I__11562 (
            .O(N__59615),
            .I(N__59607));
    LocalMux I__11561 (
            .O(N__59612),
            .I(\pid_side.error_i_acumm_preregZ0Z_6 ));
    LocalMux I__11560 (
            .O(N__59607),
            .I(\pid_side.error_i_acumm_preregZ0Z_6 ));
    InMux I__11559 (
            .O(N__59602),
            .I(N__59597));
    InMux I__11558 (
            .O(N__59601),
            .I(N__59591));
    InMux I__11557 (
            .O(N__59600),
            .I(N__59591));
    LocalMux I__11556 (
            .O(N__59597),
            .I(N__59588));
    InMux I__11555 (
            .O(N__59596),
            .I(N__59585));
    LocalMux I__11554 (
            .O(N__59591),
            .I(N__59582));
    Span4Mux_v I__11553 (
            .O(N__59588),
            .I(N__59579));
    LocalMux I__11552 (
            .O(N__59585),
            .I(N__59576));
    Odrv4 I__11551 (
            .O(N__59582),
            .I(\pid_side.error_i_acumm_preregZ0Z_4 ));
    Odrv4 I__11550 (
            .O(N__59579),
            .I(\pid_side.error_i_acumm_preregZ0Z_4 ));
    Odrv12 I__11549 (
            .O(N__59576),
            .I(\pid_side.error_i_acumm_preregZ0Z_4 ));
    CascadeMux I__11548 (
            .O(N__59569),
            .I(\pid_side.error_i_acumm_13_0_a2_2_2_2_cascade_ ));
    CascadeMux I__11547 (
            .O(N__59566),
            .I(N__59563));
    InMux I__11546 (
            .O(N__59563),
            .I(N__59556));
    InMux I__11545 (
            .O(N__59562),
            .I(N__59556));
    InMux I__11544 (
            .O(N__59561),
            .I(N__59553));
    LocalMux I__11543 (
            .O(N__59556),
            .I(N__59550));
    LocalMux I__11542 (
            .O(N__59553),
            .I(\pid_side.N_255 ));
    Odrv12 I__11541 (
            .O(N__59550),
            .I(\pid_side.N_255 ));
    InMux I__11540 (
            .O(N__59545),
            .I(N__59539));
    InMux I__11539 (
            .O(N__59544),
            .I(N__59539));
    LocalMux I__11538 (
            .O(N__59539),
            .I(N__59535));
    InMux I__11537 (
            .O(N__59538),
            .I(N__59532));
    Odrv4 I__11536 (
            .O(N__59535),
            .I(\pid_side.error_i_acumm_13_i_0_tz_7 ));
    LocalMux I__11535 (
            .O(N__59532),
            .I(\pid_side.error_i_acumm_13_i_0_tz_7 ));
    CascadeMux I__11534 (
            .O(N__59527),
            .I(N__59524));
    InMux I__11533 (
            .O(N__59524),
            .I(N__59521));
    LocalMux I__11532 (
            .O(N__59521),
            .I(N__59518));
    Odrv12 I__11531 (
            .O(N__59518),
            .I(\pid_side.error_i_acumm_preregZ0Z_1 ));
    InMux I__11530 (
            .O(N__59515),
            .I(N__59512));
    LocalMux I__11529 (
            .O(N__59512),
            .I(\pid_side.N_181 ));
    CascadeMux I__11528 (
            .O(N__59509),
            .I(\pid_side.N_483_cascade_ ));
    InMux I__11527 (
            .O(N__59506),
            .I(N__59503));
    LocalMux I__11526 (
            .O(N__59503),
            .I(\pid_side.error_i_acumm_13_0_a2_2_4_2 ));
    InMux I__11525 (
            .O(N__59500),
            .I(N__59496));
    InMux I__11524 (
            .O(N__59499),
            .I(N__59493));
    LocalMux I__11523 (
            .O(N__59496),
            .I(N__59487));
    LocalMux I__11522 (
            .O(N__59493),
            .I(N__59487));
    InMux I__11521 (
            .O(N__59492),
            .I(N__59484));
    Odrv4 I__11520 (
            .O(N__59487),
            .I(\pid_side.error_i_acumm_preregZ0Z_9 ));
    LocalMux I__11519 (
            .O(N__59484),
            .I(\pid_side.error_i_acumm_preregZ0Z_9 ));
    InMux I__11518 (
            .O(N__59479),
            .I(N__59476));
    LocalMux I__11517 (
            .O(N__59476),
            .I(N__59472));
    InMux I__11516 (
            .O(N__59475),
            .I(N__59469));
    Span4Mux_v I__11515 (
            .O(N__59472),
            .I(N__59465));
    LocalMux I__11514 (
            .O(N__59469),
            .I(N__59462));
    InMux I__11513 (
            .O(N__59468),
            .I(N__59459));
    Odrv4 I__11512 (
            .O(N__59465),
            .I(\pid_side.error_i_acumm_preregZ0Z_8 ));
    Odrv4 I__11511 (
            .O(N__59462),
            .I(\pid_side.error_i_acumm_preregZ0Z_8 ));
    LocalMux I__11510 (
            .O(N__59459),
            .I(\pid_side.error_i_acumm_preregZ0Z_8 ));
    CascadeMux I__11509 (
            .O(N__59452),
            .I(N__59447));
    InMux I__11508 (
            .O(N__59451),
            .I(N__59444));
    InMux I__11507 (
            .O(N__59450),
            .I(N__59441));
    InMux I__11506 (
            .O(N__59447),
            .I(N__59438));
    LocalMux I__11505 (
            .O(N__59444),
            .I(\pid_side.N_217 ));
    LocalMux I__11504 (
            .O(N__59441),
            .I(\pid_side.N_217 ));
    LocalMux I__11503 (
            .O(N__59438),
            .I(\pid_side.N_217 ));
    InMux I__11502 (
            .O(N__59431),
            .I(N__59427));
    InMux I__11501 (
            .O(N__59430),
            .I(N__59423));
    LocalMux I__11500 (
            .O(N__59427),
            .I(N__59420));
    InMux I__11499 (
            .O(N__59426),
            .I(N__59417));
    LocalMux I__11498 (
            .O(N__59423),
            .I(\pid_side.error_i_acumm_preregZ0Z_7 ));
    Odrv4 I__11497 (
            .O(N__59420),
            .I(\pid_side.error_i_acumm_preregZ0Z_7 ));
    LocalMux I__11496 (
            .O(N__59417),
            .I(\pid_side.error_i_acumm_preregZ0Z_7 ));
    SRMux I__11495 (
            .O(N__59410),
            .I(N__59406));
    SRMux I__11494 (
            .O(N__59409),
            .I(N__59403));
    LocalMux I__11493 (
            .O(N__59406),
            .I(N__59400));
    LocalMux I__11492 (
            .O(N__59403),
            .I(N__59396));
    Span4Mux_v I__11491 (
            .O(N__59400),
            .I(N__59392));
    SRMux I__11490 (
            .O(N__59399),
            .I(N__59389));
    Span4Mux_v I__11489 (
            .O(N__59396),
            .I(N__59386));
    SRMux I__11488 (
            .O(N__59395),
            .I(N__59383));
    Span4Mux_s3_v I__11487 (
            .O(N__59392),
            .I(N__59378));
    LocalMux I__11486 (
            .O(N__59389),
            .I(N__59378));
    Span4Mux_h I__11485 (
            .O(N__59386),
            .I(N__59373));
    LocalMux I__11484 (
            .O(N__59383),
            .I(N__59373));
    Sp12to4 I__11483 (
            .O(N__59378),
            .I(N__59370));
    Span4Mux_h I__11482 (
            .O(N__59373),
            .I(N__59367));
    Odrv12 I__11481 (
            .O(N__59370),
            .I(\pid_side.un1_reset_0_i_3 ));
    Odrv4 I__11480 (
            .O(N__59367),
            .I(\pid_side.un1_reset_0_i_3 ));
    InMux I__11479 (
            .O(N__59362),
            .I(N__59356));
    InMux I__11478 (
            .O(N__59361),
            .I(N__59356));
    LocalMux I__11477 (
            .O(N__59356),
            .I(\pid_side.N_251 ));
    InMux I__11476 (
            .O(N__59353),
            .I(N__59350));
    LocalMux I__11475 (
            .O(N__59350),
            .I(\pid_side.un1_reset_i_a2_5 ));
    InMux I__11474 (
            .O(N__59347),
            .I(N__59344));
    LocalMux I__11473 (
            .O(N__59344),
            .I(\pid_side.N_291 ));
    InMux I__11472 (
            .O(N__59341),
            .I(N__59338));
    LocalMux I__11471 (
            .O(N__59338),
            .I(\pid_side.un1_reset_i_o3_0 ));
    CascadeMux I__11470 (
            .O(N__59335),
            .I(\pid_side.N_631_cascade_ ));
    InMux I__11469 (
            .O(N__59332),
            .I(N__59328));
    InMux I__11468 (
            .O(N__59331),
            .I(N__59325));
    LocalMux I__11467 (
            .O(N__59328),
            .I(N__59320));
    LocalMux I__11466 (
            .O(N__59325),
            .I(N__59320));
    Span4Mux_v I__11465 (
            .O(N__59320),
            .I(N__59317));
    Span4Mux_h I__11464 (
            .O(N__59317),
            .I(N__59314));
    Odrv4 I__11463 (
            .O(N__59314),
            .I(side_order_4));
    CascadeMux I__11462 (
            .O(N__59311),
            .I(\pid_side.un1_reset_i_a2_3_4_cascade_ ));
    CascadeMux I__11461 (
            .O(N__59308),
            .I(N__59304));
    InMux I__11460 (
            .O(N__59307),
            .I(N__59301));
    InMux I__11459 (
            .O(N__59304),
            .I(N__59298));
    LocalMux I__11458 (
            .O(N__59301),
            .I(\pid_side.N_593 ));
    LocalMux I__11457 (
            .O(N__59298),
            .I(\pid_side.N_593 ));
    CascadeMux I__11456 (
            .O(N__59293),
            .I(\pid_side.N_593_cascade_ ));
    InMux I__11455 (
            .O(N__59290),
            .I(N__59287));
    LocalMux I__11454 (
            .O(N__59287),
            .I(N__59284));
    Span4Mux_v I__11453 (
            .O(N__59284),
            .I(N__59280));
    InMux I__11452 (
            .O(N__59283),
            .I(N__59277));
    Sp12to4 I__11451 (
            .O(N__59280),
            .I(N__59272));
    LocalMux I__11450 (
            .O(N__59277),
            .I(N__59272));
    Span12Mux_h I__11449 (
            .O(N__59272),
            .I(N__59269));
    Odrv12 I__11448 (
            .O(N__59269),
            .I(side_order_5));
    InMux I__11447 (
            .O(N__59266),
            .I(N__59263));
    LocalMux I__11446 (
            .O(N__59263),
            .I(N__59260));
    Odrv4 I__11445 (
            .O(N__59260),
            .I(\pid_side.N_11_i ));
    CascadeMux I__11444 (
            .O(N__59257),
            .I(N__59246));
    CascadeMux I__11443 (
            .O(N__59256),
            .I(N__59243));
    CascadeMux I__11442 (
            .O(N__59255),
            .I(N__59238));
    InMux I__11441 (
            .O(N__59254),
            .I(N__59230));
    InMux I__11440 (
            .O(N__59253),
            .I(N__59230));
    InMux I__11439 (
            .O(N__59252),
            .I(N__59230));
    InMux I__11438 (
            .O(N__59251),
            .I(N__59217));
    InMux I__11437 (
            .O(N__59250),
            .I(N__59217));
    InMux I__11436 (
            .O(N__59249),
            .I(N__59217));
    InMux I__11435 (
            .O(N__59246),
            .I(N__59217));
    InMux I__11434 (
            .O(N__59243),
            .I(N__59217));
    InMux I__11433 (
            .O(N__59242),
            .I(N__59217));
    InMux I__11432 (
            .O(N__59241),
            .I(N__59210));
    InMux I__11431 (
            .O(N__59238),
            .I(N__59210));
    InMux I__11430 (
            .O(N__59237),
            .I(N__59210));
    LocalMux I__11429 (
            .O(N__59230),
            .I(N__59207));
    LocalMux I__11428 (
            .O(N__59217),
            .I(\pid_side.N_386 ));
    LocalMux I__11427 (
            .O(N__59210),
            .I(\pid_side.N_386 ));
    Odrv4 I__11426 (
            .O(N__59207),
            .I(\pid_side.N_386 ));
    CascadeMux I__11425 (
            .O(N__59200),
            .I(N__59195));
    InMux I__11424 (
            .O(N__59199),
            .I(N__59190));
    InMux I__11423 (
            .O(N__59198),
            .I(N__59181));
    InMux I__11422 (
            .O(N__59195),
            .I(N__59181));
    InMux I__11421 (
            .O(N__59194),
            .I(N__59181));
    InMux I__11420 (
            .O(N__59193),
            .I(N__59181));
    LocalMux I__11419 (
            .O(N__59190),
            .I(\pid_side.N_631 ));
    LocalMux I__11418 (
            .O(N__59181),
            .I(\pid_side.N_631 ));
    InMux I__11417 (
            .O(N__59176),
            .I(N__59172));
    InMux I__11416 (
            .O(N__59175),
            .I(N__59169));
    LocalMux I__11415 (
            .O(N__59172),
            .I(N__59166));
    LocalMux I__11414 (
            .O(N__59169),
            .I(N__59163));
    Span4Mux_v I__11413 (
            .O(N__59166),
            .I(N__59160));
    Span4Mux_h I__11412 (
            .O(N__59163),
            .I(N__59157));
    Span4Mux_h I__11411 (
            .O(N__59160),
            .I(N__59154));
    Odrv4 I__11410 (
            .O(N__59157),
            .I(side_order_0));
    Odrv4 I__11409 (
            .O(N__59154),
            .I(side_order_0));
    CEMux I__11408 (
            .O(N__59149),
            .I(N__59145));
    CEMux I__11407 (
            .O(N__59148),
            .I(N__59142));
    LocalMux I__11406 (
            .O(N__59145),
            .I(N__59138));
    LocalMux I__11405 (
            .O(N__59142),
            .I(N__59135));
    CEMux I__11404 (
            .O(N__59141),
            .I(N__59132));
    Span4Mux_v I__11403 (
            .O(N__59138),
            .I(N__59129));
    Span4Mux_v I__11402 (
            .O(N__59135),
            .I(N__59126));
    LocalMux I__11401 (
            .O(N__59132),
            .I(N__59123));
    Span4Mux_s1_v I__11400 (
            .O(N__59129),
            .I(N__59120));
    Span4Mux_h I__11399 (
            .O(N__59126),
            .I(N__59115));
    Span4Mux_h I__11398 (
            .O(N__59123),
            .I(N__59115));
    Odrv4 I__11397 (
            .O(N__59120),
            .I(\pid_side.state_0_1 ));
    Odrv4 I__11396 (
            .O(N__59115),
            .I(\pid_side.state_0_1 ));
    InMux I__11395 (
            .O(N__59110),
            .I(N__59107));
    LocalMux I__11394 (
            .O(N__59107),
            .I(\pid_side.un11lto30_i_a2_0_and ));
    InMux I__11393 (
            .O(N__59104),
            .I(N__59101));
    LocalMux I__11392 (
            .O(N__59101),
            .I(N__59098));
    Odrv4 I__11391 (
            .O(N__59098),
            .I(\pid_side.un11lto30_i_a2_2_and ));
    InMux I__11390 (
            .O(N__59095),
            .I(N__59092));
    LocalMux I__11389 (
            .O(N__59092),
            .I(\pid_side.source_pid_9_i_0_o3_0_11 ));
    InMux I__11388 (
            .O(N__59089),
            .I(bfn_14_4_0_));
    InMux I__11387 (
            .O(N__59086),
            .I(N__59083));
    LocalMux I__11386 (
            .O(N__59083),
            .I(N__59080));
    Span4Mux_v I__11385 (
            .O(N__59080),
            .I(N__59074));
    InMux I__11384 (
            .O(N__59079),
            .I(N__59071));
    InMux I__11383 (
            .O(N__59078),
            .I(N__59066));
    InMux I__11382 (
            .O(N__59077),
            .I(N__59066));
    Odrv4 I__11381 (
            .O(N__59074),
            .I(\pid_front.error_d_reg_prevZ0Z_6 ));
    LocalMux I__11380 (
            .O(N__59071),
            .I(\pid_front.error_d_reg_prevZ0Z_6 ));
    LocalMux I__11379 (
            .O(N__59066),
            .I(\pid_front.error_d_reg_prevZ0Z_6 ));
    InMux I__11378 (
            .O(N__59059),
            .I(N__59056));
    LocalMux I__11377 (
            .O(N__59056),
            .I(N__59053));
    Span4Mux_h I__11376 (
            .O(N__59053),
            .I(N__59050));
    Sp12to4 I__11375 (
            .O(N__59050),
            .I(N__59047));
    Span12Mux_v I__11374 (
            .O(N__59047),
            .I(N__59044));
    Odrv12 I__11373 (
            .O(N__59044),
            .I(\pid_front.O_0_5 ));
    CascadeMux I__11372 (
            .O(N__59041),
            .I(N__59036));
    CascadeMux I__11371 (
            .O(N__59040),
            .I(N__59033));
    InMux I__11370 (
            .O(N__59039),
            .I(N__59030));
    InMux I__11369 (
            .O(N__59036),
            .I(N__59025));
    InMux I__11368 (
            .O(N__59033),
            .I(N__59025));
    LocalMux I__11367 (
            .O(N__59030),
            .I(\pid_front.error_p_regZ0Z_1 ));
    LocalMux I__11366 (
            .O(N__59025),
            .I(\pid_front.error_p_regZ0Z_1 ));
    CascadeMux I__11365 (
            .O(N__59020),
            .I(\pid_front.un1_pid_prereg_9_0_cascade_ ));
    CascadeMux I__11364 (
            .O(N__59017),
            .I(N__59014));
    InMux I__11363 (
            .O(N__59014),
            .I(N__59011));
    LocalMux I__11362 (
            .O(N__59011),
            .I(N__59008));
    Odrv12 I__11361 (
            .O(N__59008),
            .I(\pid_front.error_d_reg_prev_esr_RNIMRLTZ0Z_0 ));
    InMux I__11360 (
            .O(N__59005),
            .I(N__59002));
    LocalMux I__11359 (
            .O(N__59002),
            .I(N__58999));
    Span12Mux_s3_v I__11358 (
            .O(N__58999),
            .I(N__58996));
    Span12Mux_h I__11357 (
            .O(N__58996),
            .I(N__58993));
    Odrv12 I__11356 (
            .O(N__58993),
            .I(\pid_front.O_4 ));
    InMux I__11355 (
            .O(N__58990),
            .I(N__58982));
    InMux I__11354 (
            .O(N__58989),
            .I(N__58982));
    InMux I__11353 (
            .O(N__58988),
            .I(N__58977));
    InMux I__11352 (
            .O(N__58987),
            .I(N__58977));
    LocalMux I__11351 (
            .O(N__58982),
            .I(\pid_front.error_d_reg_prevZ0Z_0 ));
    LocalMux I__11350 (
            .O(N__58977),
            .I(\pid_front.error_d_reg_prevZ0Z_0 ));
    InMux I__11349 (
            .O(N__58972),
            .I(N__58969));
    LocalMux I__11348 (
            .O(N__58969),
            .I(N__58966));
    Span4Mux_v I__11347 (
            .O(N__58966),
            .I(N__58963));
    Odrv4 I__11346 (
            .O(N__58963),
            .I(\pid_front.error_d_reg_prev_esr_RNIAHDKZ0Z_0 ));
    InMux I__11345 (
            .O(N__58960),
            .I(N__58957));
    LocalMux I__11344 (
            .O(N__58957),
            .I(N__58954));
    Odrv12 I__11343 (
            .O(N__58954),
            .I(\pid_front.N_5_0 ));
    CascadeMux I__11342 (
            .O(N__58951),
            .I(\pid_front.error_p_reg_esr_RNI6D5L7Z0Z_12_cascade_ ));
    InMux I__11341 (
            .O(N__58948),
            .I(N__58945));
    LocalMux I__11340 (
            .O(N__58945),
            .I(N__58941));
    InMux I__11339 (
            .O(N__58944),
            .I(N__58938));
    Sp12to4 I__11338 (
            .O(N__58941),
            .I(N__58933));
    LocalMux I__11337 (
            .O(N__58938),
            .I(N__58933));
    Odrv12 I__11336 (
            .O(N__58933),
            .I(\pid_front.un1_pid_prereg_0_axb_14 ));
    InMux I__11335 (
            .O(N__58930),
            .I(N__58927));
    LocalMux I__11334 (
            .O(N__58927),
            .I(N__58924));
    Span12Mux_s4_v I__11333 (
            .O(N__58924),
            .I(N__58921));
    Span12Mux_h I__11332 (
            .O(N__58921),
            .I(N__58918));
    Odrv12 I__11331 (
            .O(N__58918),
            .I(\pid_front.O_3 ));
    InMux I__11330 (
            .O(N__58915),
            .I(N__58906));
    InMux I__11329 (
            .O(N__58914),
            .I(N__58906));
    InMux I__11328 (
            .O(N__58913),
            .I(N__58899));
    InMux I__11327 (
            .O(N__58912),
            .I(N__58899));
    InMux I__11326 (
            .O(N__58911),
            .I(N__58899));
    LocalMux I__11325 (
            .O(N__58906),
            .I(\pid_front.error_d_regZ0Z_0 ));
    LocalMux I__11324 (
            .O(N__58899),
            .I(\pid_front.error_d_regZ0Z_0 ));
    InMux I__11323 (
            .O(N__58894),
            .I(N__58891));
    LocalMux I__11322 (
            .O(N__58891),
            .I(\pid_front.pid_preregZ0Z_28 ));
    InMux I__11321 (
            .O(N__58888),
            .I(\pid_front.un1_pid_prereg_0_cry_27 ));
    InMux I__11320 (
            .O(N__58885),
            .I(N__58882));
    LocalMux I__11319 (
            .O(N__58882),
            .I(\pid_front.pid_preregZ0Z_29 ));
    InMux I__11318 (
            .O(N__58879),
            .I(\pid_front.un1_pid_prereg_0_cry_28 ));
    InMux I__11317 (
            .O(N__58876),
            .I(\pid_front.un1_pid_prereg_0_cry_29 ));
    CascadeMux I__11316 (
            .O(N__58873),
            .I(N__58868));
    InMux I__11315 (
            .O(N__58872),
            .I(N__58863));
    InMux I__11314 (
            .O(N__58871),
            .I(N__58855));
    InMux I__11313 (
            .O(N__58868),
            .I(N__58855));
    InMux I__11312 (
            .O(N__58867),
            .I(N__58855));
    InMux I__11311 (
            .O(N__58866),
            .I(N__58852));
    LocalMux I__11310 (
            .O(N__58863),
            .I(N__58849));
    InMux I__11309 (
            .O(N__58862),
            .I(N__58846));
    LocalMux I__11308 (
            .O(N__58855),
            .I(N__58843));
    LocalMux I__11307 (
            .O(N__58852),
            .I(N__58840));
    Span4Mux_h I__11306 (
            .O(N__58849),
            .I(N__58836));
    LocalMux I__11305 (
            .O(N__58846),
            .I(N__58829));
    Span4Mux_v I__11304 (
            .O(N__58843),
            .I(N__58829));
    Span4Mux_h I__11303 (
            .O(N__58840),
            .I(N__58829));
    InMux I__11302 (
            .O(N__58839),
            .I(N__58826));
    Odrv4 I__11301 (
            .O(N__58836),
            .I(\pid_front.pid_preregZ0Z_30 ));
    Odrv4 I__11300 (
            .O(N__58829),
            .I(\pid_front.pid_preregZ0Z_30 ));
    LocalMux I__11299 (
            .O(N__58826),
            .I(\pid_front.pid_preregZ0Z_30 ));
    CascadeMux I__11298 (
            .O(N__58819),
            .I(\pid_front.N_2358_i_cascade_ ));
    InMux I__11297 (
            .O(N__58816),
            .I(N__58813));
    LocalMux I__11296 (
            .O(N__58813),
            .I(\pid_front.error_p_reg_esr_RNI6B6FZ0Z_6 ));
    InMux I__11295 (
            .O(N__58810),
            .I(N__58807));
    LocalMux I__11294 (
            .O(N__58807),
            .I(\pid_front.error_p_reg_esr_RNIBG6F_0Z0Z_7 ));
    CascadeMux I__11293 (
            .O(N__58804),
            .I(\pid_front.error_p_reg_esr_RNI6B6FZ0Z_6_cascade_ ));
    InMux I__11292 (
            .O(N__58801),
            .I(N__58798));
    LocalMux I__11291 (
            .O(N__58798),
            .I(N__58795));
    Odrv4 I__11290 (
            .O(N__58795),
            .I(\pid_front.error_p_reg_esr_RNI3K9L1_0Z0Z_6 ));
    CascadeMux I__11289 (
            .O(N__58792),
            .I(\pid_front.error_p_reg_esr_RNIMVC9Z0Z_6_cascade_ ));
    InMux I__11288 (
            .O(N__58789),
            .I(N__58786));
    LocalMux I__11287 (
            .O(N__58786),
            .I(\pid_front.error_p_reg_esr_RNI80EDDZ0Z_17 ));
    InMux I__11286 (
            .O(N__58783),
            .I(N__58780));
    LocalMux I__11285 (
            .O(N__58780),
            .I(N__58777));
    Span4Mux_h I__11284 (
            .O(N__58777),
            .I(N__58774));
    Odrv4 I__11283 (
            .O(N__58774),
            .I(\pid_front.pid_preregZ0Z_20 ));
    InMux I__11282 (
            .O(N__58771),
            .I(\pid_front.un1_pid_prereg_0_cry_19 ));
    InMux I__11281 (
            .O(N__58768),
            .I(N__58765));
    LocalMux I__11280 (
            .O(N__58765),
            .I(\pid_front.error_p_reg_esr_RNIRNJEDZ0Z_18 ));
    CascadeMux I__11279 (
            .O(N__58762),
            .I(N__58759));
    InMux I__11278 (
            .O(N__58759),
            .I(N__58756));
    LocalMux I__11277 (
            .O(N__58756),
            .I(N__58753));
    Odrv4 I__11276 (
            .O(N__58753),
            .I(\pid_front.error_p_reg_esr_RNIQOPM6Z0Z_18 ));
    InMux I__11275 (
            .O(N__58750),
            .I(N__58747));
    LocalMux I__11274 (
            .O(N__58747),
            .I(N__58744));
    Span4Mux_h I__11273 (
            .O(N__58744),
            .I(N__58741));
    Odrv4 I__11272 (
            .O(N__58741),
            .I(\pid_front.pid_preregZ0Z_21 ));
    InMux I__11271 (
            .O(N__58738),
            .I(\pid_front.un1_pid_prereg_0_cry_20 ));
    CascadeMux I__11270 (
            .O(N__58735),
            .I(N__58732));
    InMux I__11269 (
            .O(N__58732),
            .I(N__58729));
    LocalMux I__11268 (
            .O(N__58729),
            .I(\pid_front.error_p_reg_esr_RNI1VPN6Z0Z_19 ));
    InMux I__11267 (
            .O(N__58726),
            .I(N__58723));
    LocalMux I__11266 (
            .O(N__58723),
            .I(N__58720));
    Span4Mux_h I__11265 (
            .O(N__58720),
            .I(N__58717));
    Odrv4 I__11264 (
            .O(N__58717),
            .I(\pid_front.pid_preregZ0Z_22 ));
    InMux I__11263 (
            .O(N__58714),
            .I(\pid_front.un1_pid_prereg_0_cry_21 ));
    CascadeMux I__11262 (
            .O(N__58711),
            .I(N__58708));
    InMux I__11261 (
            .O(N__58708),
            .I(N__58705));
    LocalMux I__11260 (
            .O(N__58705),
            .I(N__58702));
    Span4Mux_h I__11259 (
            .O(N__58702),
            .I(N__58699));
    Odrv4 I__11258 (
            .O(N__58699),
            .I(\pid_front.pid_preregZ0Z_23 ));
    InMux I__11257 (
            .O(N__58696),
            .I(bfn_13_26_0_));
    InMux I__11256 (
            .O(N__58693),
            .I(N__58690));
    LocalMux I__11255 (
            .O(N__58690),
            .I(\pid_front.pid_preregZ0Z_24 ));
    InMux I__11254 (
            .O(N__58687),
            .I(\pid_front.un1_pid_prereg_0_cry_23 ));
    InMux I__11253 (
            .O(N__58684),
            .I(N__58681));
    LocalMux I__11252 (
            .O(N__58681),
            .I(\pid_front.pid_preregZ0Z_25 ));
    InMux I__11251 (
            .O(N__58678),
            .I(\pid_front.un1_pid_prereg_0_cry_24 ));
    InMux I__11250 (
            .O(N__58675),
            .I(N__58672));
    LocalMux I__11249 (
            .O(N__58672),
            .I(\pid_front.pid_preregZ0Z_26 ));
    InMux I__11248 (
            .O(N__58669),
            .I(\pid_front.un1_pid_prereg_0_cry_25 ));
    CascadeMux I__11247 (
            .O(N__58666),
            .I(N__58663));
    InMux I__11246 (
            .O(N__58663),
            .I(N__58660));
    LocalMux I__11245 (
            .O(N__58660),
            .I(\pid_front.pid_preregZ0Z_27 ));
    InMux I__11244 (
            .O(N__58657),
            .I(\pid_front.un1_pid_prereg_0_cry_26 ));
    InMux I__11243 (
            .O(N__58654),
            .I(N__58650));
    CascadeMux I__11242 (
            .O(N__58653),
            .I(N__58646));
    LocalMux I__11241 (
            .O(N__58650),
            .I(N__58643));
    InMux I__11240 (
            .O(N__58649),
            .I(N__58638));
    InMux I__11239 (
            .O(N__58646),
            .I(N__58638));
    Sp12to4 I__11238 (
            .O(N__58643),
            .I(N__58635));
    LocalMux I__11237 (
            .O(N__58638),
            .I(N__58632));
    Span12Mux_v I__11236 (
            .O(N__58635),
            .I(N__58629));
    Span4Mux_h I__11235 (
            .O(N__58632),
            .I(N__58626));
    Odrv12 I__11234 (
            .O(N__58629),
            .I(\pid_front.pid_preregZ0Z_11 ));
    Odrv4 I__11233 (
            .O(N__58626),
            .I(\pid_front.pid_preregZ0Z_11 ));
    InMux I__11232 (
            .O(N__58621),
            .I(\pid_front.un1_pid_prereg_0_cry_10 ));
    CascadeMux I__11231 (
            .O(N__58618),
            .I(N__58614));
    InMux I__11230 (
            .O(N__58617),
            .I(N__58611));
    InMux I__11229 (
            .O(N__58614),
            .I(N__58608));
    LocalMux I__11228 (
            .O(N__58611),
            .I(N__58601));
    LocalMux I__11227 (
            .O(N__58608),
            .I(N__58601));
    InMux I__11226 (
            .O(N__58607),
            .I(N__58596));
    InMux I__11225 (
            .O(N__58606),
            .I(N__58596));
    Odrv4 I__11224 (
            .O(N__58601),
            .I(\pid_front.pid_preregZ0Z_12 ));
    LocalMux I__11223 (
            .O(N__58596),
            .I(\pid_front.pid_preregZ0Z_12 ));
    InMux I__11222 (
            .O(N__58591),
            .I(\pid_front.un1_pid_prereg_0_cry_11 ));
    CascadeMux I__11221 (
            .O(N__58588),
            .I(N__58585));
    InMux I__11220 (
            .O(N__58585),
            .I(N__58579));
    InMux I__11219 (
            .O(N__58584),
            .I(N__58579));
    LocalMux I__11218 (
            .O(N__58579),
            .I(N__58575));
    InMux I__11217 (
            .O(N__58578),
            .I(N__58572));
    Span4Mux_h I__11216 (
            .O(N__58575),
            .I(N__58567));
    LocalMux I__11215 (
            .O(N__58572),
            .I(N__58564));
    InMux I__11214 (
            .O(N__58571),
            .I(N__58559));
    InMux I__11213 (
            .O(N__58570),
            .I(N__58559));
    Odrv4 I__11212 (
            .O(N__58567),
            .I(\pid_front.pid_preregZ0Z_13 ));
    Odrv4 I__11211 (
            .O(N__58564),
            .I(\pid_front.pid_preregZ0Z_13 ));
    LocalMux I__11210 (
            .O(N__58559),
            .I(\pid_front.pid_preregZ0Z_13 ));
    InMux I__11209 (
            .O(N__58552),
            .I(\pid_front.un1_pid_prereg_0_cry_12 ));
    InMux I__11208 (
            .O(N__58549),
            .I(N__58546));
    LocalMux I__11207 (
            .O(N__58546),
            .I(\pid_front.un1_pid_prereg_0_cry_13_THRU_CO ));
    InMux I__11206 (
            .O(N__58543),
            .I(\pid_front.un1_pid_prereg_0_cry_13 ));
    InMux I__11205 (
            .O(N__58540),
            .I(N__58535));
    CascadeMux I__11204 (
            .O(N__58539),
            .I(N__58532));
    CascadeMux I__11203 (
            .O(N__58538),
            .I(N__58529));
    LocalMux I__11202 (
            .O(N__58535),
            .I(N__58526));
    InMux I__11201 (
            .O(N__58532),
            .I(N__58521));
    InMux I__11200 (
            .O(N__58529),
            .I(N__58521));
    Odrv4 I__11199 (
            .O(N__58526),
            .I(\pid_front.pid_preregZ0Z_15 ));
    LocalMux I__11198 (
            .O(N__58521),
            .I(\pid_front.pid_preregZ0Z_15 ));
    InMux I__11197 (
            .O(N__58516),
            .I(bfn_13_25_0_));
    InMux I__11196 (
            .O(N__58513),
            .I(N__58510));
    LocalMux I__11195 (
            .O(N__58510),
            .I(\pid_front.pid_preregZ0Z_16 ));
    InMux I__11194 (
            .O(N__58507),
            .I(\pid_front.un1_pid_prereg_0_cry_15 ));
    InMux I__11193 (
            .O(N__58504),
            .I(N__58501));
    LocalMux I__11192 (
            .O(N__58501),
            .I(\pid_front.pid_preregZ0Z_17 ));
    InMux I__11191 (
            .O(N__58498),
            .I(\pid_front.un1_pid_prereg_0_cry_16 ));
    InMux I__11190 (
            .O(N__58495),
            .I(N__58492));
    LocalMux I__11189 (
            .O(N__58492),
            .I(\pid_front.pid_preregZ0Z_18 ));
    InMux I__11188 (
            .O(N__58489),
            .I(\pid_front.un1_pid_prereg_0_cry_17 ));
    CascadeMux I__11187 (
            .O(N__58486),
            .I(N__58483));
    InMux I__11186 (
            .O(N__58483),
            .I(N__58480));
    LocalMux I__11185 (
            .O(N__58480),
            .I(\pid_front.pid_preregZ0Z_19 ));
    InMux I__11184 (
            .O(N__58477),
            .I(\pid_front.un1_pid_prereg_0_cry_18 ));
    InMux I__11183 (
            .O(N__58474),
            .I(\pid_front.un1_pid_prereg_0_cry_2 ));
    InMux I__11182 (
            .O(N__58471),
            .I(N__58468));
    LocalMux I__11181 (
            .O(N__58468),
            .I(N__58465));
    Sp12to4 I__11180 (
            .O(N__58465),
            .I(N__58460));
    InMux I__11179 (
            .O(N__58464),
            .I(N__58454));
    InMux I__11178 (
            .O(N__58463),
            .I(N__58454));
    Span12Mux_v I__11177 (
            .O(N__58460),
            .I(N__58451));
    InMux I__11176 (
            .O(N__58459),
            .I(N__58448));
    LocalMux I__11175 (
            .O(N__58454),
            .I(N__58445));
    Odrv12 I__11174 (
            .O(N__58451),
            .I(\pid_front.pid_preregZ0Z_4 ));
    LocalMux I__11173 (
            .O(N__58448),
            .I(\pid_front.pid_preregZ0Z_4 ));
    Odrv4 I__11172 (
            .O(N__58445),
            .I(\pid_front.pid_preregZ0Z_4 ));
    InMux I__11171 (
            .O(N__58438),
            .I(\pid_front.un1_pid_prereg_0_cry_3 ));
    InMux I__11170 (
            .O(N__58435),
            .I(N__58432));
    LocalMux I__11169 (
            .O(N__58432),
            .I(N__58426));
    InMux I__11168 (
            .O(N__58431),
            .I(N__58421));
    InMux I__11167 (
            .O(N__58430),
            .I(N__58421));
    InMux I__11166 (
            .O(N__58429),
            .I(N__58418));
    Span4Mux_v I__11165 (
            .O(N__58426),
            .I(N__58413));
    LocalMux I__11164 (
            .O(N__58421),
            .I(N__58413));
    LocalMux I__11163 (
            .O(N__58418),
            .I(\pid_front.pid_preregZ0Z_5 ));
    Odrv4 I__11162 (
            .O(N__58413),
            .I(\pid_front.pid_preregZ0Z_5 ));
    InMux I__11161 (
            .O(N__58408),
            .I(\pid_front.un1_pid_prereg_0_cry_4 ));
    InMux I__11160 (
            .O(N__58405),
            .I(N__58402));
    LocalMux I__11159 (
            .O(N__58402),
            .I(N__58398));
    InMux I__11158 (
            .O(N__58401),
            .I(N__58395));
    Sp12to4 I__11157 (
            .O(N__58398),
            .I(N__58391));
    LocalMux I__11156 (
            .O(N__58395),
            .I(N__58388));
    InMux I__11155 (
            .O(N__58394),
            .I(N__58385));
    Span12Mux_v I__11154 (
            .O(N__58391),
            .I(N__58382));
    Span4Mux_v I__11153 (
            .O(N__58388),
            .I(N__58377));
    LocalMux I__11152 (
            .O(N__58385),
            .I(N__58377));
    Odrv12 I__11151 (
            .O(N__58382),
            .I(\pid_front.pid_preregZ0Z_6 ));
    Odrv4 I__11150 (
            .O(N__58377),
            .I(\pid_front.pid_preregZ0Z_6 ));
    InMux I__11149 (
            .O(N__58372),
            .I(\pid_front.un1_pid_prereg_0_cry_5 ));
    InMux I__11148 (
            .O(N__58369),
            .I(N__58365));
    CascadeMux I__11147 (
            .O(N__58368),
            .I(N__58361));
    LocalMux I__11146 (
            .O(N__58365),
            .I(N__58358));
    CascadeMux I__11145 (
            .O(N__58364),
            .I(N__58355));
    InMux I__11144 (
            .O(N__58361),
            .I(N__58352));
    Span4Mux_h I__11143 (
            .O(N__58358),
            .I(N__58349));
    InMux I__11142 (
            .O(N__58355),
            .I(N__58346));
    LocalMux I__11141 (
            .O(N__58352),
            .I(N__58343));
    Sp12to4 I__11140 (
            .O(N__58349),
            .I(N__58340));
    LocalMux I__11139 (
            .O(N__58346),
            .I(N__58335));
    Span4Mux_v I__11138 (
            .O(N__58343),
            .I(N__58335));
    Odrv12 I__11137 (
            .O(N__58340),
            .I(\pid_front.pid_preregZ0Z_7 ));
    Odrv4 I__11136 (
            .O(N__58335),
            .I(\pid_front.pid_preregZ0Z_7 ));
    InMux I__11135 (
            .O(N__58330),
            .I(bfn_13_24_0_));
    InMux I__11134 (
            .O(N__58327),
            .I(N__58323));
    InMux I__11133 (
            .O(N__58326),
            .I(N__58320));
    LocalMux I__11132 (
            .O(N__58323),
            .I(N__58317));
    LocalMux I__11131 (
            .O(N__58320),
            .I(N__58314));
    Span4Mux_h I__11130 (
            .O(N__58317),
            .I(N__58311));
    Odrv4 I__11129 (
            .O(N__58314),
            .I(\pid_front.error_p_reg_esr_RNI3K9L1Z0Z_6 ));
    Odrv4 I__11128 (
            .O(N__58311),
            .I(\pid_front.error_p_reg_esr_RNI3K9L1Z0Z_6 ));
    CascadeMux I__11127 (
            .O(N__58306),
            .I(N__58303));
    InMux I__11126 (
            .O(N__58303),
            .I(N__58300));
    LocalMux I__11125 (
            .O(N__58300),
            .I(\pid_front.error_p_reg_esr_RNIS0F23Z0Z_7 ));
    CascadeMux I__11124 (
            .O(N__58297),
            .I(N__58294));
    InMux I__11123 (
            .O(N__58294),
            .I(N__58291));
    LocalMux I__11122 (
            .O(N__58291),
            .I(N__58288));
    Sp12to4 I__11121 (
            .O(N__58288),
            .I(N__58285));
    Span12Mux_s8_v I__11120 (
            .O(N__58285),
            .I(N__58280));
    InMux I__11119 (
            .O(N__58284),
            .I(N__58275));
    InMux I__11118 (
            .O(N__58283),
            .I(N__58275));
    Span12Mux_v I__11117 (
            .O(N__58280),
            .I(N__58272));
    LocalMux I__11116 (
            .O(N__58275),
            .I(N__58269));
    Odrv12 I__11115 (
            .O(N__58272),
            .I(\pid_front.pid_preregZ0Z_8 ));
    Odrv12 I__11114 (
            .O(N__58269),
            .I(\pid_front.pid_preregZ0Z_8 ));
    InMux I__11113 (
            .O(N__58264),
            .I(\pid_front.un1_pid_prereg_0_cry_7 ));
    InMux I__11112 (
            .O(N__58261),
            .I(N__58258));
    LocalMux I__11111 (
            .O(N__58258),
            .I(\pid_front.error_p_reg_esr_RNIV7CQ2Z0Z_8 ));
    CascadeMux I__11110 (
            .O(N__58255),
            .I(N__58251));
    InMux I__11109 (
            .O(N__58254),
            .I(N__58248));
    InMux I__11108 (
            .O(N__58251),
            .I(N__58245));
    LocalMux I__11107 (
            .O(N__58248),
            .I(\pid_front.error_p_reg_esr_RNIPC5D1Z0Z_7 ));
    LocalMux I__11106 (
            .O(N__58245),
            .I(\pid_front.error_p_reg_esr_RNIPC5D1Z0Z_7 ));
    InMux I__11105 (
            .O(N__58240),
            .I(N__58237));
    LocalMux I__11104 (
            .O(N__58237),
            .I(N__58234));
    Span4Mux_v I__11103 (
            .O(N__58234),
            .I(N__58231));
    Span4Mux_v I__11102 (
            .O(N__58231),
            .I(N__58226));
    InMux I__11101 (
            .O(N__58230),
            .I(N__58221));
    InMux I__11100 (
            .O(N__58229),
            .I(N__58221));
    Span4Mux_v I__11099 (
            .O(N__58226),
            .I(N__58218));
    LocalMux I__11098 (
            .O(N__58221),
            .I(N__58215));
    Odrv4 I__11097 (
            .O(N__58218),
            .I(\pid_front.pid_preregZ0Z_9 ));
    Odrv4 I__11096 (
            .O(N__58215),
            .I(\pid_front.pid_preregZ0Z_9 ));
    InMux I__11095 (
            .O(N__58210),
            .I(\pid_front.un1_pid_prereg_0_cry_8 ));
    InMux I__11094 (
            .O(N__58207),
            .I(N__58204));
    LocalMux I__11093 (
            .O(N__58204),
            .I(N__58201));
    Sp12to4 I__11092 (
            .O(N__58201),
            .I(N__58196));
    InMux I__11091 (
            .O(N__58200),
            .I(N__58191));
    InMux I__11090 (
            .O(N__58199),
            .I(N__58191));
    Span12Mux_v I__11089 (
            .O(N__58196),
            .I(N__58188));
    LocalMux I__11088 (
            .O(N__58191),
            .I(N__58185));
    Odrv12 I__11087 (
            .O(N__58188),
            .I(\pid_front.pid_preregZ0Z_10 ));
    Odrv4 I__11086 (
            .O(N__58185),
            .I(\pid_front.pid_preregZ0Z_10 ));
    InMux I__11085 (
            .O(N__58180),
            .I(\pid_front.un1_pid_prereg_0_cry_9 ));
    InMux I__11084 (
            .O(N__58177),
            .I(N__58174));
    LocalMux I__11083 (
            .O(N__58174),
            .I(\pid_front.state_RNIPKTDZ0Z_0 ));
    CascadeMux I__11082 (
            .O(N__58171),
            .I(\pid_front.state_RNIPKTDZ0Z_0_cascade_ ));
    InMux I__11081 (
            .O(N__58168),
            .I(\pid_front.un1_pid_prereg_0_cry_0_c_THRU_CO ));
    InMux I__11080 (
            .O(N__58165),
            .I(N__58162));
    LocalMux I__11079 (
            .O(N__58162),
            .I(N__58159));
    Span4Mux_h I__11078 (
            .O(N__58159),
            .I(N__58156));
    Sp12to4 I__11077 (
            .O(N__58156),
            .I(N__58151));
    InMux I__11076 (
            .O(N__58155),
            .I(N__58146));
    InMux I__11075 (
            .O(N__58154),
            .I(N__58146));
    Odrv12 I__11074 (
            .O(N__58151),
            .I(\pid_front.pid_preregZ0Z_1 ));
    LocalMux I__11073 (
            .O(N__58146),
            .I(\pid_front.pid_preregZ0Z_1 ));
    InMux I__11072 (
            .O(N__58141),
            .I(\pid_front.un1_pid_prereg_0_cry_0 ));
    InMux I__11071 (
            .O(N__58138),
            .I(N__58135));
    LocalMux I__11070 (
            .O(N__58135),
            .I(N__58132));
    Span4Mux_h I__11069 (
            .O(N__58132),
            .I(N__58129));
    Odrv4 I__11068 (
            .O(N__58129),
            .I(\pid_front.error_d_reg_prev_esr_RNID19M1Z0Z_1 ));
    InMux I__11067 (
            .O(N__58126),
            .I(\pid_front.un1_pid_prereg_0_cry_1 ));
    InMux I__11066 (
            .O(N__58123),
            .I(N__58117));
    InMux I__11065 (
            .O(N__58122),
            .I(N__58117));
    LocalMux I__11064 (
            .O(N__58117),
            .I(drone_H_disp_front_11));
    CascadeMux I__11063 (
            .O(N__58114),
            .I(N__58111));
    InMux I__11062 (
            .O(N__58111),
            .I(N__58105));
    InMux I__11061 (
            .O(N__58110),
            .I(N__58105));
    LocalMux I__11060 (
            .O(N__58105),
            .I(front_command_7));
    CascadeMux I__11059 (
            .O(N__58102),
            .I(N__58099));
    InMux I__11058 (
            .O(N__58099),
            .I(N__58096));
    LocalMux I__11057 (
            .O(N__58096),
            .I(N__58093));
    Odrv4 I__11056 (
            .O(N__58093),
            .I(\pid_front.error_axbZ0Z_7 ));
    CascadeMux I__11055 (
            .O(N__58090),
            .I(N__58087));
    InMux I__11054 (
            .O(N__58087),
            .I(N__58082));
    InMux I__11053 (
            .O(N__58086),
            .I(N__58077));
    InMux I__11052 (
            .O(N__58085),
            .I(N__58077));
    LocalMux I__11051 (
            .O(N__58082),
            .I(drone_H_disp_front_12));
    LocalMux I__11050 (
            .O(N__58077),
            .I(drone_H_disp_front_12));
    InMux I__11049 (
            .O(N__58072),
            .I(N__58069));
    LocalMux I__11048 (
            .O(N__58069),
            .I(N__58066));
    Odrv4 I__11047 (
            .O(N__58066),
            .I(drone_H_disp_front_i_12));
    InMux I__11046 (
            .O(N__58063),
            .I(N__58060));
    LocalMux I__11045 (
            .O(N__58060),
            .I(\pid_front.un1_reset_i_a2_5 ));
    InMux I__11044 (
            .O(N__58057),
            .I(N__58054));
    LocalMux I__11043 (
            .O(N__58054),
            .I(N__58051));
    Odrv4 I__11042 (
            .O(N__58051),
            .I(\pid_front.source_pid10lt4_0 ));
    InMux I__11041 (
            .O(N__58048),
            .I(N__58045));
    LocalMux I__11040 (
            .O(N__58045),
            .I(N__58042));
    Odrv4 I__11039 (
            .O(N__58042),
            .I(\pid_front.un1_reset_i_a2_4 ));
    CascadeMux I__11038 (
            .O(N__58039),
            .I(\pid_front.N_162_cascade_ ));
    InMux I__11037 (
            .O(N__58036),
            .I(N__58030));
    InMux I__11036 (
            .O(N__58035),
            .I(N__58025));
    InMux I__11035 (
            .O(N__58034),
            .I(N__58020));
    InMux I__11034 (
            .O(N__58033),
            .I(N__58020));
    LocalMux I__11033 (
            .O(N__58030),
            .I(N__58017));
    InMux I__11032 (
            .O(N__58029),
            .I(N__58013));
    InMux I__11031 (
            .O(N__58028),
            .I(N__58008));
    LocalMux I__11030 (
            .O(N__58025),
            .I(N__58003));
    LocalMux I__11029 (
            .O(N__58020),
            .I(N__58003));
    Span4Mux_v I__11028 (
            .O(N__58017),
            .I(N__58000));
    InMux I__11027 (
            .O(N__58016),
            .I(N__57997));
    LocalMux I__11026 (
            .O(N__58013),
            .I(N__57994));
    InMux I__11025 (
            .O(N__58012),
            .I(N__57991));
    InMux I__11024 (
            .O(N__58011),
            .I(N__57988));
    LocalMux I__11023 (
            .O(N__58008),
            .I(N__57983));
    Span4Mux_h I__11022 (
            .O(N__58003),
            .I(N__57983));
    Span4Mux_h I__11021 (
            .O(N__58000),
            .I(N__57980));
    LocalMux I__11020 (
            .O(N__57997),
            .I(N__57977));
    Span4Mux_h I__11019 (
            .O(N__57994),
            .I(N__57968));
    LocalMux I__11018 (
            .O(N__57991),
            .I(N__57968));
    LocalMux I__11017 (
            .O(N__57988),
            .I(N__57968));
    Span4Mux_v I__11016 (
            .O(N__57983),
            .I(N__57968));
    Span4Mux_v I__11015 (
            .O(N__57980),
            .I(N__57965));
    Span4Mux_h I__11014 (
            .O(N__57977),
            .I(N__57962));
    Span4Mux_v I__11013 (
            .O(N__57968),
            .I(N__57959));
    Odrv4 I__11012 (
            .O(N__57965),
            .I(uart_drone_data_3));
    Odrv4 I__11011 (
            .O(N__57962),
            .I(uart_drone_data_3));
    Odrv4 I__11010 (
            .O(N__57959),
            .I(uart_drone_data_3));
    InMux I__11009 (
            .O(N__57952),
            .I(N__57949));
    LocalMux I__11008 (
            .O(N__57949),
            .I(N__57943));
    InMux I__11007 (
            .O(N__57948),
            .I(N__57935));
    InMux I__11006 (
            .O(N__57947),
            .I(N__57932));
    InMux I__11005 (
            .O(N__57946),
            .I(N__57929));
    Span4Mux_h I__11004 (
            .O(N__57943),
            .I(N__57926));
    InMux I__11003 (
            .O(N__57942),
            .I(N__57921));
    InMux I__11002 (
            .O(N__57941),
            .I(N__57921));
    InMux I__11001 (
            .O(N__57940),
            .I(N__57918));
    InMux I__11000 (
            .O(N__57939),
            .I(N__57915));
    InMux I__10999 (
            .O(N__57938),
            .I(N__57912));
    LocalMux I__10998 (
            .O(N__57935),
            .I(N__57907));
    LocalMux I__10997 (
            .O(N__57932),
            .I(N__57907));
    LocalMux I__10996 (
            .O(N__57929),
            .I(N__57902));
    Span4Mux_v I__10995 (
            .O(N__57926),
            .I(N__57902));
    LocalMux I__10994 (
            .O(N__57921),
            .I(N__57899));
    LocalMux I__10993 (
            .O(N__57918),
            .I(N__57896));
    LocalMux I__10992 (
            .O(N__57915),
            .I(N__57885));
    LocalMux I__10991 (
            .O(N__57912),
            .I(N__57885));
    Span4Mux_h I__10990 (
            .O(N__57907),
            .I(N__57885));
    Span4Mux_v I__10989 (
            .O(N__57902),
            .I(N__57885));
    Span4Mux_v I__10988 (
            .O(N__57899),
            .I(N__57885));
    Span4Mux_v I__10987 (
            .O(N__57896),
            .I(N__57882));
    Span4Mux_v I__10986 (
            .O(N__57885),
            .I(N__57879));
    Odrv4 I__10985 (
            .O(N__57882),
            .I(uart_drone_data_4));
    Odrv4 I__10984 (
            .O(N__57879),
            .I(uart_drone_data_4));
    InMux I__10983 (
            .O(N__57874),
            .I(N__57865));
    InMux I__10982 (
            .O(N__57873),
            .I(N__57862));
    InMux I__10981 (
            .O(N__57872),
            .I(N__57859));
    InMux I__10980 (
            .O(N__57871),
            .I(N__57856));
    InMux I__10979 (
            .O(N__57870),
            .I(N__57853));
    InMux I__10978 (
            .O(N__57869),
            .I(N__57850));
    InMux I__10977 (
            .O(N__57868),
            .I(N__57847));
    LocalMux I__10976 (
            .O(N__57865),
            .I(N__57844));
    LocalMux I__10975 (
            .O(N__57862),
            .I(N__57837));
    LocalMux I__10974 (
            .O(N__57859),
            .I(N__57837));
    LocalMux I__10973 (
            .O(N__57856),
            .I(N__57837));
    LocalMux I__10972 (
            .O(N__57853),
            .I(N__57834));
    LocalMux I__10971 (
            .O(N__57850),
            .I(N__57825));
    LocalMux I__10970 (
            .O(N__57847),
            .I(N__57825));
    Span4Mux_h I__10969 (
            .O(N__57844),
            .I(N__57825));
    Span4Mux_v I__10968 (
            .O(N__57837),
            .I(N__57825));
    Span4Mux_v I__10967 (
            .O(N__57834),
            .I(N__57822));
    Span4Mux_v I__10966 (
            .O(N__57825),
            .I(N__57819));
    Odrv4 I__10965 (
            .O(N__57822),
            .I(uart_drone_data_5));
    Odrv4 I__10964 (
            .O(N__57819),
            .I(uart_drone_data_5));
    InMux I__10963 (
            .O(N__57814),
            .I(N__57810));
    CascadeMux I__10962 (
            .O(N__57813),
            .I(N__57807));
    LocalMux I__10961 (
            .O(N__57810),
            .I(N__57804));
    InMux I__10960 (
            .O(N__57807),
            .I(N__57801));
    Span4Mux_h I__10959 (
            .O(N__57804),
            .I(N__57798));
    LocalMux I__10958 (
            .O(N__57801),
            .I(drone_H_disp_front_13));
    Odrv4 I__10957 (
            .O(N__57798),
            .I(drone_H_disp_front_13));
    CascadeMux I__10956 (
            .O(N__57793),
            .I(N__57786));
    InMux I__10955 (
            .O(N__57792),
            .I(N__57782));
    InMux I__10954 (
            .O(N__57791),
            .I(N__57778));
    InMux I__10953 (
            .O(N__57790),
            .I(N__57775));
    InMux I__10952 (
            .O(N__57789),
            .I(N__57772));
    InMux I__10951 (
            .O(N__57786),
            .I(N__57769));
    InMux I__10950 (
            .O(N__57785),
            .I(N__57766));
    LocalMux I__10949 (
            .O(N__57782),
            .I(N__57763));
    InMux I__10948 (
            .O(N__57781),
            .I(N__57760));
    LocalMux I__10947 (
            .O(N__57778),
            .I(N__57751));
    LocalMux I__10946 (
            .O(N__57775),
            .I(N__57751));
    LocalMux I__10945 (
            .O(N__57772),
            .I(N__57751));
    LocalMux I__10944 (
            .O(N__57769),
            .I(N__57751));
    LocalMux I__10943 (
            .O(N__57766),
            .I(N__57748));
    Span4Mux_h I__10942 (
            .O(N__57763),
            .I(N__57743));
    LocalMux I__10941 (
            .O(N__57760),
            .I(N__57743));
    Span12Mux_v I__10940 (
            .O(N__57751),
            .I(N__57740));
    Odrv12 I__10939 (
            .O(N__57748),
            .I(uart_drone_data_7));
    Odrv4 I__10938 (
            .O(N__57743),
            .I(uart_drone_data_7));
    Odrv12 I__10937 (
            .O(N__57740),
            .I(uart_drone_data_7));
    InMux I__10936 (
            .O(N__57733),
            .I(N__57730));
    LocalMux I__10935 (
            .O(N__57730),
            .I(drone_H_disp_front_15));
    InMux I__10934 (
            .O(N__57727),
            .I(N__57724));
    LocalMux I__10933 (
            .O(N__57724),
            .I(N__57718));
    InMux I__10932 (
            .O(N__57723),
            .I(N__57715));
    InMux I__10931 (
            .O(N__57722),
            .I(N__57712));
    InMux I__10930 (
            .O(N__57721),
            .I(N__57704));
    Span4Mux_v I__10929 (
            .O(N__57718),
            .I(N__57697));
    LocalMux I__10928 (
            .O(N__57715),
            .I(N__57697));
    LocalMux I__10927 (
            .O(N__57712),
            .I(N__57697));
    InMux I__10926 (
            .O(N__57711),
            .I(N__57694));
    InMux I__10925 (
            .O(N__57710),
            .I(N__57689));
    InMux I__10924 (
            .O(N__57709),
            .I(N__57689));
    InMux I__10923 (
            .O(N__57708),
            .I(N__57684));
    InMux I__10922 (
            .O(N__57707),
            .I(N__57684));
    LocalMux I__10921 (
            .O(N__57704),
            .I(N__57681));
    Span4Mux_v I__10920 (
            .O(N__57697),
            .I(N__57678));
    LocalMux I__10919 (
            .O(N__57694),
            .I(N__57669));
    LocalMux I__10918 (
            .O(N__57689),
            .I(N__57669));
    LocalMux I__10917 (
            .O(N__57684),
            .I(N__57669));
    Span12Mux_h I__10916 (
            .O(N__57681),
            .I(N__57669));
    Odrv4 I__10915 (
            .O(N__57678),
            .I(uart_drone_data_0));
    Odrv12 I__10914 (
            .O(N__57669),
            .I(uart_drone_data_0));
    InMux I__10913 (
            .O(N__57664),
            .I(N__57661));
    LocalMux I__10912 (
            .O(N__57661),
            .I(N__57658));
    Odrv12 I__10911 (
            .O(N__57658),
            .I(\dron_frame_decoder_1.drone_H_disp_front_8 ));
    CEMux I__10910 (
            .O(N__57655),
            .I(N__57652));
    LocalMux I__10909 (
            .O(N__57652),
            .I(N__57649));
    Span4Mux_v I__10908 (
            .O(N__57649),
            .I(N__57645));
    CEMux I__10907 (
            .O(N__57648),
            .I(N__57642));
    Span4Mux_v I__10906 (
            .O(N__57645),
            .I(N__57636));
    LocalMux I__10905 (
            .O(N__57642),
            .I(N__57636));
    CEMux I__10904 (
            .O(N__57641),
            .I(N__57633));
    Span4Mux_v I__10903 (
            .O(N__57636),
            .I(N__57630));
    LocalMux I__10902 (
            .O(N__57633),
            .I(N__57627));
    Span4Mux_h I__10901 (
            .O(N__57630),
            .I(N__57624));
    Span4Mux_h I__10900 (
            .O(N__57627),
            .I(N__57621));
    Odrv4 I__10899 (
            .O(N__57624),
            .I(\dron_frame_decoder_1.N_700_0 ));
    Odrv4 I__10898 (
            .O(N__57621),
            .I(\dron_frame_decoder_1.N_700_0 ));
    InMux I__10897 (
            .O(N__57616),
            .I(N__57613));
    LocalMux I__10896 (
            .O(N__57613),
            .I(N__57607));
    InMux I__10895 (
            .O(N__57612),
            .I(N__57604));
    InMux I__10894 (
            .O(N__57611),
            .I(N__57599));
    InMux I__10893 (
            .O(N__57610),
            .I(N__57599));
    Sp12to4 I__10892 (
            .O(N__57607),
            .I(N__57596));
    LocalMux I__10891 (
            .O(N__57604),
            .I(N__57591));
    LocalMux I__10890 (
            .O(N__57599),
            .I(N__57591));
    Span12Mux_v I__10889 (
            .O(N__57596),
            .I(N__57588));
    Span4Mux_v I__10888 (
            .O(N__57591),
            .I(N__57585));
    Odrv12 I__10887 (
            .O(N__57588),
            .I(\pid_alt.error_i_acumm_preregZ0Z_21 ));
    Odrv4 I__10886 (
            .O(N__57585),
            .I(\pid_alt.error_i_acumm_preregZ0Z_21 ));
    InMux I__10885 (
            .O(N__57580),
            .I(N__57577));
    LocalMux I__10884 (
            .O(N__57577),
            .I(N__57574));
    Span4Mux_h I__10883 (
            .O(N__57574),
            .I(N__57571));
    Span4Mux_h I__10882 (
            .O(N__57571),
            .I(N__57568));
    Span4Mux_h I__10881 (
            .O(N__57568),
            .I(N__57565));
    Odrv4 I__10880 (
            .O(N__57565),
            .I(\pid_alt.N_545 ));
    InMux I__10879 (
            .O(N__57562),
            .I(N__57559));
    LocalMux I__10878 (
            .O(N__57559),
            .I(N__57554));
    InMux I__10877 (
            .O(N__57558),
            .I(N__57549));
    InMux I__10876 (
            .O(N__57557),
            .I(N__57549));
    Odrv12 I__10875 (
            .O(N__57554),
            .I(\pid_alt.error_i_acumm7lto13 ));
    LocalMux I__10874 (
            .O(N__57549),
            .I(\pid_alt.error_i_acumm7lto13 ));
    InMux I__10873 (
            .O(N__57544),
            .I(N__57541));
    LocalMux I__10872 (
            .O(N__57541),
            .I(N__57538));
    Span4Mux_h I__10871 (
            .O(N__57538),
            .I(N__57535));
    Span4Mux_h I__10870 (
            .O(N__57535),
            .I(N__57532));
    Span4Mux_h I__10869 (
            .O(N__57532),
            .I(N__57529));
    Odrv4 I__10868 (
            .O(N__57529),
            .I(\pid_alt.error_i_acummZ0Z_13 ));
    CEMux I__10867 (
            .O(N__57526),
            .I(N__57523));
    LocalMux I__10866 (
            .O(N__57523),
            .I(N__57520));
    Span4Mux_v I__10865 (
            .O(N__57520),
            .I(N__57517));
    Span4Mux_h I__10864 (
            .O(N__57517),
            .I(N__57513));
    CEMux I__10863 (
            .O(N__57516),
            .I(N__57510));
    Span4Mux_h I__10862 (
            .O(N__57513),
            .I(N__57504));
    LocalMux I__10861 (
            .O(N__57510),
            .I(N__57504));
    CEMux I__10860 (
            .O(N__57509),
            .I(N__57501));
    Span4Mux_h I__10859 (
            .O(N__57504),
            .I(N__57498));
    LocalMux I__10858 (
            .O(N__57501),
            .I(N__57495));
    Odrv4 I__10857 (
            .O(N__57498),
            .I(\pid_alt.N_72_i_0 ));
    Odrv4 I__10856 (
            .O(N__57495),
            .I(\pid_alt.N_72_i_0 ));
    SRMux I__10855 (
            .O(N__57490),
            .I(N__57486));
    SRMux I__10854 (
            .O(N__57489),
            .I(N__57482));
    LocalMux I__10853 (
            .O(N__57486),
            .I(N__57479));
    SRMux I__10852 (
            .O(N__57485),
            .I(N__57475));
    LocalMux I__10851 (
            .O(N__57482),
            .I(N__57472));
    Span4Mux_v I__10850 (
            .O(N__57479),
            .I(N__57469));
    SRMux I__10849 (
            .O(N__57478),
            .I(N__57466));
    LocalMux I__10848 (
            .O(N__57475),
            .I(N__57463));
    Span4Mux_v I__10847 (
            .O(N__57472),
            .I(N__57460));
    Span4Mux_v I__10846 (
            .O(N__57469),
            .I(N__57457));
    LocalMux I__10845 (
            .O(N__57466),
            .I(N__57454));
    Span4Mux_h I__10844 (
            .O(N__57463),
            .I(N__57451));
    Span4Mux_h I__10843 (
            .O(N__57460),
            .I(N__57448));
    Span4Mux_h I__10842 (
            .O(N__57457),
            .I(N__57443));
    Span4Mux_h I__10841 (
            .O(N__57454),
            .I(N__57443));
    Odrv4 I__10840 (
            .O(N__57451),
            .I(\pid_alt.un1_reset_1_0_i ));
    Odrv4 I__10839 (
            .O(N__57448),
            .I(\pid_alt.un1_reset_1_0_i ));
    Odrv4 I__10838 (
            .O(N__57443),
            .I(\pid_alt.un1_reset_1_0_i ));
    InMux I__10837 (
            .O(N__57436),
            .I(N__57433));
    LocalMux I__10836 (
            .O(N__57433),
            .I(N__57430));
    Span4Mux_h I__10835 (
            .O(N__57430),
            .I(N__57427));
    Odrv4 I__10834 (
            .O(N__57427),
            .I(\pid_front.error_axb_8_l_ofx_0 ));
    InMux I__10833 (
            .O(N__57424),
            .I(N__57421));
    LocalMux I__10832 (
            .O(N__57421),
            .I(dron_frame_decoder_1_source_H_disp_front_fast_0));
    CEMux I__10831 (
            .O(N__57418),
            .I(N__57415));
    LocalMux I__10830 (
            .O(N__57415),
            .I(N__57409));
    CEMux I__10829 (
            .O(N__57414),
            .I(N__57406));
    CEMux I__10828 (
            .O(N__57413),
            .I(N__57403));
    CEMux I__10827 (
            .O(N__57412),
            .I(N__57400));
    Span4Mux_v I__10826 (
            .O(N__57409),
            .I(N__57396));
    LocalMux I__10825 (
            .O(N__57406),
            .I(N__57393));
    LocalMux I__10824 (
            .O(N__57403),
            .I(N__57390));
    LocalMux I__10823 (
            .O(N__57400),
            .I(N__57387));
    CEMux I__10822 (
            .O(N__57399),
            .I(N__57384));
    Span4Mux_h I__10821 (
            .O(N__57396),
            .I(N__57379));
    Span4Mux_h I__10820 (
            .O(N__57393),
            .I(N__57379));
    Span4Mux_v I__10819 (
            .O(N__57390),
            .I(N__57374));
    Span4Mux_h I__10818 (
            .O(N__57387),
            .I(N__57374));
    LocalMux I__10817 (
            .O(N__57384),
            .I(N__57371));
    Span4Mux_h I__10816 (
            .O(N__57379),
            .I(N__57368));
    Span4Mux_h I__10815 (
            .O(N__57374),
            .I(N__57365));
    Sp12to4 I__10814 (
            .O(N__57371),
            .I(N__57362));
    Span4Mux_h I__10813 (
            .O(N__57368),
            .I(N__57359));
    Span4Mux_h I__10812 (
            .O(N__57365),
            .I(N__57356));
    Odrv12 I__10811 (
            .O(N__57362),
            .I(\dron_frame_decoder_1.N_708_0 ));
    Odrv4 I__10810 (
            .O(N__57359),
            .I(\dron_frame_decoder_1.N_708_0 ));
    Odrv4 I__10809 (
            .O(N__57356),
            .I(\dron_frame_decoder_1.N_708_0 ));
    CascadeMux I__10808 (
            .O(N__57349),
            .I(\pid_front.N_510_cascade_ ));
    CascadeMux I__10807 (
            .O(N__57346),
            .I(\pid_front.N_596_cascade_ ));
    InMux I__10806 (
            .O(N__57343),
            .I(N__57340));
    LocalMux I__10805 (
            .O(N__57340),
            .I(N__57337));
    Span4Mux_h I__10804 (
            .O(N__57337),
            .I(N__57334));
    Odrv4 I__10803 (
            .O(N__57334),
            .I(\pid_front.m9_2_03_3_i_0_o2_1 ));
    CascadeMux I__10802 (
            .O(N__57331),
            .I(\pid_front.m9_2_03_3_i_3_cascade_ ));
    InMux I__10801 (
            .O(N__57328),
            .I(N__57322));
    InMux I__10800 (
            .O(N__57327),
            .I(N__57314));
    InMux I__10799 (
            .O(N__57326),
            .I(N__57311));
    InMux I__10798 (
            .O(N__57325),
            .I(N__57308));
    LocalMux I__10797 (
            .O(N__57322),
            .I(N__57305));
    InMux I__10796 (
            .O(N__57321),
            .I(N__57300));
    InMux I__10795 (
            .O(N__57320),
            .I(N__57300));
    InMux I__10794 (
            .O(N__57319),
            .I(N__57297));
    InMux I__10793 (
            .O(N__57318),
            .I(N__57294));
    InMux I__10792 (
            .O(N__57317),
            .I(N__57291));
    LocalMux I__10791 (
            .O(N__57314),
            .I(N__57288));
    LocalMux I__10790 (
            .O(N__57311),
            .I(N__57279));
    LocalMux I__10789 (
            .O(N__57308),
            .I(N__57279));
    Span4Mux_h I__10788 (
            .O(N__57305),
            .I(N__57279));
    LocalMux I__10787 (
            .O(N__57300),
            .I(N__57279));
    LocalMux I__10786 (
            .O(N__57297),
            .I(N__57276));
    LocalMux I__10785 (
            .O(N__57294),
            .I(N__57267));
    LocalMux I__10784 (
            .O(N__57291),
            .I(N__57267));
    Span4Mux_h I__10783 (
            .O(N__57288),
            .I(N__57267));
    Span4Mux_v I__10782 (
            .O(N__57279),
            .I(N__57267));
    Span4Mux_h I__10781 (
            .O(N__57276),
            .I(N__57264));
    Span4Mux_v I__10780 (
            .O(N__57267),
            .I(N__57261));
    Odrv4 I__10779 (
            .O(N__57264),
            .I(uart_drone_data_1));
    Odrv4 I__10778 (
            .O(N__57261),
            .I(uart_drone_data_1));
    InMux I__10777 (
            .O(N__57256),
            .I(N__57253));
    LocalMux I__10776 (
            .O(N__57253),
            .I(drone_H_disp_side_1));
    InMux I__10775 (
            .O(N__57250),
            .I(N__57245));
    InMux I__10774 (
            .O(N__57249),
            .I(N__57239));
    InMux I__10773 (
            .O(N__57248),
            .I(N__57236));
    LocalMux I__10772 (
            .O(N__57245),
            .I(N__57233));
    InMux I__10771 (
            .O(N__57244),
            .I(N__57230));
    InMux I__10770 (
            .O(N__57243),
            .I(N__57227));
    InMux I__10769 (
            .O(N__57242),
            .I(N__57223));
    LocalMux I__10768 (
            .O(N__57239),
            .I(N__57218));
    LocalMux I__10767 (
            .O(N__57236),
            .I(N__57218));
    Span4Mux_v I__10766 (
            .O(N__57233),
            .I(N__57213));
    LocalMux I__10765 (
            .O(N__57230),
            .I(N__57213));
    LocalMux I__10764 (
            .O(N__57227),
            .I(N__57210));
    InMux I__10763 (
            .O(N__57226),
            .I(N__57207));
    LocalMux I__10762 (
            .O(N__57223),
            .I(N__57202));
    Span4Mux_v I__10761 (
            .O(N__57218),
            .I(N__57202));
    Span4Mux_v I__10760 (
            .O(N__57213),
            .I(N__57199));
    Sp12to4 I__10759 (
            .O(N__57210),
            .I(N__57194));
    LocalMux I__10758 (
            .O(N__57207),
            .I(N__57194));
    Span4Mux_v I__10757 (
            .O(N__57202),
            .I(N__57191));
    Odrv4 I__10756 (
            .O(N__57199),
            .I(uart_drone_data_2));
    Odrv12 I__10755 (
            .O(N__57194),
            .I(uart_drone_data_2));
    Odrv4 I__10754 (
            .O(N__57191),
            .I(uart_drone_data_2));
    InMux I__10753 (
            .O(N__57184),
            .I(N__57181));
    LocalMux I__10752 (
            .O(N__57181),
            .I(drone_H_disp_side_2));
    InMux I__10751 (
            .O(N__57178),
            .I(N__57175));
    LocalMux I__10750 (
            .O(N__57175),
            .I(drone_H_disp_side_3));
    InMux I__10749 (
            .O(N__57172),
            .I(N__57169));
    LocalMux I__10748 (
            .O(N__57169),
            .I(\dron_frame_decoder_1.drone_H_disp_side_4 ));
    InMux I__10747 (
            .O(N__57166),
            .I(N__57163));
    LocalMux I__10746 (
            .O(N__57163),
            .I(\dron_frame_decoder_1.drone_H_disp_side_5 ));
    CascadeMux I__10745 (
            .O(N__57160),
            .I(N__57156));
    CascadeMux I__10744 (
            .O(N__57159),
            .I(N__57152));
    InMux I__10743 (
            .O(N__57156),
            .I(N__57144));
    InMux I__10742 (
            .O(N__57155),
            .I(N__57141));
    InMux I__10741 (
            .O(N__57152),
            .I(N__57138));
    InMux I__10740 (
            .O(N__57151),
            .I(N__57134));
    InMux I__10739 (
            .O(N__57150),
            .I(N__57131));
    InMux I__10738 (
            .O(N__57149),
            .I(N__57128));
    InMux I__10737 (
            .O(N__57148),
            .I(N__57125));
    InMux I__10736 (
            .O(N__57147),
            .I(N__57122));
    LocalMux I__10735 (
            .O(N__57144),
            .I(N__57115));
    LocalMux I__10734 (
            .O(N__57141),
            .I(N__57115));
    LocalMux I__10733 (
            .O(N__57138),
            .I(N__57115));
    InMux I__10732 (
            .O(N__57137),
            .I(N__57112));
    LocalMux I__10731 (
            .O(N__57134),
            .I(N__57109));
    LocalMux I__10730 (
            .O(N__57131),
            .I(N__57106));
    LocalMux I__10729 (
            .O(N__57128),
            .I(N__57097));
    LocalMux I__10728 (
            .O(N__57125),
            .I(N__57097));
    LocalMux I__10727 (
            .O(N__57122),
            .I(N__57097));
    Span4Mux_h I__10726 (
            .O(N__57115),
            .I(N__57097));
    LocalMux I__10725 (
            .O(N__57112),
            .I(N__57088));
    Span4Mux_h I__10724 (
            .O(N__57109),
            .I(N__57088));
    Span4Mux_h I__10723 (
            .O(N__57106),
            .I(N__57088));
    Span4Mux_v I__10722 (
            .O(N__57097),
            .I(N__57088));
    Span4Mux_v I__10721 (
            .O(N__57088),
            .I(N__57085));
    Odrv4 I__10720 (
            .O(N__57085),
            .I(uart_drone_data_6));
    InMux I__10719 (
            .O(N__57082),
            .I(N__57079));
    LocalMux I__10718 (
            .O(N__57079),
            .I(\dron_frame_decoder_1.drone_H_disp_side_6 ));
    CEMux I__10717 (
            .O(N__57076),
            .I(N__57073));
    LocalMux I__10716 (
            .O(N__57073),
            .I(N__57069));
    CEMux I__10715 (
            .O(N__57072),
            .I(N__57066));
    Span4Mux_h I__10714 (
            .O(N__57069),
            .I(N__57063));
    LocalMux I__10713 (
            .O(N__57066),
            .I(N__57060));
    Span4Mux_h I__10712 (
            .O(N__57063),
            .I(N__57057));
    Odrv4 I__10711 (
            .O(N__57060),
            .I(\dron_frame_decoder_1.N_724_0 ));
    Odrv4 I__10710 (
            .O(N__57057),
            .I(\dron_frame_decoder_1.N_724_0 ));
    CascadeMux I__10709 (
            .O(N__57052),
            .I(\pid_side.error_i_reg_esr_RNO_6Z0Z_12_cascade_ ));
    InMux I__10708 (
            .O(N__57049),
            .I(N__57046));
    LocalMux I__10707 (
            .O(N__57046),
            .I(\dron_frame_decoder_1.drone_H_disp_front_7 ));
    InMux I__10706 (
            .O(N__57043),
            .I(N__57040));
    LocalMux I__10705 (
            .O(N__57040),
            .I(N__57037));
    Odrv4 I__10704 (
            .O(N__57037),
            .I(drone_H_disp_front_i_7));
    CascadeMux I__10703 (
            .O(N__57034),
            .I(N__57031));
    InMux I__10702 (
            .O(N__57031),
            .I(N__57028));
    LocalMux I__10701 (
            .O(N__57028),
            .I(N__57025));
    Odrv4 I__10700 (
            .O(N__57025),
            .I(drone_H_disp_front_i_8));
    InMux I__10699 (
            .O(N__57022),
            .I(N__57019));
    LocalMux I__10698 (
            .O(N__57019),
            .I(\dron_frame_decoder_1.drone_H_disp_front_9 ));
    InMux I__10697 (
            .O(N__57016),
            .I(N__57013));
    LocalMux I__10696 (
            .O(N__57013),
            .I(N__57010));
    Odrv4 I__10695 (
            .O(N__57010),
            .I(drone_H_disp_front_i_9));
    InMux I__10694 (
            .O(N__57007),
            .I(N__57004));
    LocalMux I__10693 (
            .O(N__57004),
            .I(N__57000));
    InMux I__10692 (
            .O(N__57003),
            .I(N__56997));
    Odrv4 I__10691 (
            .O(N__57000),
            .I(\uart_drone.data_AuxZ0Z_6 ));
    LocalMux I__10690 (
            .O(N__56997),
            .I(\uart_drone.data_AuxZ0Z_6 ));
    InMux I__10689 (
            .O(N__56992),
            .I(N__56988));
    CascadeMux I__10688 (
            .O(N__56991),
            .I(N__56985));
    LocalMux I__10687 (
            .O(N__56988),
            .I(N__56982));
    InMux I__10686 (
            .O(N__56985),
            .I(N__56979));
    Odrv4 I__10685 (
            .O(N__56982),
            .I(\uart_drone.data_AuxZ0Z_7 ));
    LocalMux I__10684 (
            .O(N__56979),
            .I(\uart_drone.data_AuxZ0Z_7 ));
    CEMux I__10683 (
            .O(N__56974),
            .I(N__56971));
    LocalMux I__10682 (
            .O(N__56971),
            .I(N__56968));
    Span4Mux_v I__10681 (
            .O(N__56968),
            .I(N__56965));
    Span4Mux_h I__10680 (
            .O(N__56965),
            .I(N__56962));
    Span4Mux_h I__10679 (
            .O(N__56962),
            .I(N__56959));
    Odrv4 I__10678 (
            .O(N__56959),
            .I(\uart_drone.data_rdyc_1_0 ));
    SRMux I__10677 (
            .O(N__56956),
            .I(N__56953));
    LocalMux I__10676 (
            .O(N__56953),
            .I(N__56950));
    Span4Mux_v I__10675 (
            .O(N__56950),
            .I(N__56946));
    InMux I__10674 (
            .O(N__56949),
            .I(N__56943));
    Odrv4 I__10673 (
            .O(N__56946),
            .I(\uart_drone.timer_Count_RNIES9Q1Z0Z_2 ));
    LocalMux I__10672 (
            .O(N__56943),
            .I(\uart_drone.timer_Count_RNIES9Q1Z0Z_2 ));
    InMux I__10671 (
            .O(N__56938),
            .I(N__56935));
    LocalMux I__10670 (
            .O(N__56935),
            .I(\pid_front.error_cry_2_c_RNIFP8GZ0Z1 ));
    CascadeMux I__10669 (
            .O(N__56932),
            .I(\pid_front.m26_2_03_0_m2_ns_1_cascade_ ));
    CascadeMux I__10668 (
            .O(N__56929),
            .I(\pid_front.m27_2_03_0_0_cascade_ ));
    InMux I__10667 (
            .O(N__56926),
            .I(N__56923));
    LocalMux I__10666 (
            .O(N__56923),
            .I(\pid_front.N_253 ));
    InMux I__10665 (
            .O(N__56920),
            .I(N__56917));
    LocalMux I__10664 (
            .O(N__56917),
            .I(N__56914));
    Span4Mux_h I__10663 (
            .O(N__56914),
            .I(N__56911));
    Odrv4 I__10662 (
            .O(N__56911),
            .I(\uart_drone.data_Auxce_0_6 ));
    InMux I__10661 (
            .O(N__56908),
            .I(N__56884));
    InMux I__10660 (
            .O(N__56907),
            .I(N__56884));
    InMux I__10659 (
            .O(N__56906),
            .I(N__56884));
    InMux I__10658 (
            .O(N__56905),
            .I(N__56884));
    InMux I__10657 (
            .O(N__56904),
            .I(N__56884));
    InMux I__10656 (
            .O(N__56903),
            .I(N__56884));
    InMux I__10655 (
            .O(N__56902),
            .I(N__56884));
    InMux I__10654 (
            .O(N__56901),
            .I(N__56884));
    LocalMux I__10653 (
            .O(N__56884),
            .I(N__56881));
    Odrv4 I__10652 (
            .O(N__56881),
            .I(\uart_drone.un1_state_2_0 ));
    IoInMux I__10651 (
            .O(N__56878),
            .I(N__56873));
    InMux I__10650 (
            .O(N__56877),
            .I(N__56870));
    CascadeMux I__10649 (
            .O(N__56876),
            .I(N__56863));
    LocalMux I__10648 (
            .O(N__56873),
            .I(N__56859));
    LocalMux I__10647 (
            .O(N__56870),
            .I(N__56856));
    CascadeMux I__10646 (
            .O(N__56869),
            .I(N__56849));
    CascadeMux I__10645 (
            .O(N__56868),
            .I(N__56846));
    CascadeMux I__10644 (
            .O(N__56867),
            .I(N__56843));
    CascadeMux I__10643 (
            .O(N__56866),
            .I(N__56840));
    InMux I__10642 (
            .O(N__56863),
            .I(N__56837));
    InMux I__10641 (
            .O(N__56862),
            .I(N__56834));
    Span4Mux_s3_v I__10640 (
            .O(N__56859),
            .I(N__56831));
    Span4Mux_h I__10639 (
            .O(N__56856),
            .I(N__56828));
    InMux I__10638 (
            .O(N__56855),
            .I(N__56810));
    InMux I__10637 (
            .O(N__56854),
            .I(N__56810));
    InMux I__10636 (
            .O(N__56853),
            .I(N__56810));
    InMux I__10635 (
            .O(N__56852),
            .I(N__56810));
    InMux I__10634 (
            .O(N__56849),
            .I(N__56810));
    InMux I__10633 (
            .O(N__56846),
            .I(N__56810));
    InMux I__10632 (
            .O(N__56843),
            .I(N__56810));
    InMux I__10631 (
            .O(N__56840),
            .I(N__56810));
    LocalMux I__10630 (
            .O(N__56837),
            .I(N__56805));
    LocalMux I__10629 (
            .O(N__56834),
            .I(N__56805));
    Span4Mux_v I__10628 (
            .O(N__56831),
            .I(N__56802));
    Span4Mux_v I__10627 (
            .O(N__56828),
            .I(N__56799));
    InMux I__10626 (
            .O(N__56827),
            .I(N__56795));
    LocalMux I__10625 (
            .O(N__56810),
            .I(N__56792));
    Span4Mux_v I__10624 (
            .O(N__56805),
            .I(N__56789));
    Span4Mux_h I__10623 (
            .O(N__56802),
            .I(N__56784));
    Span4Mux_v I__10622 (
            .O(N__56799),
            .I(N__56784));
    InMux I__10621 (
            .O(N__56798),
            .I(N__56781));
    LocalMux I__10620 (
            .O(N__56795),
            .I(debug_CH0_16A_c));
    Odrv4 I__10619 (
            .O(N__56792),
            .I(debug_CH0_16A_c));
    Odrv4 I__10618 (
            .O(N__56789),
            .I(debug_CH0_16A_c));
    Odrv4 I__10617 (
            .O(N__56784),
            .I(debug_CH0_16A_c));
    LocalMux I__10616 (
            .O(N__56781),
            .I(debug_CH0_16A_c));
    CascadeMux I__10615 (
            .O(N__56770),
            .I(N__56766));
    InMux I__10614 (
            .O(N__56769),
            .I(N__56763));
    InMux I__10613 (
            .O(N__56766),
            .I(N__56760));
    LocalMux I__10612 (
            .O(N__56763),
            .I(N__56757));
    LocalMux I__10611 (
            .O(N__56760),
            .I(N__56751));
    Span4Mux_v I__10610 (
            .O(N__56757),
            .I(N__56751));
    InMux I__10609 (
            .O(N__56756),
            .I(N__56748));
    Odrv4 I__10608 (
            .O(N__56751),
            .I(\uart_drone.N_152 ));
    LocalMux I__10607 (
            .O(N__56748),
            .I(\uart_drone.N_152 ));
    SRMux I__10606 (
            .O(N__56743),
            .I(N__56740));
    LocalMux I__10605 (
            .O(N__56740),
            .I(N__56737));
    Span4Mux_v I__10604 (
            .O(N__56737),
            .I(N__56734));
    Odrv4 I__10603 (
            .O(N__56734),
            .I(\uart_drone.state_RNIOU0NZ0Z_4 ));
    InMux I__10602 (
            .O(N__56731),
            .I(N__56728));
    LocalMux I__10601 (
            .O(N__56728),
            .I(N__56724));
    InMux I__10600 (
            .O(N__56727),
            .I(N__56721));
    Odrv4 I__10599 (
            .O(N__56724),
            .I(\uart_drone.data_AuxZ0Z_0 ));
    LocalMux I__10598 (
            .O(N__56721),
            .I(\uart_drone.data_AuxZ0Z_0 ));
    InMux I__10597 (
            .O(N__56716),
            .I(N__56712));
    CascadeMux I__10596 (
            .O(N__56715),
            .I(N__56709));
    LocalMux I__10595 (
            .O(N__56712),
            .I(N__56706));
    InMux I__10594 (
            .O(N__56709),
            .I(N__56703));
    Odrv4 I__10593 (
            .O(N__56706),
            .I(\uart_drone.data_AuxZ0Z_1 ));
    LocalMux I__10592 (
            .O(N__56703),
            .I(\uart_drone.data_AuxZ0Z_1 ));
    InMux I__10591 (
            .O(N__56698),
            .I(N__56695));
    LocalMux I__10590 (
            .O(N__56695),
            .I(N__56691));
    InMux I__10589 (
            .O(N__56694),
            .I(N__56688));
    Odrv4 I__10588 (
            .O(N__56691),
            .I(\uart_drone.data_AuxZ0Z_2 ));
    LocalMux I__10587 (
            .O(N__56688),
            .I(\uart_drone.data_AuxZ0Z_2 ));
    InMux I__10586 (
            .O(N__56683),
            .I(N__56679));
    CascadeMux I__10585 (
            .O(N__56682),
            .I(N__56676));
    LocalMux I__10584 (
            .O(N__56679),
            .I(N__56673));
    InMux I__10583 (
            .O(N__56676),
            .I(N__56670));
    Odrv4 I__10582 (
            .O(N__56673),
            .I(\uart_drone.data_AuxZ0Z_3 ));
    LocalMux I__10581 (
            .O(N__56670),
            .I(\uart_drone.data_AuxZ0Z_3 ));
    InMux I__10580 (
            .O(N__56665),
            .I(N__56662));
    LocalMux I__10579 (
            .O(N__56662),
            .I(N__56658));
    InMux I__10578 (
            .O(N__56661),
            .I(N__56655));
    Odrv4 I__10577 (
            .O(N__56658),
            .I(\uart_drone.data_AuxZ0Z_4 ));
    LocalMux I__10576 (
            .O(N__56655),
            .I(\uart_drone.data_AuxZ0Z_4 ));
    InMux I__10575 (
            .O(N__56650),
            .I(N__56646));
    CascadeMux I__10574 (
            .O(N__56649),
            .I(N__56643));
    LocalMux I__10573 (
            .O(N__56646),
            .I(N__56640));
    InMux I__10572 (
            .O(N__56643),
            .I(N__56637));
    Odrv4 I__10571 (
            .O(N__56640),
            .I(\uart_drone.data_AuxZ0Z_5 ));
    LocalMux I__10570 (
            .O(N__56637),
            .I(\uart_drone.data_AuxZ0Z_5 ));
    InMux I__10569 (
            .O(N__56632),
            .I(N__56623));
    InMux I__10568 (
            .O(N__56631),
            .I(N__56623));
    InMux I__10567 (
            .O(N__56630),
            .I(N__56623));
    LocalMux I__10566 (
            .O(N__56623),
            .I(N__56617));
    InMux I__10565 (
            .O(N__56622),
            .I(N__56612));
    InMux I__10564 (
            .O(N__56621),
            .I(N__56612));
    CascadeMux I__10563 (
            .O(N__56620),
            .I(N__56607));
    Span4Mux_v I__10562 (
            .O(N__56617),
            .I(N__56601));
    LocalMux I__10561 (
            .O(N__56612),
            .I(N__56601));
    InMux I__10560 (
            .O(N__56611),
            .I(N__56596));
    InMux I__10559 (
            .O(N__56610),
            .I(N__56596));
    InMux I__10558 (
            .O(N__56607),
            .I(N__56589));
    InMux I__10557 (
            .O(N__56606),
            .I(N__56589));
    Span4Mux_h I__10556 (
            .O(N__56601),
            .I(N__56586));
    LocalMux I__10555 (
            .O(N__56596),
            .I(N__56583));
    InMux I__10554 (
            .O(N__56595),
            .I(N__56578));
    InMux I__10553 (
            .O(N__56594),
            .I(N__56578));
    LocalMux I__10552 (
            .O(N__56589),
            .I(\uart_drone.bit_CountZ0Z_0 ));
    Odrv4 I__10551 (
            .O(N__56586),
            .I(\uart_drone.bit_CountZ0Z_0 ));
    Odrv12 I__10550 (
            .O(N__56583),
            .I(\uart_drone.bit_CountZ0Z_0 ));
    LocalMux I__10549 (
            .O(N__56578),
            .I(\uart_drone.bit_CountZ0Z_0 ));
    CascadeMux I__10548 (
            .O(N__56569),
            .I(N__56566));
    InMux I__10547 (
            .O(N__56566),
            .I(N__56557));
    InMux I__10546 (
            .O(N__56565),
            .I(N__56557));
    InMux I__10545 (
            .O(N__56564),
            .I(N__56557));
    LocalMux I__10544 (
            .O(N__56557),
            .I(N__56551));
    InMux I__10543 (
            .O(N__56556),
            .I(N__56546));
    InMux I__10542 (
            .O(N__56555),
            .I(N__56546));
    CascadeMux I__10541 (
            .O(N__56554),
            .I(N__56540));
    Span4Mux_v I__10540 (
            .O(N__56551),
            .I(N__56534));
    LocalMux I__10539 (
            .O(N__56546),
            .I(N__56534));
    InMux I__10538 (
            .O(N__56545),
            .I(N__56529));
    InMux I__10537 (
            .O(N__56544),
            .I(N__56529));
    CascadeMux I__10536 (
            .O(N__56543),
            .I(N__56526));
    InMux I__10535 (
            .O(N__56540),
            .I(N__56521));
    InMux I__10534 (
            .O(N__56539),
            .I(N__56521));
    Span4Mux_h I__10533 (
            .O(N__56534),
            .I(N__56518));
    LocalMux I__10532 (
            .O(N__56529),
            .I(N__56515));
    InMux I__10531 (
            .O(N__56526),
            .I(N__56512));
    LocalMux I__10530 (
            .O(N__56521),
            .I(\uart_drone.bit_CountZ0Z_1 ));
    Odrv4 I__10529 (
            .O(N__56518),
            .I(\uart_drone.bit_CountZ0Z_1 ));
    Odrv12 I__10528 (
            .O(N__56515),
            .I(\uart_drone.bit_CountZ0Z_1 ));
    LocalMux I__10527 (
            .O(N__56512),
            .I(\uart_drone.bit_CountZ0Z_1 ));
    InMux I__10526 (
            .O(N__56503),
            .I(N__56494));
    InMux I__10525 (
            .O(N__56502),
            .I(N__56494));
    InMux I__10524 (
            .O(N__56501),
            .I(N__56494));
    LocalMux I__10523 (
            .O(N__56494),
            .I(N__56488));
    InMux I__10522 (
            .O(N__56493),
            .I(N__56483));
    InMux I__10521 (
            .O(N__56492),
            .I(N__56483));
    CascadeMux I__10520 (
            .O(N__56491),
            .I(N__56480));
    Span4Mux_v I__10519 (
            .O(N__56488),
            .I(N__56473));
    LocalMux I__10518 (
            .O(N__56483),
            .I(N__56473));
    InMux I__10517 (
            .O(N__56480),
            .I(N__56468));
    InMux I__10516 (
            .O(N__56479),
            .I(N__56468));
    InMux I__10515 (
            .O(N__56478),
            .I(N__56464));
    Span4Mux_h I__10514 (
            .O(N__56473),
            .I(N__56461));
    LocalMux I__10513 (
            .O(N__56468),
            .I(N__56458));
    InMux I__10512 (
            .O(N__56467),
            .I(N__56455));
    LocalMux I__10511 (
            .O(N__56464),
            .I(\uart_drone.bit_CountZ0Z_2 ));
    Odrv4 I__10510 (
            .O(N__56461),
            .I(\uart_drone.bit_CountZ0Z_2 ));
    Odrv12 I__10509 (
            .O(N__56458),
            .I(\uart_drone.bit_CountZ0Z_2 ));
    LocalMux I__10508 (
            .O(N__56455),
            .I(\uart_drone.bit_CountZ0Z_2 ));
    InMux I__10507 (
            .O(N__56446),
            .I(N__56443));
    LocalMux I__10506 (
            .O(N__56443),
            .I(\uart_drone.data_Auxce_0_0_0 ));
    InMux I__10505 (
            .O(N__56440),
            .I(N__56437));
    LocalMux I__10504 (
            .O(N__56437),
            .I(\uart_drone.data_Auxce_0_1 ));
    InMux I__10503 (
            .O(N__56434),
            .I(N__56431));
    LocalMux I__10502 (
            .O(N__56431),
            .I(N__56428));
    Odrv12 I__10501 (
            .O(N__56428),
            .I(\uart_drone.data_Auxce_0_0_2 ));
    InMux I__10500 (
            .O(N__56425),
            .I(N__56422));
    LocalMux I__10499 (
            .O(N__56422),
            .I(N__56419));
    Odrv4 I__10498 (
            .O(N__56419),
            .I(\uart_drone.data_Auxce_0_3 ));
    InMux I__10497 (
            .O(N__56416),
            .I(N__56413));
    LocalMux I__10496 (
            .O(N__56413),
            .I(N__56410));
    Odrv12 I__10495 (
            .O(N__56410),
            .I(\uart_drone.data_Auxce_0_0_4 ));
    InMux I__10494 (
            .O(N__56407),
            .I(N__56404));
    LocalMux I__10493 (
            .O(N__56404),
            .I(\uart_drone.data_Auxce_0_5 ));
    InMux I__10492 (
            .O(N__56401),
            .I(N__56398));
    LocalMux I__10491 (
            .O(N__56398),
            .I(N__56395));
    Span4Mux_h I__10490 (
            .O(N__56395),
            .I(N__56391));
    InMux I__10489 (
            .O(N__56394),
            .I(N__56388));
    Odrv4 I__10488 (
            .O(N__56391),
            .I(\pid_side.N_603 ));
    LocalMux I__10487 (
            .O(N__56388),
            .I(\pid_side.N_603 ));
    CascadeMux I__10486 (
            .O(N__56383),
            .I(\pid_side.N_181_cascade_ ));
    CascadeMux I__10485 (
            .O(N__56380),
            .I(\pid_side.error_i_acumm_13_i_0_1_3_cascade_ ));
    CascadeMux I__10484 (
            .O(N__56377),
            .I(\pid_side.error_i_acumm_13_i_0_3_cascade_ ));
    InMux I__10483 (
            .O(N__56374),
            .I(N__56368));
    InMux I__10482 (
            .O(N__56373),
            .I(N__56368));
    LocalMux I__10481 (
            .O(N__56368),
            .I(N__56365));
    Odrv4 I__10480 (
            .O(N__56365),
            .I(\pid_side.N_177 ));
    InMux I__10479 (
            .O(N__56362),
            .I(N__56359));
    LocalMux I__10478 (
            .O(N__56359),
            .I(\pid_side.N_544 ));
    CascadeMux I__10477 (
            .O(N__56356),
            .I(\pid_side.N_233_cascade_ ));
    CascadeMux I__10476 (
            .O(N__56353),
            .I(\pid_side.N_251_cascade_ ));
    CascadeMux I__10475 (
            .O(N__56350),
            .I(\pid_side.N_531_cascade_ ));
    CascadeMux I__10474 (
            .O(N__56347),
            .I(\pid_side.N_544_cascade_ ));
    IoInMux I__10473 (
            .O(N__56344),
            .I(N__56341));
    LocalMux I__10472 (
            .O(N__56341),
            .I(N__56338));
    IoSpan4Mux I__10471 (
            .O(N__56338),
            .I(N__56335));
    Span4Mux_s1_v I__10470 (
            .O(N__56335),
            .I(N__56332));
    Odrv4 I__10469 (
            .O(N__56332),
            .I(\pid_side.state_0_0 ));
    CascadeMux I__10468 (
            .O(N__56329),
            .I(\pid_side.source_pid_9_i_0_o3_0_11_cascade_ ));
    CascadeMux I__10467 (
            .O(N__56326),
            .I(N__56320));
    CascadeMux I__10466 (
            .O(N__56325),
            .I(N__56317));
    CascadeMux I__10465 (
            .O(N__56324),
            .I(N__56313));
    CascadeMux I__10464 (
            .O(N__56323),
            .I(N__56310));
    InMux I__10463 (
            .O(N__56320),
            .I(N__56284));
    InMux I__10462 (
            .O(N__56317),
            .I(N__56284));
    InMux I__10461 (
            .O(N__56316),
            .I(N__56284));
    InMux I__10460 (
            .O(N__56313),
            .I(N__56284));
    InMux I__10459 (
            .O(N__56310),
            .I(N__56284));
    InMux I__10458 (
            .O(N__56309),
            .I(N__56284));
    InMux I__10457 (
            .O(N__56308),
            .I(N__56275));
    InMux I__10456 (
            .O(N__56307),
            .I(N__56275));
    InMux I__10455 (
            .O(N__56306),
            .I(N__56275));
    InMux I__10454 (
            .O(N__56305),
            .I(N__56275));
    InMux I__10453 (
            .O(N__56304),
            .I(N__56271));
    InMux I__10452 (
            .O(N__56303),
            .I(N__56262));
    InMux I__10451 (
            .O(N__56302),
            .I(N__56262));
    InMux I__10450 (
            .O(N__56301),
            .I(N__56262));
    InMux I__10449 (
            .O(N__56300),
            .I(N__56255));
    InMux I__10448 (
            .O(N__56299),
            .I(N__56255));
    InMux I__10447 (
            .O(N__56298),
            .I(N__56255));
    InMux I__10446 (
            .O(N__56297),
            .I(N__56252));
    LocalMux I__10445 (
            .O(N__56284),
            .I(N__56246));
    LocalMux I__10444 (
            .O(N__56275),
            .I(N__56246));
    InMux I__10443 (
            .O(N__56274),
            .I(N__56243));
    LocalMux I__10442 (
            .O(N__56271),
            .I(N__56233));
    InMux I__10441 (
            .O(N__56270),
            .I(N__56228));
    InMux I__10440 (
            .O(N__56269),
            .I(N__56228));
    LocalMux I__10439 (
            .O(N__56262),
            .I(N__56225));
    LocalMux I__10438 (
            .O(N__56255),
            .I(N__56220));
    LocalMux I__10437 (
            .O(N__56252),
            .I(N__56220));
    CascadeMux I__10436 (
            .O(N__56251),
            .I(N__56217));
    Span4Mux_s2_v I__10435 (
            .O(N__56246),
            .I(N__56212));
    LocalMux I__10434 (
            .O(N__56243),
            .I(N__56209));
    InMux I__10433 (
            .O(N__56242),
            .I(N__56206));
    InMux I__10432 (
            .O(N__56241),
            .I(N__56193));
    InMux I__10431 (
            .O(N__56240),
            .I(N__56193));
    InMux I__10430 (
            .O(N__56239),
            .I(N__56193));
    InMux I__10429 (
            .O(N__56238),
            .I(N__56193));
    InMux I__10428 (
            .O(N__56237),
            .I(N__56193));
    InMux I__10427 (
            .O(N__56236),
            .I(N__56193));
    Span4Mux_h I__10426 (
            .O(N__56233),
            .I(N__56190));
    LocalMux I__10425 (
            .O(N__56228),
            .I(N__56185));
    Span4Mux_h I__10424 (
            .O(N__56225),
            .I(N__56185));
    Span4Mux_h I__10423 (
            .O(N__56220),
            .I(N__56182));
    InMux I__10422 (
            .O(N__56217),
            .I(N__56175));
    InMux I__10421 (
            .O(N__56216),
            .I(N__56175));
    InMux I__10420 (
            .O(N__56215),
            .I(N__56175));
    Span4Mux_v I__10419 (
            .O(N__56212),
            .I(N__56172));
    Span4Mux_h I__10418 (
            .O(N__56209),
            .I(N__56169));
    LocalMux I__10417 (
            .O(N__56206),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    LocalMux I__10416 (
            .O(N__56193),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    Odrv4 I__10415 (
            .O(N__56190),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    Odrv4 I__10414 (
            .O(N__56185),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    Odrv4 I__10413 (
            .O(N__56182),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    LocalMux I__10412 (
            .O(N__56175),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    Odrv4 I__10411 (
            .O(N__56172),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    Odrv4 I__10410 (
            .O(N__56169),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    InMux I__10409 (
            .O(N__56152),
            .I(N__56149));
    LocalMux I__10408 (
            .O(N__56149),
            .I(N__56146));
    Span4Mux_h I__10407 (
            .O(N__56146),
            .I(N__56143));
    Odrv4 I__10406 (
            .O(N__56143),
            .I(\ppm_encoder_1.N_267_i ));
    CascadeMux I__10405 (
            .O(N__56140),
            .I(N__56137));
    InMux I__10404 (
            .O(N__56137),
            .I(N__56134));
    LocalMux I__10403 (
            .O(N__56134),
            .I(N__56131));
    Span4Mux_v I__10402 (
            .O(N__56131),
            .I(N__56128));
    Odrv4 I__10401 (
            .O(N__56128),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_12_1 ));
    InMux I__10400 (
            .O(N__56125),
            .I(N__56122));
    LocalMux I__10399 (
            .O(N__56122),
            .I(N__56119));
    Span4Mux_h I__10398 (
            .O(N__56119),
            .I(N__56116));
    Span4Mux_h I__10397 (
            .O(N__56116),
            .I(N__56113));
    Odrv4 I__10396 (
            .O(N__56113),
            .I(\ppm_encoder_1.un2_throttle_iv_0_2_12 ));
    CascadeMux I__10395 (
            .O(N__56110),
            .I(N__56107));
    InMux I__10394 (
            .O(N__56107),
            .I(N__56104));
    LocalMux I__10393 (
            .O(N__56104),
            .I(N__56101));
    Span4Mux_v I__10392 (
            .O(N__56101),
            .I(N__56097));
    InMux I__10391 (
            .O(N__56100),
            .I(N__56094));
    Sp12to4 I__10390 (
            .O(N__56097),
            .I(N__56089));
    LocalMux I__10389 (
            .O(N__56094),
            .I(N__56089));
    Odrv12 I__10388 (
            .O(N__56089),
            .I(\ppm_encoder_1.N_267_i_i ));
    CascadeMux I__10387 (
            .O(N__56086),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_12_cascade_ ));
    InMux I__10386 (
            .O(N__56083),
            .I(N__56080));
    LocalMux I__10385 (
            .O(N__56080),
            .I(N__56077));
    Span4Mux_h I__10384 (
            .O(N__56077),
            .I(N__56074));
    Odrv4 I__10383 (
            .O(N__56074),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_RNI1TA86Z0Z_2 ));
    CascadeMux I__10382 (
            .O(N__56071),
            .I(\pid_side.error_i_acumm_13_i_o2_0_7_3_cascade_ ));
    CascadeMux I__10381 (
            .O(N__56068),
            .I(\pid_side.un1_reset_i_a2_4_cascade_ ));
    CascadeMux I__10380 (
            .O(N__56065),
            .I(\pid_side.N_342_cascade_ ));
    CascadeMux I__10379 (
            .O(N__56062),
            .I(\pid_side.un1_reset_0_i_3_cascade_ ));
    InMux I__10378 (
            .O(N__56059),
            .I(N__56056));
    LocalMux I__10377 (
            .O(N__56056),
            .I(N__56052));
    InMux I__10376 (
            .O(N__56055),
            .I(N__56049));
    Span4Mux_v I__10375 (
            .O(N__56052),
            .I(N__56044));
    LocalMux I__10374 (
            .O(N__56049),
            .I(N__56044));
    Span4Mux_h I__10373 (
            .O(N__56044),
            .I(N__56041));
    Span4Mux_v I__10372 (
            .O(N__56041),
            .I(N__56038));
    Odrv4 I__10371 (
            .O(N__56038),
            .I(side_order_1));
    InMux I__10370 (
            .O(N__56035),
            .I(N__56032));
    LocalMux I__10369 (
            .O(N__56032),
            .I(N__56028));
    InMux I__10368 (
            .O(N__56031),
            .I(N__56025));
    Span4Mux_h I__10367 (
            .O(N__56028),
            .I(N__56022));
    LocalMux I__10366 (
            .O(N__56025),
            .I(N__56019));
    Span4Mux_h I__10365 (
            .O(N__56022),
            .I(N__56016));
    Span12Mux_h I__10364 (
            .O(N__56019),
            .I(N__56013));
    Odrv4 I__10363 (
            .O(N__56016),
            .I(side_order_2));
    Odrv12 I__10362 (
            .O(N__56013),
            .I(side_order_2));
    InMux I__10361 (
            .O(N__56008),
            .I(N__56005));
    LocalMux I__10360 (
            .O(N__56005),
            .I(N__56001));
    InMux I__10359 (
            .O(N__56004),
            .I(N__55998));
    Span4Mux_h I__10358 (
            .O(N__56001),
            .I(N__55995));
    LocalMux I__10357 (
            .O(N__55998),
            .I(N__55992));
    Span4Mux_v I__10356 (
            .O(N__55995),
            .I(N__55989));
    Span12Mux_v I__10355 (
            .O(N__55992),
            .I(N__55986));
    Odrv4 I__10354 (
            .O(N__55989),
            .I(side_order_3));
    Odrv12 I__10353 (
            .O(N__55986),
            .I(side_order_3));
    CascadeMux I__10352 (
            .O(N__55981),
            .I(\pid_front.error_d_reg_prev_esr_RNIQHN6Z0Z_1_cascade_ ));
    CascadeMux I__10351 (
            .O(N__55978),
            .I(\pid_front.error_p_reg_esr_RNI2BC9_0Z0Z_1_cascade_ ));
    InMux I__10350 (
            .O(N__55975),
            .I(N__55972));
    LocalMux I__10349 (
            .O(N__55972),
            .I(\pid_front.error_p_reg_esr_RNI2BC9Z0Z_1 ));
    InMux I__10348 (
            .O(N__55969),
            .I(N__55966));
    LocalMux I__10347 (
            .O(N__55966),
            .I(N__55963));
    Span12Mux_h I__10346 (
            .O(N__55963),
            .I(N__55960));
    Span12Mux_v I__10345 (
            .O(N__55960),
            .I(N__55957));
    Odrv12 I__10344 (
            .O(N__55957),
            .I(\pid_front.O_0_10 ));
    CascadeMux I__10343 (
            .O(N__55954),
            .I(\pid_front.un1_pid_prereg_0_10_cascade_ ));
    InMux I__10342 (
            .O(N__55951),
            .I(N__55947));
    InMux I__10341 (
            .O(N__55950),
            .I(N__55944));
    LocalMux I__10340 (
            .O(N__55947),
            .I(\pid_front.un1_pid_prereg_0_8 ));
    LocalMux I__10339 (
            .O(N__55944),
            .I(\pid_front.un1_pid_prereg_0_8 ));
    CascadeMux I__10338 (
            .O(N__55939),
            .I(\pid_front.un1_pid_prereg_0_8_cascade_ ));
    InMux I__10337 (
            .O(N__55936),
            .I(N__55930));
    InMux I__10336 (
            .O(N__55935),
            .I(N__55930));
    LocalMux I__10335 (
            .O(N__55930),
            .I(\pid_front.un1_pid_prereg_0_9 ));
    InMux I__10334 (
            .O(N__55927),
            .I(N__55923));
    InMux I__10333 (
            .O(N__55926),
            .I(N__55920));
    LocalMux I__10332 (
            .O(N__55923),
            .I(N__55917));
    LocalMux I__10331 (
            .O(N__55920),
            .I(N__55914));
    Span4Mux_h I__10330 (
            .O(N__55917),
            .I(N__55909));
    Span4Mux_h I__10329 (
            .O(N__55914),
            .I(N__55909));
    Odrv4 I__10328 (
            .O(N__55909),
            .I(\pid_front.un11lto30_i_a2_5_and ));
    InMux I__10327 (
            .O(N__55906),
            .I(N__55903));
    LocalMux I__10326 (
            .O(N__55903),
            .I(N__55900));
    Odrv4 I__10325 (
            .O(N__55900),
            .I(\pid_front.N_2364_i ));
    CascadeMux I__10324 (
            .O(N__55897),
            .I(N__55894));
    InMux I__10323 (
            .O(N__55894),
            .I(N__55890));
    InMux I__10322 (
            .O(N__55893),
            .I(N__55887));
    LocalMux I__10321 (
            .O(N__55890),
            .I(N__55884));
    LocalMux I__10320 (
            .O(N__55887),
            .I(N__55881));
    Span4Mux_h I__10319 (
            .O(N__55884),
            .I(N__55878));
    Span4Mux_v I__10318 (
            .O(N__55881),
            .I(N__55875));
    Span4Mux_h I__10317 (
            .O(N__55878),
            .I(N__55872));
    Span4Mux_v I__10316 (
            .O(N__55875),
            .I(N__55869));
    Span4Mux_v I__10315 (
            .O(N__55872),
            .I(N__55866));
    Sp12to4 I__10314 (
            .O(N__55869),
            .I(N__55863));
    Span4Mux_v I__10313 (
            .O(N__55866),
            .I(N__55860));
    Odrv12 I__10312 (
            .O(N__55863),
            .I(\pid_front.error_p_regZ0Z_7 ));
    Odrv4 I__10311 (
            .O(N__55860),
            .I(\pid_front.error_p_regZ0Z_7 ));
    CascadeMux I__10310 (
            .O(N__55855),
            .I(\pid_front.error_p_reg_esr_RNIBG6F_0Z0Z_7_cascade_ ));
    InMux I__10309 (
            .O(N__55852),
            .I(N__55848));
    CascadeMux I__10308 (
            .O(N__55851),
            .I(N__55845));
    LocalMux I__10307 (
            .O(N__55848),
            .I(N__55842));
    InMux I__10306 (
            .O(N__55845),
            .I(N__55839));
    Sp12to4 I__10305 (
            .O(N__55842),
            .I(N__55834));
    LocalMux I__10304 (
            .O(N__55839),
            .I(N__55834));
    Odrv12 I__10303 (
            .O(N__55834),
            .I(\pid_front.un11lto30_i_a2_6_and ));
    CascadeMux I__10302 (
            .O(N__55831),
            .I(\pid_front.error_p_reg_esr_RNIGL6FZ0Z_8_cascade_ ));
    InMux I__10301 (
            .O(N__55828),
            .I(N__55824));
    InMux I__10300 (
            .O(N__55827),
            .I(N__55821));
    LocalMux I__10299 (
            .O(N__55824),
            .I(N__55818));
    LocalMux I__10298 (
            .O(N__55821),
            .I(N__55815));
    Span4Mux_h I__10297 (
            .O(N__55818),
            .I(N__55812));
    Odrv4 I__10296 (
            .O(N__55815),
            .I(\pid_front.un11lto30_i_a2_3_and ));
    Odrv4 I__10295 (
            .O(N__55812),
            .I(\pid_front.un11lto30_i_a2_3_and ));
    InMux I__10294 (
            .O(N__55807),
            .I(N__55804));
    LocalMux I__10293 (
            .O(N__55804),
            .I(N__55801));
    Odrv4 I__10292 (
            .O(N__55801),
            .I(\pid_front.un11lto30_i_a2_2_and ));
    InMux I__10291 (
            .O(N__55798),
            .I(N__55795));
    LocalMux I__10290 (
            .O(N__55795),
            .I(N__55789));
    InMux I__10289 (
            .O(N__55794),
            .I(N__55782));
    InMux I__10288 (
            .O(N__55793),
            .I(N__55782));
    InMux I__10287 (
            .O(N__55792),
            .I(N__55782));
    Odrv4 I__10286 (
            .O(N__55789),
            .I(\pid_front.pid_preregZ0Z_14 ));
    LocalMux I__10285 (
            .O(N__55782),
            .I(\pid_front.pid_preregZ0Z_14 ));
    InMux I__10284 (
            .O(N__55777),
            .I(N__55774));
    LocalMux I__10283 (
            .O(N__55774),
            .I(\pid_front.source_pid_9_i_0_o3_0_11 ));
    CascadeMux I__10282 (
            .O(N__55771),
            .I(\pid_front.source_pid_9_i_0_o3_0_11_cascade_ ));
    InMux I__10281 (
            .O(N__55768),
            .I(N__55765));
    LocalMux I__10280 (
            .O(N__55765),
            .I(N__55761));
    InMux I__10279 (
            .O(N__55764),
            .I(N__55758));
    Odrv4 I__10278 (
            .O(N__55761),
            .I(\pid_front.N_175 ));
    LocalMux I__10277 (
            .O(N__55758),
            .I(\pid_front.N_175 ));
    CascadeMux I__10276 (
            .O(N__55753),
            .I(\pid_front.un1_pid_prereg_0_9_cascade_ ));
    InMux I__10275 (
            .O(N__55750),
            .I(N__55747));
    LocalMux I__10274 (
            .O(N__55747),
            .I(N__55744));
    Span4Mux_v I__10273 (
            .O(N__55744),
            .I(N__55740));
    InMux I__10272 (
            .O(N__55743),
            .I(N__55737));
    Span4Mux_v I__10271 (
            .O(N__55740),
            .I(N__55734));
    LocalMux I__10270 (
            .O(N__55737),
            .I(N__55731));
    Span4Mux_v I__10269 (
            .O(N__55734),
            .I(N__55728));
    Span12Mux_s9_v I__10268 (
            .O(N__55731),
            .I(N__55725));
    Span4Mux_h I__10267 (
            .O(N__55728),
            .I(N__55722));
    Span12Mux_v I__10266 (
            .O(N__55725),
            .I(N__55719));
    Odrv4 I__10265 (
            .O(N__55722),
            .I(front_order_13));
    Odrv12 I__10264 (
            .O(N__55719),
            .I(front_order_13));
    InMux I__10263 (
            .O(N__55714),
            .I(N__55708));
    InMux I__10262 (
            .O(N__55713),
            .I(N__55708));
    LocalMux I__10261 (
            .O(N__55708),
            .I(\pid_front.N_277 ));
    InMux I__10260 (
            .O(N__55705),
            .I(N__55702));
    LocalMux I__10259 (
            .O(N__55702),
            .I(N__55698));
    InMux I__10258 (
            .O(N__55701),
            .I(N__55695));
    Span4Mux_h I__10257 (
            .O(N__55698),
            .I(N__55692));
    LocalMux I__10256 (
            .O(N__55695),
            .I(N__55689));
    Span4Mux_h I__10255 (
            .O(N__55692),
            .I(N__55686));
    Span4Mux_v I__10254 (
            .O(N__55689),
            .I(N__55683));
    Sp12to4 I__10253 (
            .O(N__55686),
            .I(N__55680));
    Span4Mux_v I__10252 (
            .O(N__55683),
            .I(N__55677));
    Span12Mux_s9_v I__10251 (
            .O(N__55680),
            .I(N__55674));
    Span4Mux_v I__10250 (
            .O(N__55677),
            .I(N__55671));
    Span12Mux_v I__10249 (
            .O(N__55674),
            .I(N__55668));
    Span4Mux_v I__10248 (
            .O(N__55671),
            .I(N__55665));
    Odrv12 I__10247 (
            .O(N__55668),
            .I(front_order_12));
    Odrv4 I__10246 (
            .O(N__55665),
            .I(front_order_12));
    CascadeMux I__10245 (
            .O(N__55660),
            .I(\pid_front.N_2364_i_cascade_ ));
    InMux I__10244 (
            .O(N__55657),
            .I(N__55654));
    LocalMux I__10243 (
            .O(N__55654),
            .I(\pid_front.error_p_reg_esr_RNIBG6FZ0Z_7 ));
    InMux I__10242 (
            .O(N__55651),
            .I(N__55645));
    InMux I__10241 (
            .O(N__55650),
            .I(N__55645));
    LocalMux I__10240 (
            .O(N__55645),
            .I(\pid_front.error_p_reg_esr_RNIGL6F_0Z0Z_8 ));
    CascadeMux I__10239 (
            .O(N__55642),
            .I(\pid_front.error_p_reg_esr_RNIBG6FZ0Z_7_cascade_ ));
    CascadeMux I__10238 (
            .O(N__55639),
            .I(N__55635));
    InMux I__10237 (
            .O(N__55638),
            .I(N__55627));
    InMux I__10236 (
            .O(N__55635),
            .I(N__55627));
    InMux I__10235 (
            .O(N__55634),
            .I(N__55627));
    LocalMux I__10234 (
            .O(N__55627),
            .I(\pid_front.error_d_reg_prevZ0Z_7 ));
    CascadeMux I__10233 (
            .O(N__55624),
            .I(N__55621));
    InMux I__10232 (
            .O(N__55621),
            .I(N__55615));
    InMux I__10231 (
            .O(N__55620),
            .I(N__55615));
    LocalMux I__10230 (
            .O(N__55615),
            .I(N__55612));
    Span4Mux_v I__10229 (
            .O(N__55612),
            .I(N__55609));
    Span4Mux_h I__10228 (
            .O(N__55609),
            .I(N__55606));
    Span4Mux_v I__10227 (
            .O(N__55606),
            .I(N__55603));
    Odrv4 I__10226 (
            .O(N__55603),
            .I(\pid_front.error_p_regZ0Z_8 ));
    CEMux I__10225 (
            .O(N__55600),
            .I(N__55597));
    LocalMux I__10224 (
            .O(N__55597),
            .I(N__55594));
    Span4Mux_v I__10223 (
            .O(N__55594),
            .I(N__55591));
    Span4Mux_h I__10222 (
            .O(N__55591),
            .I(N__55588));
    Span4Mux_h I__10221 (
            .O(N__55588),
            .I(N__55585));
    Odrv4 I__10220 (
            .O(N__55585),
            .I(\Commands_frame_decoder.source_CH3data_1_sqmuxa_0 ));
    InMux I__10219 (
            .O(N__55582),
            .I(N__55576));
    InMux I__10218 (
            .O(N__55581),
            .I(N__55576));
    LocalMux I__10217 (
            .O(N__55576),
            .I(N__55573));
    Odrv4 I__10216 (
            .O(N__55573),
            .I(drone_H_disp_front_14));
    InMux I__10215 (
            .O(N__55570),
            .I(N__55567));
    LocalMux I__10214 (
            .O(N__55567),
            .I(N__55564));
    Span4Mux_h I__10213 (
            .O(N__55564),
            .I(N__55561));
    Odrv4 I__10212 (
            .O(N__55561),
            .I(\dron_frame_decoder_1.drone_H_disp_front_10 ));
    InMux I__10211 (
            .O(N__55558),
            .I(N__55554));
    InMux I__10210 (
            .O(N__55557),
            .I(N__55551));
    LocalMux I__10209 (
            .O(N__55554),
            .I(N__55548));
    LocalMux I__10208 (
            .O(N__55551),
            .I(N__55545));
    Odrv4 I__10207 (
            .O(N__55548),
            .I(\pid_front.un11lto30_i_a2_4_and ));
    Odrv4 I__10206 (
            .O(N__55545),
            .I(\pid_front.un11lto30_i_a2_4_and ));
    CascadeMux I__10205 (
            .O(N__55540),
            .I(\pid_front.N_175_cascade_ ));
    CascadeMux I__10204 (
            .O(N__55537),
            .I(N__55534));
    InMux I__10203 (
            .O(N__55534),
            .I(N__55530));
    InMux I__10202 (
            .O(N__55533),
            .I(N__55527));
    LocalMux I__10201 (
            .O(N__55530),
            .I(N__55522));
    LocalMux I__10200 (
            .O(N__55527),
            .I(N__55522));
    Odrv4 I__10199 (
            .O(N__55522),
            .I(\pid_front.N_593 ));
    CascadeMux I__10198 (
            .O(N__55519),
            .I(\pid_front.N_277_cascade_ ));
    InMux I__10197 (
            .O(N__55516),
            .I(N__55513));
    LocalMux I__10196 (
            .O(N__55513),
            .I(\pid_front.N_291 ));
    CascadeMux I__10195 (
            .O(N__55510),
            .I(\pid_front.un1_reset_i_o3_0_cascade_ ));
    InMux I__10194 (
            .O(N__55507),
            .I(N__55504));
    LocalMux I__10193 (
            .O(N__55504),
            .I(\pid_front.N_342 ));
    CascadeMux I__10192 (
            .O(N__55501),
            .I(\pid_front.un1_reset_0_i_3_cascade_ ));
    CascadeMux I__10191 (
            .O(N__55498),
            .I(N__55495));
    InMux I__10190 (
            .O(N__55495),
            .I(N__55492));
    LocalMux I__10189 (
            .O(N__55492),
            .I(drone_H_disp_front_i_13));
    InMux I__10188 (
            .O(N__55489),
            .I(\pid_front.error_cry_9 ));
    InMux I__10187 (
            .O(N__55486),
            .I(\pid_front.error_cry_10 ));
    CascadeMux I__10186 (
            .O(N__55483),
            .I(N__55480));
    InMux I__10185 (
            .O(N__55480),
            .I(N__55477));
    LocalMux I__10184 (
            .O(N__55477),
            .I(N__55474));
    Odrv4 I__10183 (
            .O(N__55474),
            .I(front_command_0));
    CascadeMux I__10182 (
            .O(N__55471),
            .I(N__55468));
    InMux I__10181 (
            .O(N__55468),
            .I(N__55465));
    LocalMux I__10180 (
            .O(N__55465),
            .I(N__55462));
    Odrv4 I__10179 (
            .O(N__55462),
            .I(front_command_1));
    CascadeMux I__10178 (
            .O(N__55459),
            .I(N__55456));
    InMux I__10177 (
            .O(N__55456),
            .I(N__55453));
    LocalMux I__10176 (
            .O(N__55453),
            .I(N__55450));
    Odrv4 I__10175 (
            .O(N__55450),
            .I(front_command_2));
    CascadeMux I__10174 (
            .O(N__55447),
            .I(N__55444));
    InMux I__10173 (
            .O(N__55444),
            .I(N__55441));
    LocalMux I__10172 (
            .O(N__55441),
            .I(N__55438));
    Odrv4 I__10171 (
            .O(N__55438),
            .I(front_command_3));
    InMux I__10170 (
            .O(N__55435),
            .I(N__55432));
    LocalMux I__10169 (
            .O(N__55432),
            .I(front_command_4));
    CascadeMux I__10168 (
            .O(N__55429),
            .I(N__55426));
    InMux I__10167 (
            .O(N__55426),
            .I(N__55423));
    LocalMux I__10166 (
            .O(N__55423),
            .I(front_command_5));
    CascadeMux I__10165 (
            .O(N__55420),
            .I(N__55417));
    InMux I__10164 (
            .O(N__55417),
            .I(N__55414));
    LocalMux I__10163 (
            .O(N__55414),
            .I(N__55411));
    Odrv4 I__10162 (
            .O(N__55411),
            .I(front_command_6));
    InMux I__10161 (
            .O(N__55408),
            .I(N__55405));
    LocalMux I__10160 (
            .O(N__55405),
            .I(drone_H_disp_front_i_5));
    InMux I__10159 (
            .O(N__55402),
            .I(\pid_front.error_cry_0_0 ));
    InMux I__10158 (
            .O(N__55399),
            .I(N__55396));
    LocalMux I__10157 (
            .O(N__55396),
            .I(drone_H_disp_front_i_6));
    InMux I__10156 (
            .O(N__55393),
            .I(\pid_front.error_cry_1_0 ));
    InMux I__10155 (
            .O(N__55390),
            .I(\pid_front.error_cry_2_0 ));
    InMux I__10154 (
            .O(N__55387),
            .I(bfn_12_19_0_));
    InMux I__10153 (
            .O(N__55384),
            .I(\pid_front.error_cry_4 ));
    InMux I__10152 (
            .O(N__55381),
            .I(N__55378));
    LocalMux I__10151 (
            .O(N__55378),
            .I(drone_H_disp_front_i_10));
    InMux I__10150 (
            .O(N__55375),
            .I(\pid_front.error_cry_5 ));
    InMux I__10149 (
            .O(N__55372),
            .I(\pid_front.error_cry_6 ));
    InMux I__10148 (
            .O(N__55369),
            .I(\pid_front.error_cry_7 ));
    InMux I__10147 (
            .O(N__55366),
            .I(\pid_front.error_cry_8 ));
    InMux I__10146 (
            .O(N__55363),
            .I(N__55360));
    LocalMux I__10145 (
            .O(N__55360),
            .I(drone_H_disp_front_2));
    InMux I__10144 (
            .O(N__55357),
            .I(N__55354));
    LocalMux I__10143 (
            .O(N__55354),
            .I(N__55351));
    Odrv4 I__10142 (
            .O(N__55351),
            .I(\dron_frame_decoder_1.drone_H_disp_front_4 ));
    InMux I__10141 (
            .O(N__55348),
            .I(N__55345));
    LocalMux I__10140 (
            .O(N__55345),
            .I(\pid_front.error_axb_0 ));
    InMux I__10139 (
            .O(N__55342),
            .I(N__55339));
    LocalMux I__10138 (
            .O(N__55339),
            .I(\pid_front.error_axbZ0Z_1 ));
    InMux I__10137 (
            .O(N__55336),
            .I(\pid_front.error_cry_0 ));
    InMux I__10136 (
            .O(N__55333),
            .I(N__55330));
    LocalMux I__10135 (
            .O(N__55330),
            .I(\pid_front.error_axbZ0Z_2 ));
    InMux I__10134 (
            .O(N__55327),
            .I(\pid_front.error_cry_1 ));
    InMux I__10133 (
            .O(N__55324),
            .I(N__55321));
    LocalMux I__10132 (
            .O(N__55321),
            .I(\pid_front.error_axbZ0Z_3 ));
    InMux I__10131 (
            .O(N__55318),
            .I(\pid_front.error_cry_2 ));
    InMux I__10130 (
            .O(N__55315),
            .I(N__55312));
    LocalMux I__10129 (
            .O(N__55312),
            .I(drone_H_disp_front_i_4));
    InMux I__10128 (
            .O(N__55309),
            .I(\pid_front.error_cry_3 ));
    CascadeMux I__10127 (
            .O(N__55306),
            .I(\pid_front.m64_i_o2_0_cascade_ ));
    CascadeMux I__10126 (
            .O(N__55303),
            .I(\pid_front.error_i_reg_esr_RNO_4_0_14_cascade_ ));
    InMux I__10125 (
            .O(N__55300),
            .I(N__55297));
    LocalMux I__10124 (
            .O(N__55297),
            .I(\pid_front.m64_i_o2_0 ));
    CascadeMux I__10123 (
            .O(N__55294),
            .I(\pid_front.m9_2_03_3_i_0_o2_0_1_cascade_ ));
    CascadeMux I__10122 (
            .O(N__55291),
            .I(\pid_front.m9_2_03_3_i_0_o2_0_cascade_ ));
    InMux I__10121 (
            .O(N__55288),
            .I(N__55285));
    LocalMux I__10120 (
            .O(N__55285),
            .I(drone_H_disp_front_3));
    InMux I__10119 (
            .O(N__55282),
            .I(N__55273));
    InMux I__10118 (
            .O(N__55281),
            .I(N__55273));
    InMux I__10117 (
            .O(N__55280),
            .I(N__55270));
    InMux I__10116 (
            .O(N__55279),
            .I(N__55264));
    InMux I__10115 (
            .O(N__55278),
            .I(N__55259));
    LocalMux I__10114 (
            .O(N__55273),
            .I(N__55248));
    LocalMux I__10113 (
            .O(N__55270),
            .I(N__55248));
    CascadeMux I__10112 (
            .O(N__55269),
            .I(N__55244));
    InMux I__10111 (
            .O(N__55268),
            .I(N__55235));
    InMux I__10110 (
            .O(N__55267),
            .I(N__55235));
    LocalMux I__10109 (
            .O(N__55264),
            .I(N__55231));
    InMux I__10108 (
            .O(N__55263),
            .I(N__55228));
    InMux I__10107 (
            .O(N__55262),
            .I(N__55225));
    LocalMux I__10106 (
            .O(N__55259),
            .I(N__55222));
    InMux I__10105 (
            .O(N__55258),
            .I(N__55219));
    InMux I__10104 (
            .O(N__55257),
            .I(N__55212));
    InMux I__10103 (
            .O(N__55256),
            .I(N__55212));
    InMux I__10102 (
            .O(N__55255),
            .I(N__55212));
    InMux I__10101 (
            .O(N__55254),
            .I(N__55209));
    InMux I__10100 (
            .O(N__55253),
            .I(N__55202));
    Span4Mux_v I__10099 (
            .O(N__55248),
            .I(N__55199));
    InMux I__10098 (
            .O(N__55247),
            .I(N__55186));
    InMux I__10097 (
            .O(N__55244),
            .I(N__55186));
    InMux I__10096 (
            .O(N__55243),
            .I(N__55186));
    InMux I__10095 (
            .O(N__55242),
            .I(N__55186));
    InMux I__10094 (
            .O(N__55241),
            .I(N__55186));
    InMux I__10093 (
            .O(N__55240),
            .I(N__55186));
    LocalMux I__10092 (
            .O(N__55235),
            .I(N__55183));
    InMux I__10091 (
            .O(N__55234),
            .I(N__55180));
    Span4Mux_v I__10090 (
            .O(N__55231),
            .I(N__55175));
    LocalMux I__10089 (
            .O(N__55228),
            .I(N__55175));
    LocalMux I__10088 (
            .O(N__55225),
            .I(N__55168));
    Span4Mux_h I__10087 (
            .O(N__55222),
            .I(N__55168));
    LocalMux I__10086 (
            .O(N__55219),
            .I(N__55168));
    LocalMux I__10085 (
            .O(N__55212),
            .I(N__55165));
    LocalMux I__10084 (
            .O(N__55209),
            .I(N__55162));
    CascadeMux I__10083 (
            .O(N__55208),
            .I(N__55159));
    InMux I__10082 (
            .O(N__55207),
            .I(N__55150));
    InMux I__10081 (
            .O(N__55206),
            .I(N__55150));
    InMux I__10080 (
            .O(N__55205),
            .I(N__55150));
    LocalMux I__10079 (
            .O(N__55202),
            .I(N__55147));
    Span4Mux_h I__10078 (
            .O(N__55199),
            .I(N__55144));
    LocalMux I__10077 (
            .O(N__55186),
            .I(N__55135));
    Span4Mux_h I__10076 (
            .O(N__55183),
            .I(N__55135));
    LocalMux I__10075 (
            .O(N__55180),
            .I(N__55135));
    Span4Mux_h I__10074 (
            .O(N__55175),
            .I(N__55135));
    Span4Mux_v I__10073 (
            .O(N__55168),
            .I(N__55128));
    Span4Mux_v I__10072 (
            .O(N__55165),
            .I(N__55128));
    Span4Mux_h I__10071 (
            .O(N__55162),
            .I(N__55128));
    InMux I__10070 (
            .O(N__55159),
            .I(N__55121));
    InMux I__10069 (
            .O(N__55158),
            .I(N__55121));
    InMux I__10068 (
            .O(N__55157),
            .I(N__55121));
    LocalMux I__10067 (
            .O(N__55150),
            .I(N__55118));
    Odrv12 I__10066 (
            .O(N__55147),
            .I(uart_pc_data_rdy));
    Odrv4 I__10065 (
            .O(N__55144),
            .I(uart_pc_data_rdy));
    Odrv4 I__10064 (
            .O(N__55135),
            .I(uart_pc_data_rdy));
    Odrv4 I__10063 (
            .O(N__55128),
            .I(uart_pc_data_rdy));
    LocalMux I__10062 (
            .O(N__55121),
            .I(uart_pc_data_rdy));
    Odrv12 I__10061 (
            .O(N__55118),
            .I(uart_pc_data_rdy));
    SRMux I__10060 (
            .O(N__55105),
            .I(N__55102));
    LocalMux I__10059 (
            .O(N__55102),
            .I(N__55098));
    SRMux I__10058 (
            .O(N__55101),
            .I(N__55095));
    Span4Mux_v I__10057 (
            .O(N__55098),
            .I(N__55092));
    LocalMux I__10056 (
            .O(N__55095),
            .I(N__55089));
    Odrv4 I__10055 (
            .O(N__55092),
            .I(\Commands_frame_decoder.un1_state57_iZ0 ));
    Odrv12 I__10054 (
            .O(N__55089),
            .I(\Commands_frame_decoder.un1_state57_iZ0 ));
    CascadeMux I__10053 (
            .O(N__55084),
            .I(\pid_side.state_RNINK4UZ0Z_0_cascade_ ));
    InMux I__10052 (
            .O(N__55081),
            .I(N__55077));
    InMux I__10051 (
            .O(N__55080),
            .I(N__55074));
    LocalMux I__10050 (
            .O(N__55077),
            .I(\reset_module_System.countZ0Z_19 ));
    LocalMux I__10049 (
            .O(N__55074),
            .I(\reset_module_System.countZ0Z_19 ));
    InMux I__10048 (
            .O(N__55069),
            .I(N__55065));
    InMux I__10047 (
            .O(N__55068),
            .I(N__55062));
    LocalMux I__10046 (
            .O(N__55065),
            .I(\reset_module_System.countZ0Z_15 ));
    LocalMux I__10045 (
            .O(N__55062),
            .I(\reset_module_System.countZ0Z_15 ));
    CascadeMux I__10044 (
            .O(N__55057),
            .I(N__55053));
    InMux I__10043 (
            .O(N__55056),
            .I(N__55050));
    InMux I__10042 (
            .O(N__55053),
            .I(N__55047));
    LocalMux I__10041 (
            .O(N__55050),
            .I(\reset_module_System.countZ0Z_21 ));
    LocalMux I__10040 (
            .O(N__55047),
            .I(\reset_module_System.countZ0Z_21 ));
    InMux I__10039 (
            .O(N__55042),
            .I(N__55038));
    InMux I__10038 (
            .O(N__55041),
            .I(N__55035));
    LocalMux I__10037 (
            .O(N__55038),
            .I(\reset_module_System.countZ0Z_13 ));
    LocalMux I__10036 (
            .O(N__55035),
            .I(\reset_module_System.countZ0Z_13 ));
    InMux I__10035 (
            .O(N__55030),
            .I(N__55019));
    InMux I__10034 (
            .O(N__55029),
            .I(N__55019));
    InMux I__10033 (
            .O(N__55028),
            .I(N__55019));
    InMux I__10032 (
            .O(N__55027),
            .I(N__55014));
    InMux I__10031 (
            .O(N__55026),
            .I(N__55014));
    LocalMux I__10030 (
            .O(N__55019),
            .I(N__55011));
    LocalMux I__10029 (
            .O(N__55014),
            .I(N__55008));
    Span4Mux_h I__10028 (
            .O(N__55011),
            .I(N__55005));
    Odrv12 I__10027 (
            .O(N__55008),
            .I(\reset_module_System.reset6_15 ));
    Odrv4 I__10026 (
            .O(N__55005),
            .I(\reset_module_System.reset6_15 ));
    InMux I__10025 (
            .O(N__55000),
            .I(N__54997));
    LocalMux I__10024 (
            .O(N__54997),
            .I(N__54993));
    InMux I__10023 (
            .O(N__54996),
            .I(N__54990));
    Span4Mux_v I__10022 (
            .O(N__54993),
            .I(N__54985));
    LocalMux I__10021 (
            .O(N__54990),
            .I(N__54985));
    Span4Mux_h I__10020 (
            .O(N__54985),
            .I(N__54982));
    Odrv4 I__10019 (
            .O(N__54982),
            .I(front_order_1));
    InMux I__10018 (
            .O(N__54979),
            .I(N__54976));
    LocalMux I__10017 (
            .O(N__54976),
            .I(N__54972));
    InMux I__10016 (
            .O(N__54975),
            .I(N__54969));
    Span4Mux_h I__10015 (
            .O(N__54972),
            .I(N__54966));
    LocalMux I__10014 (
            .O(N__54969),
            .I(N__54963));
    Span4Mux_v I__10013 (
            .O(N__54966),
            .I(N__54960));
    Span4Mux_h I__10012 (
            .O(N__54963),
            .I(N__54957));
    Odrv4 I__10011 (
            .O(N__54960),
            .I(front_order_4));
    Odrv4 I__10010 (
            .O(N__54957),
            .I(front_order_4));
    InMux I__10009 (
            .O(N__54952),
            .I(N__54949));
    LocalMux I__10008 (
            .O(N__54949),
            .I(\reset_module_System.count_1_2 ));
    CascadeMux I__10007 (
            .O(N__54946),
            .I(N__54942));
    CascadeMux I__10006 (
            .O(N__54945),
            .I(N__54937));
    InMux I__10005 (
            .O(N__54942),
            .I(N__54931));
    InMux I__10004 (
            .O(N__54941),
            .I(N__54931));
    InMux I__10003 (
            .O(N__54940),
            .I(N__54924));
    InMux I__10002 (
            .O(N__54937),
            .I(N__54924));
    InMux I__10001 (
            .O(N__54936),
            .I(N__54924));
    LocalMux I__10000 (
            .O(N__54931),
            .I(\reset_module_System.reset6_14 ));
    LocalMux I__9999 (
            .O(N__54924),
            .I(\reset_module_System.reset6_14 ));
    InMux I__9998 (
            .O(N__54919),
            .I(N__54913));
    InMux I__9997 (
            .O(N__54918),
            .I(N__54908));
    InMux I__9996 (
            .O(N__54917),
            .I(N__54908));
    InMux I__9995 (
            .O(N__54916),
            .I(N__54905));
    LocalMux I__9994 (
            .O(N__54913),
            .I(\reset_module_System.reset6_19 ));
    LocalMux I__9993 (
            .O(N__54908),
            .I(\reset_module_System.reset6_19 ));
    LocalMux I__9992 (
            .O(N__54905),
            .I(\reset_module_System.reset6_19 ));
    InMux I__9991 (
            .O(N__54898),
            .I(N__54894));
    InMux I__9990 (
            .O(N__54897),
            .I(N__54891));
    LocalMux I__9989 (
            .O(N__54894),
            .I(N__54888));
    LocalMux I__9988 (
            .O(N__54891),
            .I(\reset_module_System.countZ0Z_6 ));
    Odrv4 I__9987 (
            .O(N__54888),
            .I(\reset_module_System.countZ0Z_6 ));
    InMux I__9986 (
            .O(N__54883),
            .I(N__54879));
    InMux I__9985 (
            .O(N__54882),
            .I(N__54876));
    LocalMux I__9984 (
            .O(N__54879),
            .I(N__54871));
    LocalMux I__9983 (
            .O(N__54876),
            .I(N__54871));
    Odrv4 I__9982 (
            .O(N__54871),
            .I(\reset_module_System.countZ0Z_3 ));
    CascadeMux I__9981 (
            .O(N__54868),
            .I(N__54865));
    InMux I__9980 (
            .O(N__54865),
            .I(N__54861));
    InMux I__9979 (
            .O(N__54864),
            .I(N__54858));
    LocalMux I__9978 (
            .O(N__54861),
            .I(N__54855));
    LocalMux I__9977 (
            .O(N__54858),
            .I(\reset_module_System.countZ0Z_20 ));
    Odrv4 I__9976 (
            .O(N__54855),
            .I(\reset_module_System.countZ0Z_20 ));
    InMux I__9975 (
            .O(N__54850),
            .I(N__54846));
    InMux I__9974 (
            .O(N__54849),
            .I(N__54843));
    LocalMux I__9973 (
            .O(N__54846),
            .I(N__54840));
    LocalMux I__9972 (
            .O(N__54843),
            .I(\reset_module_System.countZ0Z_2 ));
    Odrv4 I__9971 (
            .O(N__54840),
            .I(\reset_module_System.countZ0Z_2 ));
    InMux I__9970 (
            .O(N__54835),
            .I(N__54832));
    LocalMux I__9969 (
            .O(N__54832),
            .I(\reset_module_System.reset6_11 ));
    InMux I__9968 (
            .O(N__54829),
            .I(N__54826));
    LocalMux I__9967 (
            .O(N__54826),
            .I(\pid_front.state_RNIVIRQZ0Z_0 ));
    InMux I__9966 (
            .O(N__54823),
            .I(N__54819));
    InMux I__9965 (
            .O(N__54822),
            .I(N__54816));
    LocalMux I__9964 (
            .O(N__54819),
            .I(N__54807));
    LocalMux I__9963 (
            .O(N__54816),
            .I(N__54807));
    InMux I__9962 (
            .O(N__54815),
            .I(N__54802));
    InMux I__9961 (
            .O(N__54814),
            .I(N__54802));
    InMux I__9960 (
            .O(N__54813),
            .I(N__54799));
    InMux I__9959 (
            .O(N__54812),
            .I(N__54796));
    Span4Mux_h I__9958 (
            .O(N__54807),
            .I(N__54793));
    LocalMux I__9957 (
            .O(N__54802),
            .I(\uart_drone.stateZ0Z_4 ));
    LocalMux I__9956 (
            .O(N__54799),
            .I(\uart_drone.stateZ0Z_4 ));
    LocalMux I__9955 (
            .O(N__54796),
            .I(\uart_drone.stateZ0Z_4 ));
    Odrv4 I__9954 (
            .O(N__54793),
            .I(\uart_drone.stateZ0Z_4 ));
    InMux I__9953 (
            .O(N__54784),
            .I(N__54779));
    InMux I__9952 (
            .O(N__54783),
            .I(N__54776));
    InMux I__9951 (
            .O(N__54782),
            .I(N__54769));
    LocalMux I__9950 (
            .O(N__54779),
            .I(N__54764));
    LocalMux I__9949 (
            .O(N__54776),
            .I(N__54764));
    InMux I__9948 (
            .O(N__54775),
            .I(N__54757));
    InMux I__9947 (
            .O(N__54774),
            .I(N__54757));
    InMux I__9946 (
            .O(N__54773),
            .I(N__54757));
    InMux I__9945 (
            .O(N__54772),
            .I(N__54752));
    LocalMux I__9944 (
            .O(N__54769),
            .I(N__54749));
    Span4Mux_h I__9943 (
            .O(N__54764),
            .I(N__54744));
    LocalMux I__9942 (
            .O(N__54757),
            .I(N__54744));
    InMux I__9941 (
            .O(N__54756),
            .I(N__54739));
    InMux I__9940 (
            .O(N__54755),
            .I(N__54739));
    LocalMux I__9939 (
            .O(N__54752),
            .I(\uart_drone.timer_CountZ0Z_4 ));
    Odrv12 I__9938 (
            .O(N__54749),
            .I(\uart_drone.timer_CountZ0Z_4 ));
    Odrv4 I__9937 (
            .O(N__54744),
            .I(\uart_drone.timer_CountZ0Z_4 ));
    LocalMux I__9936 (
            .O(N__54739),
            .I(\uart_drone.timer_CountZ0Z_4 ));
    CascadeMux I__9935 (
            .O(N__54730),
            .I(\uart_drone.state_srsts_0_0_0_cascade_ ));
    InMux I__9934 (
            .O(N__54727),
            .I(N__54724));
    LocalMux I__9933 (
            .O(N__54724),
            .I(N__54720));
    InMux I__9932 (
            .O(N__54723),
            .I(N__54717));
    Span4Mux_v I__9931 (
            .O(N__54720),
            .I(N__54712));
    LocalMux I__9930 (
            .O(N__54717),
            .I(N__54712));
    Odrv4 I__9929 (
            .O(N__54712),
            .I(\uart_drone.N_126_li ));
    CascadeMux I__9928 (
            .O(N__54709),
            .I(N__54706));
    InMux I__9927 (
            .O(N__54706),
            .I(N__54703));
    LocalMux I__9926 (
            .O(N__54703),
            .I(N__54700));
    Span4Mux_v I__9925 (
            .O(N__54700),
            .I(N__54696));
    InMux I__9924 (
            .O(N__54699),
            .I(N__54693));
    Odrv4 I__9923 (
            .O(N__54696),
            .I(\uart_drone.stateZ0Z_0 ));
    LocalMux I__9922 (
            .O(N__54693),
            .I(\uart_drone.stateZ0Z_0 ));
    CascadeMux I__9921 (
            .O(N__54688),
            .I(N__54685));
    InMux I__9920 (
            .O(N__54685),
            .I(N__54682));
    LocalMux I__9919 (
            .O(N__54682),
            .I(N__54679));
    Odrv4 I__9918 (
            .O(N__54679),
            .I(\pid_side.error_i_acumm_13_0_a2_3_0_2 ));
    InMux I__9917 (
            .O(N__54676),
            .I(N__54673));
    LocalMux I__9916 (
            .O(N__54673),
            .I(N__54668));
    InMux I__9915 (
            .O(N__54672),
            .I(N__54665));
    CascadeMux I__9914 (
            .O(N__54671),
            .I(N__54662));
    Span4Mux_h I__9913 (
            .O(N__54668),
            .I(N__54657));
    LocalMux I__9912 (
            .O(N__54665),
            .I(N__54657));
    InMux I__9911 (
            .O(N__54662),
            .I(N__54654));
    Span4Mux_h I__9910 (
            .O(N__54657),
            .I(N__54651));
    LocalMux I__9909 (
            .O(N__54654),
            .I(front_order_10));
    Odrv4 I__9908 (
            .O(N__54651),
            .I(front_order_10));
    InMux I__9907 (
            .O(N__54646),
            .I(N__54643));
    LocalMux I__9906 (
            .O(N__54643),
            .I(N__54638));
    InMux I__9905 (
            .O(N__54642),
            .I(N__54635));
    CascadeMux I__9904 (
            .O(N__54641),
            .I(N__54632));
    Span4Mux_v I__9903 (
            .O(N__54638),
            .I(N__54629));
    LocalMux I__9902 (
            .O(N__54635),
            .I(N__54626));
    InMux I__9901 (
            .O(N__54632),
            .I(N__54623));
    Span4Mux_h I__9900 (
            .O(N__54629),
            .I(N__54618));
    Span4Mux_v I__9899 (
            .O(N__54626),
            .I(N__54618));
    LocalMux I__9898 (
            .O(N__54623),
            .I(front_order_11));
    Odrv4 I__9897 (
            .O(N__54618),
            .I(front_order_11));
    CascadeMux I__9896 (
            .O(N__54613),
            .I(N__54610));
    InMux I__9895 (
            .O(N__54610),
            .I(N__54607));
    LocalMux I__9894 (
            .O(N__54607),
            .I(N__54604));
    Span4Mux_s1_v I__9893 (
            .O(N__54604),
            .I(N__54599));
    InMux I__9892 (
            .O(N__54603),
            .I(N__54596));
    CascadeMux I__9891 (
            .O(N__54602),
            .I(N__54593));
    Span4Mux_v I__9890 (
            .O(N__54599),
            .I(N__54590));
    LocalMux I__9889 (
            .O(N__54596),
            .I(N__54587));
    InMux I__9888 (
            .O(N__54593),
            .I(N__54584));
    Span4Mux_h I__9887 (
            .O(N__54590),
            .I(N__54581));
    Span4Mux_h I__9886 (
            .O(N__54587),
            .I(N__54578));
    LocalMux I__9885 (
            .O(N__54584),
            .I(front_order_6));
    Odrv4 I__9884 (
            .O(N__54581),
            .I(front_order_6));
    Odrv4 I__9883 (
            .O(N__54578),
            .I(front_order_6));
    InMux I__9882 (
            .O(N__54571),
            .I(N__54566));
    InMux I__9881 (
            .O(N__54570),
            .I(N__54563));
    CascadeMux I__9880 (
            .O(N__54569),
            .I(N__54560));
    LocalMux I__9879 (
            .O(N__54566),
            .I(N__54555));
    LocalMux I__9878 (
            .O(N__54563),
            .I(N__54555));
    InMux I__9877 (
            .O(N__54560),
            .I(N__54552));
    Span4Mux_h I__9876 (
            .O(N__54555),
            .I(N__54549));
    LocalMux I__9875 (
            .O(N__54552),
            .I(front_order_7));
    Odrv4 I__9874 (
            .O(N__54549),
            .I(front_order_7));
    InMux I__9873 (
            .O(N__54544),
            .I(N__54540));
    InMux I__9872 (
            .O(N__54543),
            .I(N__54537));
    LocalMux I__9871 (
            .O(N__54540),
            .I(N__54533));
    LocalMux I__9870 (
            .O(N__54537),
            .I(N__54530));
    InMux I__9869 (
            .O(N__54536),
            .I(N__54527));
    Span12Mux_s9_v I__9868 (
            .O(N__54533),
            .I(N__54524));
    Span4Mux_h I__9867 (
            .O(N__54530),
            .I(N__54521));
    LocalMux I__9866 (
            .O(N__54527),
            .I(front_order_8));
    Odrv12 I__9865 (
            .O(N__54524),
            .I(front_order_8));
    Odrv4 I__9864 (
            .O(N__54521),
            .I(front_order_8));
    CascadeMux I__9863 (
            .O(N__54514),
            .I(N__54511));
    InMux I__9862 (
            .O(N__54511),
            .I(N__54506));
    InMux I__9861 (
            .O(N__54510),
            .I(N__54503));
    CascadeMux I__9860 (
            .O(N__54509),
            .I(N__54500));
    LocalMux I__9859 (
            .O(N__54506),
            .I(N__54495));
    LocalMux I__9858 (
            .O(N__54503),
            .I(N__54495));
    InMux I__9857 (
            .O(N__54500),
            .I(N__54492));
    Span4Mux_h I__9856 (
            .O(N__54495),
            .I(N__54489));
    LocalMux I__9855 (
            .O(N__54492),
            .I(front_order_9));
    Odrv4 I__9854 (
            .O(N__54489),
            .I(front_order_9));
    InMux I__9853 (
            .O(N__54484),
            .I(N__54480));
    InMux I__9852 (
            .O(N__54483),
            .I(N__54477));
    LocalMux I__9851 (
            .O(N__54480),
            .I(N__54474));
    LocalMux I__9850 (
            .O(N__54477),
            .I(N__54470));
    Span4Mux_v I__9849 (
            .O(N__54474),
            .I(N__54467));
    InMux I__9848 (
            .O(N__54473),
            .I(N__54464));
    Span4Mux_h I__9847 (
            .O(N__54470),
            .I(N__54461));
    Span4Mux_v I__9846 (
            .O(N__54467),
            .I(N__54458));
    LocalMux I__9845 (
            .O(N__54464),
            .I(side_order_11));
    Odrv4 I__9844 (
            .O(N__54461),
            .I(side_order_11));
    Odrv4 I__9843 (
            .O(N__54458),
            .I(side_order_11));
    CascadeMux I__9842 (
            .O(N__54451),
            .I(N__54448));
    InMux I__9841 (
            .O(N__54448),
            .I(N__54444));
    InMux I__9840 (
            .O(N__54447),
            .I(N__54441));
    LocalMux I__9839 (
            .O(N__54444),
            .I(N__54438));
    LocalMux I__9838 (
            .O(N__54441),
            .I(N__54434));
    Span4Mux_h I__9837 (
            .O(N__54438),
            .I(N__54431));
    InMux I__9836 (
            .O(N__54437),
            .I(N__54428));
    Span4Mux_h I__9835 (
            .O(N__54434),
            .I(N__54425));
    Span4Mux_v I__9834 (
            .O(N__54431),
            .I(N__54422));
    LocalMux I__9833 (
            .O(N__54428),
            .I(side_order_6));
    Odrv4 I__9832 (
            .O(N__54425),
            .I(side_order_6));
    Odrv4 I__9831 (
            .O(N__54422),
            .I(side_order_6));
    InMux I__9830 (
            .O(N__54415),
            .I(N__54411));
    InMux I__9829 (
            .O(N__54414),
            .I(N__54407));
    LocalMux I__9828 (
            .O(N__54411),
            .I(N__54404));
    InMux I__9827 (
            .O(N__54410),
            .I(N__54401));
    LocalMux I__9826 (
            .O(N__54407),
            .I(N__54398));
    Span4Mux_v I__9825 (
            .O(N__54404),
            .I(N__54395));
    LocalMux I__9824 (
            .O(N__54401),
            .I(N__54390));
    Span4Mux_v I__9823 (
            .O(N__54398),
            .I(N__54390));
    Odrv4 I__9822 (
            .O(N__54395),
            .I(side_order_7));
    Odrv4 I__9821 (
            .O(N__54390),
            .I(side_order_7));
    InMux I__9820 (
            .O(N__54385),
            .I(N__54381));
    InMux I__9819 (
            .O(N__54384),
            .I(N__54378));
    LocalMux I__9818 (
            .O(N__54381),
            .I(N__54375));
    LocalMux I__9817 (
            .O(N__54378),
            .I(N__54371));
    Span4Mux_v I__9816 (
            .O(N__54375),
            .I(N__54368));
    InMux I__9815 (
            .O(N__54374),
            .I(N__54365));
    Span4Mux_v I__9814 (
            .O(N__54371),
            .I(N__54362));
    Span4Mux_h I__9813 (
            .O(N__54368),
            .I(N__54359));
    LocalMux I__9812 (
            .O(N__54365),
            .I(N__54354));
    Span4Mux_v I__9811 (
            .O(N__54362),
            .I(N__54354));
    Odrv4 I__9810 (
            .O(N__54359),
            .I(side_order_8));
    Odrv4 I__9809 (
            .O(N__54354),
            .I(side_order_8));
    InMux I__9808 (
            .O(N__54349),
            .I(N__54345));
    InMux I__9807 (
            .O(N__54348),
            .I(N__54342));
    LocalMux I__9806 (
            .O(N__54345),
            .I(N__54338));
    LocalMux I__9805 (
            .O(N__54342),
            .I(N__54335));
    InMux I__9804 (
            .O(N__54341),
            .I(N__54332));
    Span4Mux_v I__9803 (
            .O(N__54338),
            .I(N__54329));
    Span12Mux_h I__9802 (
            .O(N__54335),
            .I(N__54326));
    LocalMux I__9801 (
            .O(N__54332),
            .I(side_order_9));
    Odrv4 I__9800 (
            .O(N__54329),
            .I(side_order_9));
    Odrv12 I__9799 (
            .O(N__54326),
            .I(side_order_9));
    CascadeMux I__9798 (
            .O(N__54319),
            .I(N__54316));
    InMux I__9797 (
            .O(N__54316),
            .I(N__54312));
    InMux I__9796 (
            .O(N__54315),
            .I(N__54308));
    LocalMux I__9795 (
            .O(N__54312),
            .I(N__54305));
    InMux I__9794 (
            .O(N__54311),
            .I(N__54302));
    LocalMux I__9793 (
            .O(N__54308),
            .I(N__54299));
    Span4Mux_h I__9792 (
            .O(N__54305),
            .I(N__54296));
    LocalMux I__9791 (
            .O(N__54302),
            .I(\ppm_encoder_1.throttleZ0Z_7 ));
    Odrv12 I__9790 (
            .O(N__54299),
            .I(\ppm_encoder_1.throttleZ0Z_7 ));
    Odrv4 I__9789 (
            .O(N__54296),
            .I(\ppm_encoder_1.throttleZ0Z_7 ));
    CascadeMux I__9788 (
            .O(N__54289),
            .I(N__54284));
    InMux I__9787 (
            .O(N__54288),
            .I(N__54281));
    InMux I__9786 (
            .O(N__54287),
            .I(N__54278));
    InMux I__9785 (
            .O(N__54284),
            .I(N__54275));
    LocalMux I__9784 (
            .O(N__54281),
            .I(N__54272));
    LocalMux I__9783 (
            .O(N__54278),
            .I(N__54269));
    LocalMux I__9782 (
            .O(N__54275),
            .I(\ppm_encoder_1.aileronZ0Z_7 ));
    Odrv12 I__9781 (
            .O(N__54272),
            .I(\ppm_encoder_1.aileronZ0Z_7 ));
    Odrv12 I__9780 (
            .O(N__54269),
            .I(\ppm_encoder_1.aileronZ0Z_7 ));
    CascadeMux I__9779 (
            .O(N__54262),
            .I(N__54256));
    CascadeMux I__9778 (
            .O(N__54261),
            .I(N__54252));
    InMux I__9777 (
            .O(N__54260),
            .I(N__54246));
    InMux I__9776 (
            .O(N__54259),
            .I(N__54242));
    InMux I__9775 (
            .O(N__54256),
            .I(N__54239));
    InMux I__9774 (
            .O(N__54255),
            .I(N__54235));
    InMux I__9773 (
            .O(N__54252),
            .I(N__54232));
    CascadeMux I__9772 (
            .O(N__54251),
            .I(N__54228));
    InMux I__9771 (
            .O(N__54250),
            .I(N__54222));
    InMux I__9770 (
            .O(N__54249),
            .I(N__54222));
    LocalMux I__9769 (
            .O(N__54246),
            .I(N__54219));
    InMux I__9768 (
            .O(N__54245),
            .I(N__54216));
    LocalMux I__9767 (
            .O(N__54242),
            .I(N__54213));
    LocalMux I__9766 (
            .O(N__54239),
            .I(N__54210));
    InMux I__9765 (
            .O(N__54238),
            .I(N__54207));
    LocalMux I__9764 (
            .O(N__54235),
            .I(N__54204));
    LocalMux I__9763 (
            .O(N__54232),
            .I(N__54201));
    InMux I__9762 (
            .O(N__54231),
            .I(N__54196));
    InMux I__9761 (
            .O(N__54228),
            .I(N__54196));
    CascadeMux I__9760 (
            .O(N__54227),
            .I(N__54190));
    LocalMux I__9759 (
            .O(N__54222),
            .I(N__54187));
    Span4Mux_h I__9758 (
            .O(N__54219),
            .I(N__54182));
    LocalMux I__9757 (
            .O(N__54216),
            .I(N__54182));
    Span4Mux_v I__9756 (
            .O(N__54213),
            .I(N__54179));
    Span4Mux_v I__9755 (
            .O(N__54210),
            .I(N__54176));
    LocalMux I__9754 (
            .O(N__54207),
            .I(N__54173));
    Span4Mux_h I__9753 (
            .O(N__54204),
            .I(N__54166));
    Span4Mux_v I__9752 (
            .O(N__54201),
            .I(N__54166));
    LocalMux I__9751 (
            .O(N__54196),
            .I(N__54166));
    InMux I__9750 (
            .O(N__54195),
            .I(N__54159));
    InMux I__9749 (
            .O(N__54194),
            .I(N__54156));
    InMux I__9748 (
            .O(N__54193),
            .I(N__54151));
    InMux I__9747 (
            .O(N__54190),
            .I(N__54151));
    Span4Mux_v I__9746 (
            .O(N__54187),
            .I(N__54144));
    Span4Mux_v I__9745 (
            .O(N__54182),
            .I(N__54144));
    Span4Mux_h I__9744 (
            .O(N__54179),
            .I(N__54144));
    Span4Mux_h I__9743 (
            .O(N__54176),
            .I(N__54137));
    Span4Mux_v I__9742 (
            .O(N__54173),
            .I(N__54137));
    Span4Mux_v I__9741 (
            .O(N__54166),
            .I(N__54137));
    InMux I__9740 (
            .O(N__54165),
            .I(N__54128));
    InMux I__9739 (
            .O(N__54164),
            .I(N__54128));
    InMux I__9738 (
            .O(N__54163),
            .I(N__54128));
    InMux I__9737 (
            .O(N__54162),
            .I(N__54128));
    LocalMux I__9736 (
            .O(N__54159),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    LocalMux I__9735 (
            .O(N__54156),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    LocalMux I__9734 (
            .O(N__54151),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    Odrv4 I__9733 (
            .O(N__54144),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    Odrv4 I__9732 (
            .O(N__54137),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    LocalMux I__9731 (
            .O(N__54128),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    InMux I__9730 (
            .O(N__54115),
            .I(N__54111));
    InMux I__9729 (
            .O(N__54114),
            .I(N__54103));
    LocalMux I__9728 (
            .O(N__54111),
            .I(N__54099));
    InMux I__9727 (
            .O(N__54110),
            .I(N__54096));
    InMux I__9726 (
            .O(N__54109),
            .I(N__54093));
    InMux I__9725 (
            .O(N__54108),
            .I(N__54090));
    InMux I__9724 (
            .O(N__54107),
            .I(N__54085));
    InMux I__9723 (
            .O(N__54106),
            .I(N__54085));
    LocalMux I__9722 (
            .O(N__54103),
            .I(N__54082));
    InMux I__9721 (
            .O(N__54102),
            .I(N__54079));
    Span4Mux_h I__9720 (
            .O(N__54099),
            .I(N__54071));
    LocalMux I__9719 (
            .O(N__54096),
            .I(N__54068));
    LocalMux I__9718 (
            .O(N__54093),
            .I(N__54065));
    LocalMux I__9717 (
            .O(N__54090),
            .I(N__54060));
    LocalMux I__9716 (
            .O(N__54085),
            .I(N__54060));
    Span4Mux_h I__9715 (
            .O(N__54082),
            .I(N__54057));
    LocalMux I__9714 (
            .O(N__54079),
            .I(N__54054));
    InMux I__9713 (
            .O(N__54078),
            .I(N__54051));
    InMux I__9712 (
            .O(N__54077),
            .I(N__54042));
    InMux I__9711 (
            .O(N__54076),
            .I(N__54042));
    InMux I__9710 (
            .O(N__54075),
            .I(N__54037));
    InMux I__9709 (
            .O(N__54074),
            .I(N__54037));
    Span4Mux_h I__9708 (
            .O(N__54071),
            .I(N__54034));
    Span4Mux_s3_v I__9707 (
            .O(N__54068),
            .I(N__54031));
    Span4Mux_h I__9706 (
            .O(N__54065),
            .I(N__54026));
    Span4Mux_h I__9705 (
            .O(N__54060),
            .I(N__54026));
    Span4Mux_h I__9704 (
            .O(N__54057),
            .I(N__54019));
    Span4Mux_h I__9703 (
            .O(N__54054),
            .I(N__54019));
    LocalMux I__9702 (
            .O(N__54051),
            .I(N__54019));
    InMux I__9701 (
            .O(N__54050),
            .I(N__54010));
    InMux I__9700 (
            .O(N__54049),
            .I(N__54010));
    InMux I__9699 (
            .O(N__54048),
            .I(N__54010));
    InMux I__9698 (
            .O(N__54047),
            .I(N__54010));
    LocalMux I__9697 (
            .O(N__54042),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    LocalMux I__9696 (
            .O(N__54037),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    Odrv4 I__9695 (
            .O(N__54034),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    Odrv4 I__9694 (
            .O(N__54031),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    Odrv4 I__9693 (
            .O(N__54026),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    Odrv4 I__9692 (
            .O(N__54019),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    LocalMux I__9691 (
            .O(N__54010),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    InMux I__9690 (
            .O(N__53995),
            .I(N__53992));
    LocalMux I__9689 (
            .O(N__53992),
            .I(N__53989));
    Odrv4 I__9688 (
            .O(N__53989),
            .I(\ppm_encoder_1.pulses2count_9_i_0_7 ));
    InMux I__9687 (
            .O(N__53986),
            .I(N__53980));
    InMux I__9686 (
            .O(N__53985),
            .I(N__53976));
    CascadeMux I__9685 (
            .O(N__53984),
            .I(N__53970));
    CascadeMux I__9684 (
            .O(N__53983),
            .I(N__53967));
    LocalMux I__9683 (
            .O(N__53980),
            .I(N__53964));
    InMux I__9682 (
            .O(N__53979),
            .I(N__53961));
    LocalMux I__9681 (
            .O(N__53976),
            .I(N__53958));
    InMux I__9680 (
            .O(N__53975),
            .I(N__53955));
    InMux I__9679 (
            .O(N__53974),
            .I(N__53952));
    InMux I__9678 (
            .O(N__53973),
            .I(N__53945));
    InMux I__9677 (
            .O(N__53970),
            .I(N__53945));
    InMux I__9676 (
            .O(N__53967),
            .I(N__53945));
    Odrv4 I__9675 (
            .O(N__53964),
            .I(\uart_drone.stateZ0Z_3 ));
    LocalMux I__9674 (
            .O(N__53961),
            .I(\uart_drone.stateZ0Z_3 ));
    Odrv4 I__9673 (
            .O(N__53958),
            .I(\uart_drone.stateZ0Z_3 ));
    LocalMux I__9672 (
            .O(N__53955),
            .I(\uart_drone.stateZ0Z_3 ));
    LocalMux I__9671 (
            .O(N__53952),
            .I(\uart_drone.stateZ0Z_3 ));
    LocalMux I__9670 (
            .O(N__53945),
            .I(\uart_drone.stateZ0Z_3 ));
    InMux I__9669 (
            .O(N__53932),
            .I(N__53928));
    InMux I__9668 (
            .O(N__53931),
            .I(N__53925));
    LocalMux I__9667 (
            .O(N__53928),
            .I(N__53922));
    LocalMux I__9666 (
            .O(N__53925),
            .I(N__53917));
    Span4Mux_h I__9665 (
            .O(N__53922),
            .I(N__53917));
    Span4Mux_v I__9664 (
            .O(N__53917),
            .I(N__53914));
    Odrv4 I__9663 (
            .O(N__53914),
            .I(side_order_13));
    InMux I__9662 (
            .O(N__53911),
            .I(N__53908));
    LocalMux I__9661 (
            .O(N__53908),
            .I(N__53904));
    InMux I__9660 (
            .O(N__53907),
            .I(N__53901));
    Span4Mux_h I__9659 (
            .O(N__53904),
            .I(N__53896));
    LocalMux I__9658 (
            .O(N__53901),
            .I(N__53896));
    Span4Mux_v I__9657 (
            .O(N__53896),
            .I(N__53893));
    Odrv4 I__9656 (
            .O(N__53893),
            .I(\ppm_encoder_1.aileronZ0Z_14 ));
    CascadeMux I__9655 (
            .O(N__53890),
            .I(N__53887));
    InMux I__9654 (
            .O(N__53887),
            .I(N__53883));
    CascadeMux I__9653 (
            .O(N__53886),
            .I(N__53880));
    LocalMux I__9652 (
            .O(N__53883),
            .I(N__53877));
    InMux I__9651 (
            .O(N__53880),
            .I(N__53874));
    Span4Mux_v I__9650 (
            .O(N__53877),
            .I(N__53871));
    LocalMux I__9649 (
            .O(N__53874),
            .I(N__53868));
    Span4Mux_h I__9648 (
            .O(N__53871),
            .I(N__53865));
    Span4Mux_h I__9647 (
            .O(N__53868),
            .I(N__53862));
    Span4Mux_h I__9646 (
            .O(N__53865),
            .I(N__53859));
    Span4Mux_v I__9645 (
            .O(N__53862),
            .I(N__53856));
    Odrv4 I__9644 (
            .O(N__53859),
            .I(\ppm_encoder_1.throttleZ0Z_14 ));
    Odrv4 I__9643 (
            .O(N__53856),
            .I(\ppm_encoder_1.throttleZ0Z_14 ));
    CascadeMux I__9642 (
            .O(N__53851),
            .I(\ppm_encoder_1.pulses2count_9_i_0_14_cascade_ ));
    CascadeMux I__9641 (
            .O(N__53848),
            .I(N__53845));
    InMux I__9640 (
            .O(N__53845),
            .I(N__53842));
    LocalMux I__9639 (
            .O(N__53842),
            .I(N__53839));
    Span4Mux_s1_v I__9638 (
            .O(N__53839),
            .I(N__53836));
    Odrv4 I__9637 (
            .O(N__53836),
            .I(\ppm_encoder_1.pulses2count_9_i_1_14 ));
    InMux I__9636 (
            .O(N__53833),
            .I(N__53830));
    LocalMux I__9635 (
            .O(N__53830),
            .I(N__53827));
    Span4Mux_h I__9634 (
            .O(N__53827),
            .I(N__53824));
    Span4Mux_h I__9633 (
            .O(N__53824),
            .I(N__53821));
    Odrv4 I__9632 (
            .O(N__53821),
            .I(\ppm_encoder_1.un2_throttle_0_0_2_5 ));
    CascadeMux I__9631 (
            .O(N__53818),
            .I(N__53815));
    InMux I__9630 (
            .O(N__53815),
            .I(N__53812));
    LocalMux I__9629 (
            .O(N__53812),
            .I(\ppm_encoder_1.pulses2count_9_i_0_5 ));
    InMux I__9628 (
            .O(N__53809),
            .I(N__53802));
    InMux I__9627 (
            .O(N__53808),
            .I(N__53799));
    CascadeMux I__9626 (
            .O(N__53807),
            .I(N__53790));
    InMux I__9625 (
            .O(N__53806),
            .I(N__53782));
    InMux I__9624 (
            .O(N__53805),
            .I(N__53782));
    LocalMux I__9623 (
            .O(N__53802),
            .I(N__53776));
    LocalMux I__9622 (
            .O(N__53799),
            .I(N__53773));
    InMux I__9621 (
            .O(N__53798),
            .I(N__53768));
    InMux I__9620 (
            .O(N__53797),
            .I(N__53761));
    InMux I__9619 (
            .O(N__53796),
            .I(N__53761));
    InMux I__9618 (
            .O(N__53795),
            .I(N__53761));
    InMux I__9617 (
            .O(N__53794),
            .I(N__53754));
    InMux I__9616 (
            .O(N__53793),
            .I(N__53754));
    InMux I__9615 (
            .O(N__53790),
            .I(N__53754));
    InMux I__9614 (
            .O(N__53789),
            .I(N__53747));
    InMux I__9613 (
            .O(N__53788),
            .I(N__53747));
    InMux I__9612 (
            .O(N__53787),
            .I(N__53747));
    LocalMux I__9611 (
            .O(N__53782),
            .I(N__53744));
    InMux I__9610 (
            .O(N__53781),
            .I(N__53741));
    InMux I__9609 (
            .O(N__53780),
            .I(N__53736));
    InMux I__9608 (
            .O(N__53779),
            .I(N__53736));
    Span4Mux_v I__9607 (
            .O(N__53776),
            .I(N__53731));
    Span4Mux_v I__9606 (
            .O(N__53773),
            .I(N__53731));
    InMux I__9605 (
            .O(N__53772),
            .I(N__53726));
    InMux I__9604 (
            .O(N__53771),
            .I(N__53726));
    LocalMux I__9603 (
            .O(N__53768),
            .I(N__53721));
    LocalMux I__9602 (
            .O(N__53761),
            .I(N__53721));
    LocalMux I__9601 (
            .O(N__53754),
            .I(N__53716));
    LocalMux I__9600 (
            .O(N__53747),
            .I(N__53716));
    Span4Mux_s2_v I__9599 (
            .O(N__53744),
            .I(N__53709));
    LocalMux I__9598 (
            .O(N__53741),
            .I(N__53709));
    LocalMux I__9597 (
            .O(N__53736),
            .I(N__53709));
    Odrv4 I__9596 (
            .O(N__53731),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z2 ));
    LocalMux I__9595 (
            .O(N__53726),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z2 ));
    Odrv12 I__9594 (
            .O(N__53721),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z2 ));
    Odrv4 I__9593 (
            .O(N__53716),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z2 ));
    Odrv4 I__9592 (
            .O(N__53709),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z2 ));
    InMux I__9591 (
            .O(N__53698),
            .I(N__53687));
    CascadeMux I__9590 (
            .O(N__53697),
            .I(N__53683));
    InMux I__9589 (
            .O(N__53696),
            .I(N__53676));
    InMux I__9588 (
            .O(N__53695),
            .I(N__53673));
    InMux I__9587 (
            .O(N__53694),
            .I(N__53666));
    InMux I__9586 (
            .O(N__53693),
            .I(N__53666));
    InMux I__9585 (
            .O(N__53692),
            .I(N__53666));
    InMux I__9584 (
            .O(N__53691),
            .I(N__53661));
    InMux I__9583 (
            .O(N__53690),
            .I(N__53661));
    LocalMux I__9582 (
            .O(N__53687),
            .I(N__53657));
    InMux I__9581 (
            .O(N__53686),
            .I(N__53653));
    InMux I__9580 (
            .O(N__53683),
            .I(N__53648));
    InMux I__9579 (
            .O(N__53682),
            .I(N__53648));
    CascadeMux I__9578 (
            .O(N__53681),
            .I(N__53645));
    CascadeMux I__9577 (
            .O(N__53680),
            .I(N__53640));
    InMux I__9576 (
            .O(N__53679),
            .I(N__53635));
    LocalMux I__9575 (
            .O(N__53676),
            .I(N__53630));
    LocalMux I__9574 (
            .O(N__53673),
            .I(N__53630));
    LocalMux I__9573 (
            .O(N__53666),
            .I(N__53627));
    LocalMux I__9572 (
            .O(N__53661),
            .I(N__53622));
    InMux I__9571 (
            .O(N__53660),
            .I(N__53619));
    Span4Mux_h I__9570 (
            .O(N__53657),
            .I(N__53616));
    InMux I__9569 (
            .O(N__53656),
            .I(N__53613));
    LocalMux I__9568 (
            .O(N__53653),
            .I(N__53610));
    LocalMux I__9567 (
            .O(N__53648),
            .I(N__53607));
    InMux I__9566 (
            .O(N__53645),
            .I(N__53600));
    InMux I__9565 (
            .O(N__53644),
            .I(N__53600));
    InMux I__9564 (
            .O(N__53643),
            .I(N__53600));
    InMux I__9563 (
            .O(N__53640),
            .I(N__53593));
    InMux I__9562 (
            .O(N__53639),
            .I(N__53593));
    InMux I__9561 (
            .O(N__53638),
            .I(N__53593));
    LocalMux I__9560 (
            .O(N__53635),
            .I(N__53586));
    Span4Mux_h I__9559 (
            .O(N__53630),
            .I(N__53586));
    Span4Mux_s1_v I__9558 (
            .O(N__53627),
            .I(N__53586));
    InMux I__9557 (
            .O(N__53626),
            .I(N__53581));
    InMux I__9556 (
            .O(N__53625),
            .I(N__53581));
    Span4Mux_s2_v I__9555 (
            .O(N__53622),
            .I(N__53576));
    LocalMux I__9554 (
            .O(N__53619),
            .I(N__53576));
    Odrv4 I__9553 (
            .O(N__53616),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z2 ));
    LocalMux I__9552 (
            .O(N__53613),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z2 ));
    Odrv4 I__9551 (
            .O(N__53610),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z2 ));
    Odrv12 I__9550 (
            .O(N__53607),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z2 ));
    LocalMux I__9549 (
            .O(N__53600),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z2 ));
    LocalMux I__9548 (
            .O(N__53593),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z2 ));
    Odrv4 I__9547 (
            .O(N__53586),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z2 ));
    LocalMux I__9546 (
            .O(N__53581),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z2 ));
    Odrv4 I__9545 (
            .O(N__53576),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z2 ));
    CascadeMux I__9544 (
            .O(N__53557),
            .I(\ppm_encoder_1.N_301_cascade_ ));
    InMux I__9543 (
            .O(N__53554),
            .I(N__53551));
    LocalMux I__9542 (
            .O(N__53551),
            .I(N__53547));
    InMux I__9541 (
            .O(N__53550),
            .I(N__53544));
    Span4Mux_v I__9540 (
            .O(N__53547),
            .I(N__53541));
    LocalMux I__9539 (
            .O(N__53544),
            .I(N__53538));
    Odrv4 I__9538 (
            .O(N__53541),
            .I(\ppm_encoder_1.un2_throttle_0_2_6 ));
    Odrv12 I__9537 (
            .O(N__53538),
            .I(\ppm_encoder_1.un2_throttle_0_2_6 ));
    InMux I__9536 (
            .O(N__53533),
            .I(N__53530));
    LocalMux I__9535 (
            .O(N__53530),
            .I(N__53527));
    Span4Mux_s2_v I__9534 (
            .O(N__53527),
            .I(N__53524));
    Odrv4 I__9533 (
            .O(N__53524),
            .I(\ppm_encoder_1.pulses2count_9_0_0_6 ));
    InMux I__9532 (
            .O(N__53521),
            .I(N__53508));
    InMux I__9531 (
            .O(N__53520),
            .I(N__53508));
    InMux I__9530 (
            .O(N__53519),
            .I(N__53508));
    InMux I__9529 (
            .O(N__53518),
            .I(N__53508));
    InMux I__9528 (
            .O(N__53517),
            .I(N__53504));
    LocalMux I__9527 (
            .O(N__53508),
            .I(N__53498));
    InMux I__9526 (
            .O(N__53507),
            .I(N__53495));
    LocalMux I__9525 (
            .O(N__53504),
            .I(N__53492));
    InMux I__9524 (
            .O(N__53503),
            .I(N__53485));
    InMux I__9523 (
            .O(N__53502),
            .I(N__53485));
    InMux I__9522 (
            .O(N__53501),
            .I(N__53485));
    Span4Mux_v I__9521 (
            .O(N__53498),
            .I(N__53482));
    LocalMux I__9520 (
            .O(N__53495),
            .I(\ppm_encoder_1.N_301 ));
    Odrv4 I__9519 (
            .O(N__53492),
            .I(\ppm_encoder_1.N_301 ));
    LocalMux I__9518 (
            .O(N__53485),
            .I(\ppm_encoder_1.N_301 ));
    Odrv4 I__9517 (
            .O(N__53482),
            .I(\ppm_encoder_1.N_301 ));
    CascadeMux I__9516 (
            .O(N__53473),
            .I(N__53470));
    InMux I__9515 (
            .O(N__53470),
            .I(N__53467));
    LocalMux I__9514 (
            .O(N__53467),
            .I(N__53464));
    Span4Mux_s1_v I__9513 (
            .O(N__53464),
            .I(N__53461));
    Odrv4 I__9512 (
            .O(N__53461),
            .I(\ppm_encoder_1.pulses2count_9_i_1_7 ));
    InMux I__9511 (
            .O(N__53458),
            .I(N__53455));
    LocalMux I__9510 (
            .O(N__53455),
            .I(N__53451));
    InMux I__9509 (
            .O(N__53454),
            .I(N__53448));
    Span4Mux_h I__9508 (
            .O(N__53451),
            .I(N__53445));
    LocalMux I__9507 (
            .O(N__53448),
            .I(N__53442));
    Span4Mux_h I__9506 (
            .O(N__53445),
            .I(N__53436));
    Span4Mux_h I__9505 (
            .O(N__53442),
            .I(N__53436));
    InMux I__9504 (
            .O(N__53441),
            .I(N__53433));
    Span4Mux_v I__9503 (
            .O(N__53436),
            .I(N__53430));
    LocalMux I__9502 (
            .O(N__53433),
            .I(side_order_10));
    Odrv4 I__9501 (
            .O(N__53430),
            .I(side_order_10));
    CascadeMux I__9500 (
            .O(N__53425),
            .I(N__53422));
    InMux I__9499 (
            .O(N__53422),
            .I(N__53418));
    InMux I__9498 (
            .O(N__53421),
            .I(N__53414));
    LocalMux I__9497 (
            .O(N__53418),
            .I(N__53411));
    InMux I__9496 (
            .O(N__53417),
            .I(N__53408));
    LocalMux I__9495 (
            .O(N__53414),
            .I(\ppm_encoder_1.counterZ0Z_11 ));
    Odrv4 I__9494 (
            .O(N__53411),
            .I(\ppm_encoder_1.counterZ0Z_11 ));
    LocalMux I__9493 (
            .O(N__53408),
            .I(\ppm_encoder_1.counterZ0Z_11 ));
    InMux I__9492 (
            .O(N__53401),
            .I(\ppm_encoder_1.un1_counter_13_cry_10 ));
    CascadeMux I__9491 (
            .O(N__53398),
            .I(N__53394));
    InMux I__9490 (
            .O(N__53397),
            .I(N__53391));
    InMux I__9489 (
            .O(N__53394),
            .I(N__53387));
    LocalMux I__9488 (
            .O(N__53391),
            .I(N__53384));
    InMux I__9487 (
            .O(N__53390),
            .I(N__53381));
    LocalMux I__9486 (
            .O(N__53387),
            .I(N__53378));
    Span4Mux_s2_v I__9485 (
            .O(N__53384),
            .I(N__53375));
    LocalMux I__9484 (
            .O(N__53381),
            .I(\ppm_encoder_1.counterZ0Z_12 ));
    Odrv12 I__9483 (
            .O(N__53378),
            .I(\ppm_encoder_1.counterZ0Z_12 ));
    Odrv4 I__9482 (
            .O(N__53375),
            .I(\ppm_encoder_1.counterZ0Z_12 ));
    InMux I__9481 (
            .O(N__53368),
            .I(\ppm_encoder_1.un1_counter_13_cry_11 ));
    InMux I__9480 (
            .O(N__53365),
            .I(N__53361));
    InMux I__9479 (
            .O(N__53364),
            .I(N__53357));
    LocalMux I__9478 (
            .O(N__53361),
            .I(N__53354));
    InMux I__9477 (
            .O(N__53360),
            .I(N__53351));
    LocalMux I__9476 (
            .O(N__53357),
            .I(N__53348));
    Span4Mux_s2_v I__9475 (
            .O(N__53354),
            .I(N__53345));
    LocalMux I__9474 (
            .O(N__53351),
            .I(\ppm_encoder_1.counterZ0Z_13 ));
    Odrv4 I__9473 (
            .O(N__53348),
            .I(\ppm_encoder_1.counterZ0Z_13 ));
    Odrv4 I__9472 (
            .O(N__53345),
            .I(\ppm_encoder_1.counterZ0Z_13 ));
    InMux I__9471 (
            .O(N__53338),
            .I(\ppm_encoder_1.un1_counter_13_cry_12 ));
    InMux I__9470 (
            .O(N__53335),
            .I(N__53328));
    InMux I__9469 (
            .O(N__53334),
            .I(N__53328));
    InMux I__9468 (
            .O(N__53333),
            .I(N__53325));
    LocalMux I__9467 (
            .O(N__53328),
            .I(N__53322));
    LocalMux I__9466 (
            .O(N__53325),
            .I(\ppm_encoder_1.counterZ0Z_14 ));
    Odrv4 I__9465 (
            .O(N__53322),
            .I(\ppm_encoder_1.counterZ0Z_14 ));
    InMux I__9464 (
            .O(N__53317),
            .I(\ppm_encoder_1.un1_counter_13_cry_13 ));
    InMux I__9463 (
            .O(N__53314),
            .I(N__53307));
    InMux I__9462 (
            .O(N__53313),
            .I(N__53307));
    InMux I__9461 (
            .O(N__53312),
            .I(N__53304));
    LocalMux I__9460 (
            .O(N__53307),
            .I(N__53301));
    LocalMux I__9459 (
            .O(N__53304),
            .I(\ppm_encoder_1.counterZ0Z_15 ));
    Odrv4 I__9458 (
            .O(N__53301),
            .I(\ppm_encoder_1.counterZ0Z_15 ));
    InMux I__9457 (
            .O(N__53296),
            .I(\ppm_encoder_1.un1_counter_13_cry_14 ));
    InMux I__9456 (
            .O(N__53293),
            .I(N__53289));
    InMux I__9455 (
            .O(N__53292),
            .I(N__53286));
    LocalMux I__9454 (
            .O(N__53289),
            .I(N__53282));
    LocalMux I__9453 (
            .O(N__53286),
            .I(N__53279));
    InMux I__9452 (
            .O(N__53285),
            .I(N__53276));
    Span4Mux_s1_v I__9451 (
            .O(N__53282),
            .I(N__53271));
    Span4Mux_h I__9450 (
            .O(N__53279),
            .I(N__53271));
    LocalMux I__9449 (
            .O(N__53276),
            .I(\ppm_encoder_1.counterZ0Z_16 ));
    Odrv4 I__9448 (
            .O(N__53271),
            .I(\ppm_encoder_1.counterZ0Z_16 ));
    InMux I__9447 (
            .O(N__53266),
            .I(bfn_12_4_0_));
    CascadeMux I__9446 (
            .O(N__53263),
            .I(N__53259));
    InMux I__9445 (
            .O(N__53262),
            .I(N__53256));
    InMux I__9444 (
            .O(N__53259),
            .I(N__53252));
    LocalMux I__9443 (
            .O(N__53256),
            .I(N__53249));
    InMux I__9442 (
            .O(N__53255),
            .I(N__53246));
    LocalMux I__9441 (
            .O(N__53252),
            .I(N__53243));
    Span4Mux_h I__9440 (
            .O(N__53249),
            .I(N__53240));
    LocalMux I__9439 (
            .O(N__53246),
            .I(\ppm_encoder_1.counterZ0Z_17 ));
    Odrv4 I__9438 (
            .O(N__53243),
            .I(\ppm_encoder_1.counterZ0Z_17 ));
    Odrv4 I__9437 (
            .O(N__53240),
            .I(\ppm_encoder_1.counterZ0Z_17 ));
    InMux I__9436 (
            .O(N__53233),
            .I(\ppm_encoder_1.un1_counter_13_cry_16 ));
    InMux I__9435 (
            .O(N__53230),
            .I(\ppm_encoder_1.un1_counter_13_cry_17 ));
    InMux I__9434 (
            .O(N__53227),
            .I(N__53221));
    InMux I__9433 (
            .O(N__53226),
            .I(N__53218));
    InMux I__9432 (
            .O(N__53225),
            .I(N__53213));
    InMux I__9431 (
            .O(N__53224),
            .I(N__53213));
    LocalMux I__9430 (
            .O(N__53221),
            .I(N__53210));
    LocalMux I__9429 (
            .O(N__53218),
            .I(\ppm_encoder_1.counterZ0Z_18 ));
    LocalMux I__9428 (
            .O(N__53213),
            .I(\ppm_encoder_1.counterZ0Z_18 ));
    Odrv4 I__9427 (
            .O(N__53210),
            .I(\ppm_encoder_1.counterZ0Z_18 ));
    SRMux I__9426 (
            .O(N__53203),
            .I(N__53198));
    SRMux I__9425 (
            .O(N__53202),
            .I(N__53195));
    SRMux I__9424 (
            .O(N__53201),
            .I(N__53192));
    LocalMux I__9423 (
            .O(N__53198),
            .I(\ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83 ));
    LocalMux I__9422 (
            .O(N__53195),
            .I(\ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83 ));
    LocalMux I__9421 (
            .O(N__53192),
            .I(\ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83 ));
    InMux I__9420 (
            .O(N__53185),
            .I(N__53181));
    InMux I__9419 (
            .O(N__53184),
            .I(N__53178));
    LocalMux I__9418 (
            .O(N__53181),
            .I(N__53175));
    LocalMux I__9417 (
            .O(N__53178),
            .I(N__53172));
    Span4Mux_v I__9416 (
            .O(N__53175),
            .I(N__53169));
    Span4Mux_h I__9415 (
            .O(N__53172),
            .I(N__53166));
    Span4Mux_v I__9414 (
            .O(N__53169),
            .I(N__53163));
    Odrv4 I__9413 (
            .O(N__53166),
            .I(side_order_12));
    Odrv4 I__9412 (
            .O(N__53163),
            .I(side_order_12));
    InMux I__9411 (
            .O(N__53158),
            .I(N__53155));
    LocalMux I__9410 (
            .O(N__53155),
            .I(N__53150));
    InMux I__9409 (
            .O(N__53154),
            .I(N__53147));
    InMux I__9408 (
            .O(N__53153),
            .I(N__53144));
    Span4Mux_v I__9407 (
            .O(N__53150),
            .I(N__53141));
    LocalMux I__9406 (
            .O(N__53147),
            .I(\ppm_encoder_1.counterZ0Z_3 ));
    LocalMux I__9405 (
            .O(N__53144),
            .I(\ppm_encoder_1.counterZ0Z_3 ));
    Odrv4 I__9404 (
            .O(N__53141),
            .I(\ppm_encoder_1.counterZ0Z_3 ));
    InMux I__9403 (
            .O(N__53134),
            .I(\ppm_encoder_1.un1_counter_13_cry_2 ));
    InMux I__9402 (
            .O(N__53131),
            .I(N__53126));
    InMux I__9401 (
            .O(N__53130),
            .I(N__53123));
    InMux I__9400 (
            .O(N__53129),
            .I(N__53120));
    LocalMux I__9399 (
            .O(N__53126),
            .I(\ppm_encoder_1.counterZ0Z_4 ));
    LocalMux I__9398 (
            .O(N__53123),
            .I(\ppm_encoder_1.counterZ0Z_4 ));
    LocalMux I__9397 (
            .O(N__53120),
            .I(\ppm_encoder_1.counterZ0Z_4 ));
    InMux I__9396 (
            .O(N__53113),
            .I(\ppm_encoder_1.un1_counter_13_cry_3 ));
    InMux I__9395 (
            .O(N__53110),
            .I(N__53105));
    InMux I__9394 (
            .O(N__53109),
            .I(N__53102));
    InMux I__9393 (
            .O(N__53108),
            .I(N__53099));
    LocalMux I__9392 (
            .O(N__53105),
            .I(\ppm_encoder_1.counterZ0Z_5 ));
    LocalMux I__9391 (
            .O(N__53102),
            .I(\ppm_encoder_1.counterZ0Z_5 ));
    LocalMux I__9390 (
            .O(N__53099),
            .I(\ppm_encoder_1.counterZ0Z_5 ));
    InMux I__9389 (
            .O(N__53092),
            .I(\ppm_encoder_1.un1_counter_13_cry_4 ));
    InMux I__9388 (
            .O(N__53089),
            .I(N__53084));
    InMux I__9387 (
            .O(N__53088),
            .I(N__53081));
    InMux I__9386 (
            .O(N__53087),
            .I(N__53078));
    LocalMux I__9385 (
            .O(N__53084),
            .I(\ppm_encoder_1.counterZ0Z_6 ));
    LocalMux I__9384 (
            .O(N__53081),
            .I(\ppm_encoder_1.counterZ0Z_6 ));
    LocalMux I__9383 (
            .O(N__53078),
            .I(\ppm_encoder_1.counterZ0Z_6 ));
    InMux I__9382 (
            .O(N__53071),
            .I(\ppm_encoder_1.un1_counter_13_cry_5 ));
    CascadeMux I__9381 (
            .O(N__53068),
            .I(N__53063));
    InMux I__9380 (
            .O(N__53067),
            .I(N__53060));
    InMux I__9379 (
            .O(N__53066),
            .I(N__53057));
    InMux I__9378 (
            .O(N__53063),
            .I(N__53054));
    LocalMux I__9377 (
            .O(N__53060),
            .I(N__53051));
    LocalMux I__9376 (
            .O(N__53057),
            .I(\ppm_encoder_1.counterZ0Z_7 ));
    LocalMux I__9375 (
            .O(N__53054),
            .I(\ppm_encoder_1.counterZ0Z_7 ));
    Odrv4 I__9374 (
            .O(N__53051),
            .I(\ppm_encoder_1.counterZ0Z_7 ));
    InMux I__9373 (
            .O(N__53044),
            .I(\ppm_encoder_1.un1_counter_13_cry_6 ));
    InMux I__9372 (
            .O(N__53041),
            .I(N__53037));
    InMux I__9371 (
            .O(N__53040),
            .I(N__53033));
    LocalMux I__9370 (
            .O(N__53037),
            .I(N__53030));
    InMux I__9369 (
            .O(N__53036),
            .I(N__53027));
    LocalMux I__9368 (
            .O(N__53033),
            .I(\ppm_encoder_1.counterZ0Z_8 ));
    Odrv4 I__9367 (
            .O(N__53030),
            .I(\ppm_encoder_1.counterZ0Z_8 ));
    LocalMux I__9366 (
            .O(N__53027),
            .I(\ppm_encoder_1.counterZ0Z_8 ));
    InMux I__9365 (
            .O(N__53020),
            .I(bfn_12_3_0_));
    InMux I__9364 (
            .O(N__53017),
            .I(N__53013));
    InMux I__9363 (
            .O(N__53016),
            .I(N__53009));
    LocalMux I__9362 (
            .O(N__53013),
            .I(N__53006));
    InMux I__9361 (
            .O(N__53012),
            .I(N__53003));
    LocalMux I__9360 (
            .O(N__53009),
            .I(\ppm_encoder_1.counterZ0Z_9 ));
    Odrv4 I__9359 (
            .O(N__53006),
            .I(\ppm_encoder_1.counterZ0Z_9 ));
    LocalMux I__9358 (
            .O(N__53003),
            .I(\ppm_encoder_1.counterZ0Z_9 ));
    InMux I__9357 (
            .O(N__52996),
            .I(\ppm_encoder_1.un1_counter_13_cry_8 ));
    InMux I__9356 (
            .O(N__52993),
            .I(N__52989));
    InMux I__9355 (
            .O(N__52992),
            .I(N__52985));
    LocalMux I__9354 (
            .O(N__52989),
            .I(N__52982));
    InMux I__9353 (
            .O(N__52988),
            .I(N__52979));
    LocalMux I__9352 (
            .O(N__52985),
            .I(\ppm_encoder_1.counterZ0Z_10 ));
    Odrv4 I__9351 (
            .O(N__52982),
            .I(\ppm_encoder_1.counterZ0Z_10 ));
    LocalMux I__9350 (
            .O(N__52979),
            .I(\ppm_encoder_1.counterZ0Z_10 ));
    InMux I__9349 (
            .O(N__52972),
            .I(\ppm_encoder_1.un1_counter_13_cry_9 ));
    InMux I__9348 (
            .O(N__52969),
            .I(N__52966));
    LocalMux I__9347 (
            .O(N__52966),
            .I(\ppm_encoder_1.pulses2countZ0Z_14 ));
    CascadeMux I__9346 (
            .O(N__52963),
            .I(N__52960));
    InMux I__9345 (
            .O(N__52960),
            .I(N__52957));
    LocalMux I__9344 (
            .O(N__52957),
            .I(N__52954));
    Odrv4 I__9343 (
            .O(N__52954),
            .I(\ppm_encoder_1.pulses2countZ0Z_15 ));
    InMux I__9342 (
            .O(N__52951),
            .I(N__52948));
    LocalMux I__9341 (
            .O(N__52948),
            .I(N__52945));
    Odrv4 I__9340 (
            .O(N__52945),
            .I(\ppm_encoder_1.counter24_0_I_45_c_RNOZ0 ));
    CascadeMux I__9339 (
            .O(N__52942),
            .I(\ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_a2_18_8_cascade_ ));
    InMux I__9338 (
            .O(N__52939),
            .I(N__52933));
    InMux I__9337 (
            .O(N__52938),
            .I(N__52933));
    LocalMux I__9336 (
            .O(N__52933),
            .I(N__52930));
    Span4Mux_v I__9335 (
            .O(N__52930),
            .I(N__52927));
    Odrv4 I__9334 (
            .O(N__52927),
            .I(\ppm_encoder_1.N_486_18 ));
    InMux I__9333 (
            .O(N__52924),
            .I(N__52921));
    LocalMux I__9332 (
            .O(N__52921),
            .I(\ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_a2_18_10 ));
    InMux I__9331 (
            .O(N__52918),
            .I(N__52915));
    LocalMux I__9330 (
            .O(N__52915),
            .I(\ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_a2_18_11 ));
    InMux I__9329 (
            .O(N__52912),
            .I(N__52909));
    LocalMux I__9328 (
            .O(N__52909),
            .I(\ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_a2_18_9 ));
    CascadeMux I__9327 (
            .O(N__52906),
            .I(N__52902));
    CascadeMux I__9326 (
            .O(N__52905),
            .I(N__52896));
    InMux I__9325 (
            .O(N__52902),
            .I(N__52874));
    InMux I__9324 (
            .O(N__52901),
            .I(N__52869));
    InMux I__9323 (
            .O(N__52900),
            .I(N__52869));
    InMux I__9322 (
            .O(N__52899),
            .I(N__52856));
    InMux I__9321 (
            .O(N__52896),
            .I(N__52853));
    InMux I__9320 (
            .O(N__52895),
            .I(N__52848));
    InMux I__9319 (
            .O(N__52894),
            .I(N__52848));
    InMux I__9318 (
            .O(N__52893),
            .I(N__52841));
    InMux I__9317 (
            .O(N__52892),
            .I(N__52841));
    InMux I__9316 (
            .O(N__52891),
            .I(N__52841));
    InMux I__9315 (
            .O(N__52890),
            .I(N__52838));
    InMux I__9314 (
            .O(N__52889),
            .I(N__52833));
    InMux I__9313 (
            .O(N__52888),
            .I(N__52833));
    InMux I__9312 (
            .O(N__52887),
            .I(N__52830));
    InMux I__9311 (
            .O(N__52886),
            .I(N__52825));
    InMux I__9310 (
            .O(N__52885),
            .I(N__52825));
    InMux I__9309 (
            .O(N__52884),
            .I(N__52818));
    InMux I__9308 (
            .O(N__52883),
            .I(N__52818));
    InMux I__9307 (
            .O(N__52882),
            .I(N__52818));
    InMux I__9306 (
            .O(N__52881),
            .I(N__52813));
    InMux I__9305 (
            .O(N__52880),
            .I(N__52813));
    InMux I__9304 (
            .O(N__52879),
            .I(N__52806));
    InMux I__9303 (
            .O(N__52878),
            .I(N__52806));
    InMux I__9302 (
            .O(N__52877),
            .I(N__52806));
    LocalMux I__9301 (
            .O(N__52874),
            .I(N__52794));
    LocalMux I__9300 (
            .O(N__52869),
            .I(N__52794));
    InMux I__9299 (
            .O(N__52868),
            .I(N__52791));
    InMux I__9298 (
            .O(N__52867),
            .I(N__52782));
    InMux I__9297 (
            .O(N__52866),
            .I(N__52782));
    InMux I__9296 (
            .O(N__52865),
            .I(N__52782));
    InMux I__9295 (
            .O(N__52864),
            .I(N__52782));
    InMux I__9294 (
            .O(N__52863),
            .I(N__52771));
    InMux I__9293 (
            .O(N__52862),
            .I(N__52771));
    InMux I__9292 (
            .O(N__52861),
            .I(N__52771));
    InMux I__9291 (
            .O(N__52860),
            .I(N__52771));
    InMux I__9290 (
            .O(N__52859),
            .I(N__52771));
    LocalMux I__9289 (
            .O(N__52856),
            .I(N__52759));
    LocalMux I__9288 (
            .O(N__52853),
            .I(N__52759));
    LocalMux I__9287 (
            .O(N__52848),
            .I(N__52756));
    LocalMux I__9286 (
            .O(N__52841),
            .I(N__52743));
    LocalMux I__9285 (
            .O(N__52838),
            .I(N__52743));
    LocalMux I__9284 (
            .O(N__52833),
            .I(N__52743));
    LocalMux I__9283 (
            .O(N__52830),
            .I(N__52743));
    LocalMux I__9282 (
            .O(N__52825),
            .I(N__52743));
    LocalMux I__9281 (
            .O(N__52818),
            .I(N__52743));
    LocalMux I__9280 (
            .O(N__52813),
            .I(N__52738));
    LocalMux I__9279 (
            .O(N__52806),
            .I(N__52735));
    InMux I__9278 (
            .O(N__52805),
            .I(N__52720));
    InMux I__9277 (
            .O(N__52804),
            .I(N__52720));
    InMux I__9276 (
            .O(N__52803),
            .I(N__52720));
    InMux I__9275 (
            .O(N__52802),
            .I(N__52720));
    InMux I__9274 (
            .O(N__52801),
            .I(N__52720));
    InMux I__9273 (
            .O(N__52800),
            .I(N__52720));
    InMux I__9272 (
            .O(N__52799),
            .I(N__52720));
    Span4Mux_h I__9271 (
            .O(N__52794),
            .I(N__52713));
    LocalMux I__9270 (
            .O(N__52791),
            .I(N__52713));
    LocalMux I__9269 (
            .O(N__52782),
            .I(N__52713));
    LocalMux I__9268 (
            .O(N__52771),
            .I(N__52708));
    InMux I__9267 (
            .O(N__52770),
            .I(N__52701));
    InMux I__9266 (
            .O(N__52769),
            .I(N__52701));
    InMux I__9265 (
            .O(N__52768),
            .I(N__52701));
    InMux I__9264 (
            .O(N__52767),
            .I(N__52692));
    InMux I__9263 (
            .O(N__52766),
            .I(N__52692));
    InMux I__9262 (
            .O(N__52765),
            .I(N__52692));
    InMux I__9261 (
            .O(N__52764),
            .I(N__52692));
    Span4Mux_h I__9260 (
            .O(N__52759),
            .I(N__52685));
    Span4Mux_s1_v I__9259 (
            .O(N__52756),
            .I(N__52685));
    Span4Mux_v I__9258 (
            .O(N__52743),
            .I(N__52685));
    InMux I__9257 (
            .O(N__52742),
            .I(N__52682));
    InMux I__9256 (
            .O(N__52741),
            .I(N__52674));
    Span12Mux_v I__9255 (
            .O(N__52738),
            .I(N__52671));
    Span4Mux_s2_v I__9254 (
            .O(N__52735),
            .I(N__52664));
    LocalMux I__9253 (
            .O(N__52720),
            .I(N__52664));
    Span4Mux_v I__9252 (
            .O(N__52713),
            .I(N__52664));
    InMux I__9251 (
            .O(N__52712),
            .I(N__52659));
    InMux I__9250 (
            .O(N__52711),
            .I(N__52659));
    Span4Mux_h I__9249 (
            .O(N__52708),
            .I(N__52648));
    LocalMux I__9248 (
            .O(N__52701),
            .I(N__52648));
    LocalMux I__9247 (
            .O(N__52692),
            .I(N__52648));
    Span4Mux_h I__9246 (
            .O(N__52685),
            .I(N__52648));
    LocalMux I__9245 (
            .O(N__52682),
            .I(N__52648));
    InMux I__9244 (
            .O(N__52681),
            .I(N__52637));
    InMux I__9243 (
            .O(N__52680),
            .I(N__52637));
    InMux I__9242 (
            .O(N__52679),
            .I(N__52637));
    InMux I__9241 (
            .O(N__52678),
            .I(N__52637));
    InMux I__9240 (
            .O(N__52677),
            .I(N__52637));
    LocalMux I__9239 (
            .O(N__52674),
            .I(\ppm_encoder_1.PPM_STATE_fast_RNICIABZ0Z_0 ));
    Odrv12 I__9238 (
            .O(N__52671),
            .I(\ppm_encoder_1.PPM_STATE_fast_RNICIABZ0Z_0 ));
    Odrv4 I__9237 (
            .O(N__52664),
            .I(\ppm_encoder_1.PPM_STATE_fast_RNICIABZ0Z_0 ));
    LocalMux I__9236 (
            .O(N__52659),
            .I(\ppm_encoder_1.PPM_STATE_fast_RNICIABZ0Z_0 ));
    Odrv4 I__9235 (
            .O(N__52648),
            .I(\ppm_encoder_1.PPM_STATE_fast_RNICIABZ0Z_0 ));
    LocalMux I__9234 (
            .O(N__52637),
            .I(\ppm_encoder_1.PPM_STATE_fast_RNICIABZ0Z_0 ));
    InMux I__9233 (
            .O(N__52624),
            .I(N__52619));
    InMux I__9232 (
            .O(N__52623),
            .I(N__52616));
    InMux I__9231 (
            .O(N__52622),
            .I(N__52613));
    LocalMux I__9230 (
            .O(N__52619),
            .I(N__52610));
    LocalMux I__9229 (
            .O(N__52616),
            .I(\ppm_encoder_1.counterZ0Z_0 ));
    LocalMux I__9228 (
            .O(N__52613),
            .I(\ppm_encoder_1.counterZ0Z_0 ));
    Odrv4 I__9227 (
            .O(N__52610),
            .I(\ppm_encoder_1.counterZ0Z_0 ));
    CascadeMux I__9226 (
            .O(N__52603),
            .I(N__52600));
    InMux I__9225 (
            .O(N__52600),
            .I(N__52595));
    InMux I__9224 (
            .O(N__52599),
            .I(N__52592));
    InMux I__9223 (
            .O(N__52598),
            .I(N__52589));
    LocalMux I__9222 (
            .O(N__52595),
            .I(N__52586));
    LocalMux I__9221 (
            .O(N__52592),
            .I(\ppm_encoder_1.counterZ0Z_1 ));
    LocalMux I__9220 (
            .O(N__52589),
            .I(\ppm_encoder_1.counterZ0Z_1 ));
    Odrv4 I__9219 (
            .O(N__52586),
            .I(\ppm_encoder_1.counterZ0Z_1 ));
    InMux I__9218 (
            .O(N__52579),
            .I(\ppm_encoder_1.un1_counter_13_cry_0 ));
    InMux I__9217 (
            .O(N__52576),
            .I(N__52572));
    InMux I__9216 (
            .O(N__52575),
            .I(N__52568));
    LocalMux I__9215 (
            .O(N__52572),
            .I(N__52565));
    InMux I__9214 (
            .O(N__52571),
            .I(N__52562));
    LocalMux I__9213 (
            .O(N__52568),
            .I(N__52557));
    Span4Mux_v I__9212 (
            .O(N__52565),
            .I(N__52557));
    LocalMux I__9211 (
            .O(N__52562),
            .I(\ppm_encoder_1.counterZ0Z_2 ));
    Odrv4 I__9210 (
            .O(N__52557),
            .I(\ppm_encoder_1.counterZ0Z_2 ));
    InMux I__9209 (
            .O(N__52552),
            .I(\ppm_encoder_1.un1_counter_13_cry_1 ));
    InMux I__9208 (
            .O(N__52549),
            .I(bfn_11_23_0_));
    InMux I__9207 (
            .O(N__52546),
            .I(N__52543));
    LocalMux I__9206 (
            .O(N__52543),
            .I(\pid_front.un11lto30_i_a2_0_and ));
    CascadeMux I__9205 (
            .O(N__52540),
            .I(\pid_front.un1_reset_i_a2_3_4_cascade_ ));
    CascadeMux I__9204 (
            .O(N__52537),
            .I(\pid_front.N_593_cascade_ ));
    InMux I__9203 (
            .O(N__52534),
            .I(N__52530));
    InMux I__9202 (
            .O(N__52533),
            .I(N__52527));
    LocalMux I__9201 (
            .O(N__52530),
            .I(N__52522));
    LocalMux I__9200 (
            .O(N__52527),
            .I(N__52522));
    Sp12to4 I__9199 (
            .O(N__52522),
            .I(N__52519));
    Span12Mux_s10_v I__9198 (
            .O(N__52519),
            .I(N__52516));
    Span12Mux_v I__9197 (
            .O(N__52516),
            .I(N__52513));
    Odrv12 I__9196 (
            .O(N__52513),
            .I(front_order_5));
    InMux I__9195 (
            .O(N__52510),
            .I(N__52507));
    LocalMux I__9194 (
            .O(N__52507),
            .I(N__52504));
    Odrv4 I__9193 (
            .O(N__52504),
            .I(\pid_front.N_11_i ));
    InMux I__9192 (
            .O(N__52501),
            .I(N__52498));
    LocalMux I__9191 (
            .O(N__52498),
            .I(\dron_frame_decoder_1.drone_H_disp_front_6 ));
    InMux I__9190 (
            .O(N__52495),
            .I(N__52492));
    LocalMux I__9189 (
            .O(N__52492),
            .I(drone_H_disp_front_1));
    InMux I__9188 (
            .O(N__52489),
            .I(N__52486));
    LocalMux I__9187 (
            .O(N__52486),
            .I(\dron_frame_decoder_1.drone_altitude_11 ));
    InMux I__9186 (
            .O(N__52483),
            .I(N__52480));
    LocalMux I__9185 (
            .O(N__52480),
            .I(N__52477));
    Span4Mux_h I__9184 (
            .O(N__52477),
            .I(N__52474));
    Odrv4 I__9183 (
            .O(N__52474),
            .I(drone_altitude_i_11));
    InMux I__9182 (
            .O(N__52471),
            .I(N__52468));
    LocalMux I__9181 (
            .O(N__52468),
            .I(\dron_frame_decoder_1.drone_H_disp_front_5 ));
    CascadeMux I__9180 (
            .O(N__52465),
            .I(N__52458));
    InMux I__9179 (
            .O(N__52464),
            .I(N__52454));
    InMux I__9178 (
            .O(N__52463),
            .I(N__52445));
    InMux I__9177 (
            .O(N__52462),
            .I(N__52445));
    InMux I__9176 (
            .O(N__52461),
            .I(N__52445));
    InMux I__9175 (
            .O(N__52458),
            .I(N__52445));
    InMux I__9174 (
            .O(N__52457),
            .I(N__52442));
    LocalMux I__9173 (
            .O(N__52454),
            .I(N__52439));
    LocalMux I__9172 (
            .O(N__52445),
            .I(N__52436));
    LocalMux I__9171 (
            .O(N__52442),
            .I(N__52433));
    Span4Mux_h I__9170 (
            .O(N__52439),
            .I(N__52430));
    Odrv4 I__9169 (
            .O(N__52436),
            .I(\Commands_frame_decoder.un1_sink_data_valid_2_0 ));
    Odrv12 I__9168 (
            .O(N__52433),
            .I(\Commands_frame_decoder.un1_sink_data_valid_2_0 ));
    Odrv4 I__9167 (
            .O(N__52430),
            .I(\Commands_frame_decoder.un1_sink_data_valid_2_0 ));
    InMux I__9166 (
            .O(N__52423),
            .I(N__52420));
    LocalMux I__9165 (
            .O(N__52420),
            .I(N__52416));
    InMux I__9164 (
            .O(N__52419),
            .I(N__52413));
    Span4Mux_v I__9163 (
            .O(N__52416),
            .I(N__52410));
    LocalMux I__9162 (
            .O(N__52413),
            .I(\Commands_frame_decoder.stateZ0Z_3 ));
    Odrv4 I__9161 (
            .O(N__52410),
            .I(\Commands_frame_decoder.stateZ0Z_3 ));
    InMux I__9160 (
            .O(N__52405),
            .I(N__52402));
    LocalMux I__9159 (
            .O(N__52402),
            .I(N__52398));
    InMux I__9158 (
            .O(N__52401),
            .I(N__52395));
    Span4Mux_v I__9157 (
            .O(N__52398),
            .I(N__52390));
    LocalMux I__9156 (
            .O(N__52395),
            .I(N__52390));
    Span4Mux_h I__9155 (
            .O(N__52390),
            .I(N__52387));
    Odrv4 I__9154 (
            .O(N__52387),
            .I(\Commands_frame_decoder.source_CH2data_1_sqmuxa ));
    CascadeMux I__9153 (
            .O(N__52384),
            .I(N__52381));
    InMux I__9152 (
            .O(N__52381),
            .I(N__52375));
    InMux I__9151 (
            .O(N__52380),
            .I(N__52375));
    LocalMux I__9150 (
            .O(N__52375),
            .I(\Commands_frame_decoder.stateZ0Z_4 ));
    InMux I__9149 (
            .O(N__52372),
            .I(N__52369));
    LocalMux I__9148 (
            .O(N__52369),
            .I(N__52366));
    Span4Mux_h I__9147 (
            .O(N__52366),
            .I(N__52363));
    Span4Mux_h I__9146 (
            .O(N__52363),
            .I(N__52360));
    Odrv4 I__9145 (
            .O(N__52360),
            .I(\pid_alt.error_axbZ0Z_13 ));
    InMux I__9144 (
            .O(N__52357),
            .I(N__52354));
    LocalMux I__9143 (
            .O(N__52354),
            .I(drone_altitude_13));
    InMux I__9142 (
            .O(N__52351),
            .I(N__52348));
    LocalMux I__9141 (
            .O(N__52348),
            .I(N__52345));
    Span4Mux_h I__9140 (
            .O(N__52345),
            .I(N__52342));
    Span4Mux_h I__9139 (
            .O(N__52342),
            .I(N__52339));
    Odrv4 I__9138 (
            .O(N__52339),
            .I(\pid_alt.error_axbZ0Z_14 ));
    InMux I__9137 (
            .O(N__52336),
            .I(N__52333));
    LocalMux I__9136 (
            .O(N__52333),
            .I(drone_altitude_14));
    CEMux I__9135 (
            .O(N__52330),
            .I(N__52326));
    CEMux I__9134 (
            .O(N__52329),
            .I(N__52323));
    LocalMux I__9133 (
            .O(N__52326),
            .I(N__52320));
    LocalMux I__9132 (
            .O(N__52323),
            .I(N__52317));
    Span4Mux_v I__9131 (
            .O(N__52320),
            .I(N__52314));
    Span4Mux_v I__9130 (
            .O(N__52317),
            .I(N__52311));
    Odrv4 I__9129 (
            .O(N__52314),
            .I(\dron_frame_decoder_1.N_732_0 ));
    Odrv4 I__9128 (
            .O(N__52311),
            .I(\dron_frame_decoder_1.N_732_0 ));
    InMux I__9127 (
            .O(N__52306),
            .I(N__52303));
    LocalMux I__9126 (
            .O(N__52303),
            .I(drone_altitude_2));
    InMux I__9125 (
            .O(N__52300),
            .I(N__52297));
    LocalMux I__9124 (
            .O(N__52297),
            .I(N__52294));
    Odrv12 I__9123 (
            .O(N__52294),
            .I(\pid_alt.error_axbZ0Z_2 ));
    InMux I__9122 (
            .O(N__52291),
            .I(N__52288));
    LocalMux I__9121 (
            .O(N__52288),
            .I(drone_altitude_3));
    InMux I__9120 (
            .O(N__52285),
            .I(N__52282));
    LocalMux I__9119 (
            .O(N__52282),
            .I(N__52279));
    Odrv12 I__9118 (
            .O(N__52279),
            .I(\pid_alt.error_axbZ0Z_3 ));
    InMux I__9117 (
            .O(N__52276),
            .I(N__52273));
    LocalMux I__9116 (
            .O(N__52273),
            .I(\dron_frame_decoder_1.drone_H_disp_side_8 ));
    InMux I__9115 (
            .O(N__52270),
            .I(N__52267));
    LocalMux I__9114 (
            .O(N__52267),
            .I(\dron_frame_decoder_1.drone_H_disp_side_9 ));
    CEMux I__9113 (
            .O(N__52264),
            .I(N__52261));
    LocalMux I__9112 (
            .O(N__52261),
            .I(N__52258));
    Span4Mux_v I__9111 (
            .O(N__52258),
            .I(N__52255));
    Span4Mux_v I__9110 (
            .O(N__52255),
            .I(N__52252));
    Odrv4 I__9109 (
            .O(N__52252),
            .I(\dron_frame_decoder_1.N_716_0 ));
    IoInMux I__9108 (
            .O(N__52249),
            .I(N__52246));
    LocalMux I__9107 (
            .O(N__52246),
            .I(N__52243));
    IoSpan4Mux I__9106 (
            .O(N__52243),
            .I(N__52238));
    InMux I__9105 (
            .O(N__52242),
            .I(N__52231));
    InMux I__9104 (
            .O(N__52241),
            .I(N__52226));
    Span4Mux_s1_v I__9103 (
            .O(N__52238),
            .I(N__52222));
    InMux I__9102 (
            .O(N__52237),
            .I(N__52219));
    CascadeMux I__9101 (
            .O(N__52236),
            .I(N__52216));
    CascadeMux I__9100 (
            .O(N__52235),
            .I(N__52213));
    CascadeMux I__9099 (
            .O(N__52234),
            .I(N__52210));
    LocalMux I__9098 (
            .O(N__52231),
            .I(N__52203));
    InMux I__9097 (
            .O(N__52230),
            .I(N__52200));
    InMux I__9096 (
            .O(N__52229),
            .I(N__52197));
    LocalMux I__9095 (
            .O(N__52226),
            .I(N__52194));
    InMux I__9094 (
            .O(N__52225),
            .I(N__52191));
    Sp12to4 I__9093 (
            .O(N__52222),
            .I(N__52188));
    LocalMux I__9092 (
            .O(N__52219),
            .I(N__52185));
    InMux I__9091 (
            .O(N__52216),
            .I(N__52170));
    InMux I__9090 (
            .O(N__52213),
            .I(N__52170));
    InMux I__9089 (
            .O(N__52210),
            .I(N__52170));
    InMux I__9088 (
            .O(N__52209),
            .I(N__52170));
    InMux I__9087 (
            .O(N__52208),
            .I(N__52170));
    InMux I__9086 (
            .O(N__52207),
            .I(N__52170));
    InMux I__9085 (
            .O(N__52206),
            .I(N__52170));
    Span4Mux_h I__9084 (
            .O(N__52203),
            .I(N__52167));
    LocalMux I__9083 (
            .O(N__52200),
            .I(N__52164));
    LocalMux I__9082 (
            .O(N__52197),
            .I(N__52157));
    Span4Mux_v I__9081 (
            .O(N__52194),
            .I(N__52157));
    LocalMux I__9080 (
            .O(N__52191),
            .I(N__52157));
    Span12Mux_v I__9079 (
            .O(N__52188),
            .I(N__52154));
    Span4Mux_h I__9078 (
            .O(N__52185),
            .I(N__52151));
    LocalMux I__9077 (
            .O(N__52170),
            .I(N__52146));
    Span4Mux_h I__9076 (
            .O(N__52167),
            .I(N__52146));
    Span4Mux_v I__9075 (
            .O(N__52164),
            .I(N__52141));
    Span4Mux_v I__9074 (
            .O(N__52157),
            .I(N__52141));
    Odrv12 I__9073 (
            .O(N__52154),
            .I(debug_CH2_18A_c));
    Odrv4 I__9072 (
            .O(N__52151),
            .I(debug_CH2_18A_c));
    Odrv4 I__9071 (
            .O(N__52146),
            .I(debug_CH2_18A_c));
    Odrv4 I__9070 (
            .O(N__52141),
            .I(debug_CH2_18A_c));
    InMux I__9069 (
            .O(N__52132),
            .I(N__52129));
    LocalMux I__9068 (
            .O(N__52129),
            .I(N__52126));
    Span4Mux_v I__9067 (
            .O(N__52126),
            .I(N__52120));
    InMux I__9066 (
            .O(N__52125),
            .I(N__52113));
    InMux I__9065 (
            .O(N__52124),
            .I(N__52113));
    InMux I__9064 (
            .O(N__52123),
            .I(N__52113));
    Odrv4 I__9063 (
            .O(N__52120),
            .I(\uart_pc.data_rdyc_1 ));
    LocalMux I__9062 (
            .O(N__52113),
            .I(\uart_pc.data_rdyc_1 ));
    InMux I__9061 (
            .O(N__52108),
            .I(N__52102));
    InMux I__9060 (
            .O(N__52107),
            .I(N__52099));
    InMux I__9059 (
            .O(N__52106),
            .I(N__52094));
    InMux I__9058 (
            .O(N__52105),
            .I(N__52094));
    LocalMux I__9057 (
            .O(N__52102),
            .I(N__52091));
    LocalMux I__9056 (
            .O(N__52099),
            .I(N__52088));
    LocalMux I__9055 (
            .O(N__52094),
            .I(\Commands_frame_decoder.stateZ0Z_6 ));
    Odrv4 I__9054 (
            .O(N__52091),
            .I(\Commands_frame_decoder.stateZ0Z_6 ));
    Odrv12 I__9053 (
            .O(N__52088),
            .I(\Commands_frame_decoder.stateZ0Z_6 ));
    InMux I__9052 (
            .O(N__52081),
            .I(N__52078));
    LocalMux I__9051 (
            .O(N__52078),
            .I(N__52075));
    Span4Mux_v I__9050 (
            .O(N__52075),
            .I(N__52072));
    Sp12to4 I__9049 (
            .O(N__52072),
            .I(N__52068));
    InMux I__9048 (
            .O(N__52071),
            .I(N__52065));
    Span12Mux_s11_h I__9047 (
            .O(N__52068),
            .I(N__52062));
    LocalMux I__9046 (
            .O(N__52065),
            .I(alt_kp_4));
    Odrv12 I__9045 (
            .O(N__52062),
            .I(alt_kp_4));
    CascadeMux I__9044 (
            .O(N__52057),
            .I(N__52053));
    CascadeMux I__9043 (
            .O(N__52056),
            .I(N__52050));
    InMux I__9042 (
            .O(N__52053),
            .I(N__52046));
    InMux I__9041 (
            .O(N__52050),
            .I(N__52040));
    InMux I__9040 (
            .O(N__52049),
            .I(N__52040));
    LocalMux I__9039 (
            .O(N__52046),
            .I(N__52037));
    InMux I__9038 (
            .O(N__52045),
            .I(N__52034));
    LocalMux I__9037 (
            .O(N__52040),
            .I(\Commands_frame_decoder.stateZ0Z_7 ));
    Odrv4 I__9036 (
            .O(N__52037),
            .I(\Commands_frame_decoder.stateZ0Z_7 ));
    LocalMux I__9035 (
            .O(N__52034),
            .I(\Commands_frame_decoder.stateZ0Z_7 ));
    InMux I__9034 (
            .O(N__52027),
            .I(N__52024));
    LocalMux I__9033 (
            .O(N__52024),
            .I(N__52021));
    Span4Mux_v I__9032 (
            .O(N__52021),
            .I(N__52018));
    Span4Mux_v I__9031 (
            .O(N__52018),
            .I(N__52014));
    InMux I__9030 (
            .O(N__52017),
            .I(N__52011));
    Sp12to4 I__9029 (
            .O(N__52014),
            .I(N__52007));
    LocalMux I__9028 (
            .O(N__52011),
            .I(N__52004));
    InMux I__9027 (
            .O(N__52010),
            .I(N__52001));
    Span12Mux_h I__9026 (
            .O(N__52007),
            .I(N__51996));
    Span12Mux_s11_h I__9025 (
            .O(N__52004),
            .I(N__51996));
    LocalMux I__9024 (
            .O(N__52001),
            .I(xy_kp_4));
    Odrv12 I__9023 (
            .O(N__51996),
            .I(xy_kp_4));
    InMux I__9022 (
            .O(N__51991),
            .I(N__51987));
    InMux I__9021 (
            .O(N__51990),
            .I(N__51984));
    LocalMux I__9020 (
            .O(N__51987),
            .I(N__51981));
    LocalMux I__9019 (
            .O(N__51984),
            .I(\reset_module_System.countZ0Z_17 ));
    Odrv4 I__9018 (
            .O(N__51981),
            .I(\reset_module_System.countZ0Z_17 ));
    InMux I__9017 (
            .O(N__51976),
            .I(bfn_11_15_0_));
    InMux I__9016 (
            .O(N__51973),
            .I(N__51969));
    InMux I__9015 (
            .O(N__51972),
            .I(N__51966));
    LocalMux I__9014 (
            .O(N__51969),
            .I(N__51963));
    LocalMux I__9013 (
            .O(N__51966),
            .I(\reset_module_System.countZ0Z_18 ));
    Odrv4 I__9012 (
            .O(N__51963),
            .I(\reset_module_System.countZ0Z_18 ));
    InMux I__9011 (
            .O(N__51958),
            .I(\reset_module_System.count_1_cry_17 ));
    InMux I__9010 (
            .O(N__51955),
            .I(\reset_module_System.count_1_cry_18 ));
    InMux I__9009 (
            .O(N__51952),
            .I(\reset_module_System.count_1_cry_19 ));
    InMux I__9008 (
            .O(N__51949),
            .I(\reset_module_System.count_1_cry_20 ));
    InMux I__9007 (
            .O(N__51946),
            .I(N__51943));
    LocalMux I__9006 (
            .O(N__51943),
            .I(\dron_frame_decoder_1.drone_H_disp_side_7 ));
    InMux I__9005 (
            .O(N__51940),
            .I(N__51936));
    InMux I__9004 (
            .O(N__51939),
            .I(N__51933));
    LocalMux I__9003 (
            .O(N__51936),
            .I(N__51930));
    LocalMux I__9002 (
            .O(N__51933),
            .I(\Commands_frame_decoder.source_CH4data_1_sqmuxa ));
    Odrv4 I__9001 (
            .O(N__51930),
            .I(\Commands_frame_decoder.source_CH4data_1_sqmuxa ));
    InMux I__9000 (
            .O(N__51925),
            .I(N__51922));
    LocalMux I__8999 (
            .O(N__51922),
            .I(\dron_frame_decoder_1.drone_H_disp_side_10 ));
    InMux I__8998 (
            .O(N__51919),
            .I(\reset_module_System.count_1_cry_7 ));
    CascadeMux I__8997 (
            .O(N__51916),
            .I(N__51913));
    InMux I__8996 (
            .O(N__51913),
            .I(N__51909));
    InMux I__8995 (
            .O(N__51912),
            .I(N__51906));
    LocalMux I__8994 (
            .O(N__51909),
            .I(N__51903));
    LocalMux I__8993 (
            .O(N__51906),
            .I(\reset_module_System.countZ0Z_9 ));
    Odrv4 I__8992 (
            .O(N__51903),
            .I(\reset_module_System.countZ0Z_9 ));
    InMux I__8991 (
            .O(N__51898),
            .I(bfn_11_14_0_));
    InMux I__8990 (
            .O(N__51895),
            .I(N__51891));
    InMux I__8989 (
            .O(N__51894),
            .I(N__51888));
    LocalMux I__8988 (
            .O(N__51891),
            .I(N__51885));
    LocalMux I__8987 (
            .O(N__51888),
            .I(\reset_module_System.countZ0Z_10 ));
    Odrv4 I__8986 (
            .O(N__51885),
            .I(\reset_module_System.countZ0Z_10 ));
    InMux I__8985 (
            .O(N__51880),
            .I(\reset_module_System.count_1_cry_9 ));
    InMux I__8984 (
            .O(N__51877),
            .I(N__51873));
    InMux I__8983 (
            .O(N__51876),
            .I(N__51870));
    LocalMux I__8982 (
            .O(N__51873),
            .I(N__51867));
    LocalMux I__8981 (
            .O(N__51870),
            .I(\reset_module_System.countZ0Z_11 ));
    Odrv4 I__8980 (
            .O(N__51867),
            .I(\reset_module_System.countZ0Z_11 ));
    InMux I__8979 (
            .O(N__51862),
            .I(\reset_module_System.count_1_cry_10 ));
    CascadeMux I__8978 (
            .O(N__51859),
            .I(N__51856));
    InMux I__8977 (
            .O(N__51856),
            .I(N__51853));
    LocalMux I__8976 (
            .O(N__51853),
            .I(N__51849));
    InMux I__8975 (
            .O(N__51852),
            .I(N__51846));
    Odrv4 I__8974 (
            .O(N__51849),
            .I(\reset_module_System.countZ0Z_12 ));
    LocalMux I__8973 (
            .O(N__51846),
            .I(\reset_module_System.countZ0Z_12 ));
    InMux I__8972 (
            .O(N__51841),
            .I(\reset_module_System.count_1_cry_11 ));
    InMux I__8971 (
            .O(N__51838),
            .I(\reset_module_System.count_1_cry_12 ));
    InMux I__8970 (
            .O(N__51835),
            .I(N__51831));
    InMux I__8969 (
            .O(N__51834),
            .I(N__51828));
    LocalMux I__8968 (
            .O(N__51831),
            .I(N__51825));
    LocalMux I__8967 (
            .O(N__51828),
            .I(\reset_module_System.countZ0Z_14 ));
    Odrv4 I__8966 (
            .O(N__51825),
            .I(\reset_module_System.countZ0Z_14 ));
    InMux I__8965 (
            .O(N__51820),
            .I(\reset_module_System.count_1_cry_13 ));
    InMux I__8964 (
            .O(N__51817),
            .I(\reset_module_System.count_1_cry_14 ));
    CascadeMux I__8963 (
            .O(N__51814),
            .I(N__51811));
    InMux I__8962 (
            .O(N__51811),
            .I(N__51808));
    LocalMux I__8961 (
            .O(N__51808),
            .I(N__51804));
    InMux I__8960 (
            .O(N__51807),
            .I(N__51801));
    Odrv4 I__8959 (
            .O(N__51804),
            .I(\reset_module_System.countZ0Z_16 ));
    LocalMux I__8958 (
            .O(N__51801),
            .I(\reset_module_System.countZ0Z_16 ));
    InMux I__8957 (
            .O(N__51796),
            .I(\reset_module_System.count_1_cry_15 ));
    CascadeMux I__8956 (
            .O(N__51793),
            .I(\reset_module_System.reset6_13_cascade_ ));
    InMux I__8955 (
            .O(N__51790),
            .I(N__51787));
    LocalMux I__8954 (
            .O(N__51787),
            .I(\reset_module_System.reset6_3 ));
    InMux I__8953 (
            .O(N__51784),
            .I(N__51781));
    LocalMux I__8952 (
            .O(N__51781),
            .I(\reset_module_System.reset6_17 ));
    CascadeMux I__8951 (
            .O(N__51778),
            .I(N__51774));
    InMux I__8950 (
            .O(N__51777),
            .I(N__51765));
    InMux I__8949 (
            .O(N__51774),
            .I(N__51765));
    InMux I__8948 (
            .O(N__51773),
            .I(N__51765));
    InMux I__8947 (
            .O(N__51772),
            .I(N__51762));
    LocalMux I__8946 (
            .O(N__51765),
            .I(\reset_module_System.countZ0Z_0 ));
    LocalMux I__8945 (
            .O(N__51762),
            .I(\reset_module_System.countZ0Z_0 ));
    CascadeMux I__8944 (
            .O(N__51757),
            .I(N__51754));
    InMux I__8943 (
            .O(N__51754),
            .I(N__51749));
    InMux I__8942 (
            .O(N__51753),
            .I(N__51744));
    InMux I__8941 (
            .O(N__51752),
            .I(N__51744));
    LocalMux I__8940 (
            .O(N__51749),
            .I(N__51741));
    LocalMux I__8939 (
            .O(N__51744),
            .I(\reset_module_System.countZ0Z_1 ));
    Odrv4 I__8938 (
            .O(N__51741),
            .I(\reset_module_System.countZ0Z_1 ));
    InMux I__8937 (
            .O(N__51736),
            .I(\reset_module_System.count_1_cry_1 ));
    InMux I__8936 (
            .O(N__51733),
            .I(\reset_module_System.count_1_cry_2 ));
    InMux I__8935 (
            .O(N__51730),
            .I(N__51726));
    InMux I__8934 (
            .O(N__51729),
            .I(N__51723));
    LocalMux I__8933 (
            .O(N__51726),
            .I(\reset_module_System.countZ0Z_4 ));
    LocalMux I__8932 (
            .O(N__51723),
            .I(\reset_module_System.countZ0Z_4 ));
    InMux I__8931 (
            .O(N__51718),
            .I(\reset_module_System.count_1_cry_3 ));
    InMux I__8930 (
            .O(N__51715),
            .I(N__51711));
    InMux I__8929 (
            .O(N__51714),
            .I(N__51708));
    LocalMux I__8928 (
            .O(N__51711),
            .I(\reset_module_System.countZ0Z_5 ));
    LocalMux I__8927 (
            .O(N__51708),
            .I(\reset_module_System.countZ0Z_5 ));
    InMux I__8926 (
            .O(N__51703),
            .I(\reset_module_System.count_1_cry_4 ));
    InMux I__8925 (
            .O(N__51700),
            .I(\reset_module_System.count_1_cry_5 ));
    InMux I__8924 (
            .O(N__51697),
            .I(N__51693));
    InMux I__8923 (
            .O(N__51696),
            .I(N__51690));
    LocalMux I__8922 (
            .O(N__51693),
            .I(\reset_module_System.countZ0Z_7 ));
    LocalMux I__8921 (
            .O(N__51690),
            .I(\reset_module_System.countZ0Z_7 ));
    InMux I__8920 (
            .O(N__51685),
            .I(\reset_module_System.count_1_cry_6 ));
    InMux I__8919 (
            .O(N__51682),
            .I(N__51678));
    InMux I__8918 (
            .O(N__51681),
            .I(N__51675));
    LocalMux I__8917 (
            .O(N__51678),
            .I(\reset_module_System.countZ0Z_8 ));
    LocalMux I__8916 (
            .O(N__51675),
            .I(\reset_module_System.countZ0Z_8 ));
    CascadeMux I__8915 (
            .O(N__51670),
            .I(N__51667));
    InMux I__8914 (
            .O(N__51667),
            .I(N__51664));
    LocalMux I__8913 (
            .O(N__51664),
            .I(\uart_drone.un1_state_2_0_a3_0 ));
    CascadeMux I__8912 (
            .O(N__51661),
            .I(\reset_module_System.count_1_1_cascade_ ));
    CascadeMux I__8911 (
            .O(N__51658),
            .I(\reset_module_System.reset6_19_cascade_ ));
    IoInMux I__8910 (
            .O(N__51655),
            .I(N__51652));
    LocalMux I__8909 (
            .O(N__51652),
            .I(N__51649));
    Span4Mux_s1_v I__8908 (
            .O(N__51649),
            .I(N__51646));
    Sp12to4 I__8907 (
            .O(N__51646),
            .I(N__51643));
    Span12Mux_h I__8906 (
            .O(N__51643),
            .I(N__51640));
    Span12Mux_v I__8905 (
            .O(N__51640),
            .I(N__51637));
    Odrv12 I__8904 (
            .O(N__51637),
            .I(\reset_module_System.reset_isoZ0 ));
    CascadeMux I__8903 (
            .O(N__51634),
            .I(\uart_drone.state_srsts_i_0_2_cascade_ ));
    InMux I__8902 (
            .O(N__51631),
            .I(N__51627));
    CascadeMux I__8901 (
            .O(N__51630),
            .I(N__51623));
    LocalMux I__8900 (
            .O(N__51627),
            .I(N__51620));
    InMux I__8899 (
            .O(N__51626),
            .I(N__51615));
    InMux I__8898 (
            .O(N__51623),
            .I(N__51615));
    Span4Mux_v I__8897 (
            .O(N__51620),
            .I(N__51612));
    LocalMux I__8896 (
            .O(N__51615),
            .I(\Commands_frame_decoder.stateZ0Z_11 ));
    Odrv4 I__8895 (
            .O(N__51612),
            .I(\Commands_frame_decoder.stateZ0Z_11 ));
    CEMux I__8894 (
            .O(N__51607),
            .I(N__51604));
    LocalMux I__8893 (
            .O(N__51604),
            .I(N__51601));
    Span4Mux_v I__8892 (
            .O(N__51601),
            .I(N__51598));
    Sp12to4 I__8891 (
            .O(N__51598),
            .I(N__51595));
    Odrv12 I__8890 (
            .O(N__51595),
            .I(\Commands_frame_decoder.state_RNIRSI31Z0Z_11 ));
    CascadeMux I__8889 (
            .O(N__51592),
            .I(N__51586));
    InMux I__8888 (
            .O(N__51591),
            .I(N__51583));
    InMux I__8887 (
            .O(N__51590),
            .I(N__51578));
    InMux I__8886 (
            .O(N__51589),
            .I(N__51578));
    InMux I__8885 (
            .O(N__51586),
            .I(N__51575));
    LocalMux I__8884 (
            .O(N__51583),
            .I(\uart_drone.stateZ0Z_2 ));
    LocalMux I__8883 (
            .O(N__51578),
            .I(\uart_drone.stateZ0Z_2 ));
    LocalMux I__8882 (
            .O(N__51575),
            .I(\uart_drone.stateZ0Z_2 ));
    CascadeMux I__8881 (
            .O(N__51568),
            .I(N__51564));
    CascadeMux I__8880 (
            .O(N__51567),
            .I(N__51558));
    InMux I__8879 (
            .O(N__51564),
            .I(N__51555));
    InMux I__8878 (
            .O(N__51563),
            .I(N__51552));
    CascadeMux I__8877 (
            .O(N__51562),
            .I(N__51549));
    InMux I__8876 (
            .O(N__51561),
            .I(N__51544));
    InMux I__8875 (
            .O(N__51558),
            .I(N__51544));
    LocalMux I__8874 (
            .O(N__51555),
            .I(N__51539));
    LocalMux I__8873 (
            .O(N__51552),
            .I(N__51539));
    InMux I__8872 (
            .O(N__51549),
            .I(N__51536));
    LocalMux I__8871 (
            .O(N__51544),
            .I(N__51533));
    Span4Mux_v I__8870 (
            .O(N__51539),
            .I(N__51530));
    LocalMux I__8869 (
            .O(N__51536),
            .I(N__51527));
    Odrv4 I__8868 (
            .O(N__51533),
            .I(\uart_drone.timer_Count_0_sqmuxa ));
    Odrv4 I__8867 (
            .O(N__51530),
            .I(\uart_drone.timer_Count_0_sqmuxa ));
    Odrv4 I__8866 (
            .O(N__51527),
            .I(\uart_drone.timer_Count_0_sqmuxa ));
    InMux I__8865 (
            .O(N__51520),
            .I(N__51515));
    InMux I__8864 (
            .O(N__51519),
            .I(N__51510));
    InMux I__8863 (
            .O(N__51518),
            .I(N__51506));
    LocalMux I__8862 (
            .O(N__51515),
            .I(N__51503));
    InMux I__8861 (
            .O(N__51514),
            .I(N__51498));
    InMux I__8860 (
            .O(N__51513),
            .I(N__51498));
    LocalMux I__8859 (
            .O(N__51510),
            .I(N__51493));
    InMux I__8858 (
            .O(N__51509),
            .I(N__51490));
    LocalMux I__8857 (
            .O(N__51506),
            .I(N__51483));
    Span4Mux_h I__8856 (
            .O(N__51503),
            .I(N__51483));
    LocalMux I__8855 (
            .O(N__51498),
            .I(N__51483));
    InMux I__8854 (
            .O(N__51497),
            .I(N__51478));
    InMux I__8853 (
            .O(N__51496),
            .I(N__51478));
    Odrv12 I__8852 (
            .O(N__51493),
            .I(\uart_drone.timer_CountZ1Z_3 ));
    LocalMux I__8851 (
            .O(N__51490),
            .I(\uart_drone.timer_CountZ1Z_3 ));
    Odrv4 I__8850 (
            .O(N__51483),
            .I(\uart_drone.timer_CountZ1Z_3 ));
    LocalMux I__8849 (
            .O(N__51478),
            .I(\uart_drone.timer_CountZ1Z_3 ));
    InMux I__8848 (
            .O(N__51469),
            .I(N__51463));
    InMux I__8847 (
            .O(N__51468),
            .I(N__51463));
    LocalMux I__8846 (
            .O(N__51463),
            .I(N__51460));
    Span4Mux_h I__8845 (
            .O(N__51460),
            .I(N__51455));
    InMux I__8844 (
            .O(N__51459),
            .I(N__51450));
    InMux I__8843 (
            .O(N__51458),
            .I(N__51450));
    Odrv4 I__8842 (
            .O(N__51455),
            .I(\uart_drone.un1_state_4_0 ));
    LocalMux I__8841 (
            .O(N__51450),
            .I(\uart_drone.un1_state_4_0 ));
    InMux I__8840 (
            .O(N__51445),
            .I(N__51442));
    LocalMux I__8839 (
            .O(N__51442),
            .I(N__51437));
    InMux I__8838 (
            .O(N__51441),
            .I(N__51432));
    InMux I__8837 (
            .O(N__51440),
            .I(N__51432));
    Odrv4 I__8836 (
            .O(N__51437),
            .I(\uart_drone.stateZ0Z_1 ));
    LocalMux I__8835 (
            .O(N__51432),
            .I(\uart_drone.stateZ0Z_1 ));
    InMux I__8834 (
            .O(N__51427),
            .I(N__51424));
    LocalMux I__8833 (
            .O(N__51424),
            .I(N__51421));
    Odrv4 I__8832 (
            .O(N__51421),
            .I(\uart_drone_sync.aux_2__0__0_0 ));
    InMux I__8831 (
            .O(N__51418),
            .I(N__51415));
    LocalMux I__8830 (
            .O(N__51415),
            .I(\uart_drone_sync.aux_3__0__0_0 ));
    InMux I__8829 (
            .O(N__51412),
            .I(N__51409));
    LocalMux I__8828 (
            .O(N__51409),
            .I(N__51406));
    Odrv4 I__8827 (
            .O(N__51406),
            .I(\ppm_encoder_1.un1_aileron_cry_12_THRU_CO ));
    CascadeMux I__8826 (
            .O(N__51403),
            .I(N__51399));
    InMux I__8825 (
            .O(N__51402),
            .I(N__51396));
    InMux I__8824 (
            .O(N__51399),
            .I(N__51393));
    LocalMux I__8823 (
            .O(N__51396),
            .I(N__51390));
    LocalMux I__8822 (
            .O(N__51393),
            .I(\ppm_encoder_1.aileronZ0Z_13 ));
    Odrv12 I__8821 (
            .O(N__51390),
            .I(\ppm_encoder_1.aileronZ0Z_13 ));
    InMux I__8820 (
            .O(N__51385),
            .I(N__51382));
    LocalMux I__8819 (
            .O(N__51382),
            .I(\ppm_encoder_1.un1_elevator_cry_4_THRU_CO ));
    CascadeMux I__8818 (
            .O(N__51379),
            .I(N__51375));
    InMux I__8817 (
            .O(N__51378),
            .I(N__51360));
    InMux I__8816 (
            .O(N__51375),
            .I(N__51360));
    CascadeMux I__8815 (
            .O(N__51374),
            .I(N__51347));
    CascadeMux I__8814 (
            .O(N__51373),
            .I(N__51341));
    CascadeMux I__8813 (
            .O(N__51372),
            .I(N__51338));
    CascadeMux I__8812 (
            .O(N__51371),
            .I(N__51335));
    CascadeMux I__8811 (
            .O(N__51370),
            .I(N__51332));
    CascadeMux I__8810 (
            .O(N__51369),
            .I(N__51329));
    CascadeMux I__8809 (
            .O(N__51368),
            .I(N__51324));
    CascadeMux I__8808 (
            .O(N__51367),
            .I(N__51314));
    CascadeMux I__8807 (
            .O(N__51366),
            .I(N__51311));
    CascadeMux I__8806 (
            .O(N__51365),
            .I(N__51308));
    LocalMux I__8805 (
            .O(N__51360),
            .I(N__51305));
    InMux I__8804 (
            .O(N__51359),
            .I(N__51298));
    InMux I__8803 (
            .O(N__51358),
            .I(N__51298));
    InMux I__8802 (
            .O(N__51357),
            .I(N__51298));
    CascadeMux I__8801 (
            .O(N__51356),
            .I(N__51292));
    CascadeMux I__8800 (
            .O(N__51355),
            .I(N__51289));
    CascadeMux I__8799 (
            .O(N__51354),
            .I(N__51282));
    CascadeMux I__8798 (
            .O(N__51353),
            .I(N__51279));
    CascadeMux I__8797 (
            .O(N__51352),
            .I(N__51275));
    CascadeMux I__8796 (
            .O(N__51351),
            .I(N__51272));
    CascadeMux I__8795 (
            .O(N__51350),
            .I(N__51268));
    InMux I__8794 (
            .O(N__51347),
            .I(N__51262));
    InMux I__8793 (
            .O(N__51346),
            .I(N__51262));
    InMux I__8792 (
            .O(N__51345),
            .I(N__51246));
    InMux I__8791 (
            .O(N__51344),
            .I(N__51246));
    InMux I__8790 (
            .O(N__51341),
            .I(N__51246));
    InMux I__8789 (
            .O(N__51338),
            .I(N__51246));
    InMux I__8788 (
            .O(N__51335),
            .I(N__51246));
    InMux I__8787 (
            .O(N__51332),
            .I(N__51246));
    InMux I__8786 (
            .O(N__51329),
            .I(N__51243));
    InMux I__8785 (
            .O(N__51328),
            .I(N__51238));
    InMux I__8784 (
            .O(N__51327),
            .I(N__51238));
    InMux I__8783 (
            .O(N__51324),
            .I(N__51235));
    CascadeMux I__8782 (
            .O(N__51323),
            .I(N__51231));
    CascadeMux I__8781 (
            .O(N__51322),
            .I(N__51228));
    CascadeMux I__8780 (
            .O(N__51321),
            .I(N__51225));
    InMux I__8779 (
            .O(N__51320),
            .I(N__51219));
    InMux I__8778 (
            .O(N__51319),
            .I(N__51206));
    InMux I__8777 (
            .O(N__51318),
            .I(N__51206));
    InMux I__8776 (
            .O(N__51317),
            .I(N__51206));
    InMux I__8775 (
            .O(N__51314),
            .I(N__51206));
    InMux I__8774 (
            .O(N__51311),
            .I(N__51206));
    InMux I__8773 (
            .O(N__51308),
            .I(N__51206));
    Span4Mux_s2_v I__8772 (
            .O(N__51305),
            .I(N__51201));
    LocalMux I__8771 (
            .O(N__51298),
            .I(N__51201));
    InMux I__8770 (
            .O(N__51297),
            .I(N__51190));
    InMux I__8769 (
            .O(N__51296),
            .I(N__51190));
    InMux I__8768 (
            .O(N__51295),
            .I(N__51190));
    InMux I__8767 (
            .O(N__51292),
            .I(N__51190));
    InMux I__8766 (
            .O(N__51289),
            .I(N__51190));
    InMux I__8765 (
            .O(N__51288),
            .I(N__51177));
    InMux I__8764 (
            .O(N__51287),
            .I(N__51177));
    InMux I__8763 (
            .O(N__51286),
            .I(N__51177));
    InMux I__8762 (
            .O(N__51285),
            .I(N__51177));
    InMux I__8761 (
            .O(N__51282),
            .I(N__51177));
    InMux I__8760 (
            .O(N__51279),
            .I(N__51177));
    InMux I__8759 (
            .O(N__51278),
            .I(N__51170));
    InMux I__8758 (
            .O(N__51275),
            .I(N__51170));
    InMux I__8757 (
            .O(N__51272),
            .I(N__51170));
    InMux I__8756 (
            .O(N__51271),
            .I(N__51163));
    InMux I__8755 (
            .O(N__51268),
            .I(N__51163));
    InMux I__8754 (
            .O(N__51267),
            .I(N__51163));
    LocalMux I__8753 (
            .O(N__51262),
            .I(N__51160));
    InMux I__8752 (
            .O(N__51261),
            .I(N__51155));
    InMux I__8751 (
            .O(N__51260),
            .I(N__51155));
    InMux I__8750 (
            .O(N__51259),
            .I(N__51152));
    LocalMux I__8749 (
            .O(N__51246),
            .I(N__51149));
    LocalMux I__8748 (
            .O(N__51243),
            .I(N__51144));
    LocalMux I__8747 (
            .O(N__51238),
            .I(N__51144));
    LocalMux I__8746 (
            .O(N__51235),
            .I(N__51141));
    InMux I__8745 (
            .O(N__51234),
            .I(N__51126));
    InMux I__8744 (
            .O(N__51231),
            .I(N__51126));
    InMux I__8743 (
            .O(N__51228),
            .I(N__51126));
    InMux I__8742 (
            .O(N__51225),
            .I(N__51126));
    InMux I__8741 (
            .O(N__51224),
            .I(N__51126));
    InMux I__8740 (
            .O(N__51223),
            .I(N__51126));
    InMux I__8739 (
            .O(N__51222),
            .I(N__51126));
    LocalMux I__8738 (
            .O(N__51219),
            .I(N__51119));
    LocalMux I__8737 (
            .O(N__51206),
            .I(N__51119));
    Span4Mux_v I__8736 (
            .O(N__51201),
            .I(N__51119));
    LocalMux I__8735 (
            .O(N__51190),
            .I(N__51116));
    LocalMux I__8734 (
            .O(N__51177),
            .I(N__51113));
    LocalMux I__8733 (
            .O(N__51170),
            .I(N__51104));
    LocalMux I__8732 (
            .O(N__51163),
            .I(N__51104));
    Span4Mux_v I__8731 (
            .O(N__51160),
            .I(N__51104));
    LocalMux I__8730 (
            .O(N__51155),
            .I(N__51104));
    LocalMux I__8729 (
            .O(N__51152),
            .I(N__51097));
    Span4Mux_v I__8728 (
            .O(N__51149),
            .I(N__51097));
    Span4Mux_v I__8727 (
            .O(N__51144),
            .I(N__51097));
    Span4Mux_v I__8726 (
            .O(N__51141),
            .I(N__51090));
    LocalMux I__8725 (
            .O(N__51126),
            .I(N__51090));
    Span4Mux_h I__8724 (
            .O(N__51119),
            .I(N__51090));
    Span4Mux_h I__8723 (
            .O(N__51116),
            .I(N__51087));
    Span4Mux_v I__8722 (
            .O(N__51113),
            .I(N__51082));
    Span4Mux_v I__8721 (
            .O(N__51104),
            .I(N__51082));
    Span4Mux_h I__8720 (
            .O(N__51097),
            .I(N__51079));
    Span4Mux_h I__8719 (
            .O(N__51090),
            .I(N__51076));
    Odrv4 I__8718 (
            .O(N__51087),
            .I(pid_altitude_dv));
    Odrv4 I__8717 (
            .O(N__51082),
            .I(pid_altitude_dv));
    Odrv4 I__8716 (
            .O(N__51079),
            .I(pid_altitude_dv));
    Odrv4 I__8715 (
            .O(N__51076),
            .I(pid_altitude_dv));
    InMux I__8714 (
            .O(N__51067),
            .I(N__51064));
    LocalMux I__8713 (
            .O(N__51064),
            .I(N__51060));
    CascadeMux I__8712 (
            .O(N__51063),
            .I(N__51057));
    Span4Mux_h I__8711 (
            .O(N__51060),
            .I(N__51054));
    InMux I__8710 (
            .O(N__51057),
            .I(N__51051));
    Span4Mux_v I__8709 (
            .O(N__51054),
            .I(N__51048));
    LocalMux I__8708 (
            .O(N__51051),
            .I(\ppm_encoder_1.elevatorZ0Z_5 ));
    Odrv4 I__8707 (
            .O(N__51048),
            .I(\ppm_encoder_1.elevatorZ0Z_5 ));
    InMux I__8706 (
            .O(N__51043),
            .I(N__51040));
    LocalMux I__8705 (
            .O(N__51040),
            .I(N__51037));
    Span4Mux_h I__8704 (
            .O(N__51037),
            .I(N__51034));
    Span4Mux_v I__8703 (
            .O(N__51034),
            .I(N__51031));
    Span4Mux_v I__8702 (
            .O(N__51031),
            .I(N__51028));
    Odrv4 I__8701 (
            .O(N__51028),
            .I(\uart_drone.timer_Count_RNO_0_0_1 ));
    InMux I__8700 (
            .O(N__51025),
            .I(N__51022));
    LocalMux I__8699 (
            .O(N__51022),
            .I(N__51019));
    Span4Mux_h I__8698 (
            .O(N__51019),
            .I(N__51015));
    InMux I__8697 (
            .O(N__51018),
            .I(N__51012));
    Span4Mux_v I__8696 (
            .O(N__51015),
            .I(N__51007));
    LocalMux I__8695 (
            .O(N__51012),
            .I(N__51007));
    Span4Mux_v I__8694 (
            .O(N__51007),
            .I(N__51004));
    Odrv4 I__8693 (
            .O(N__51004),
            .I(\uart_drone.timer_CountZ1Z_1 ));
    CascadeMux I__8692 (
            .O(N__51001),
            .I(\uart_drone.N_144_1_cascade_ ));
    InMux I__8691 (
            .O(N__50998),
            .I(N__50995));
    LocalMux I__8690 (
            .O(N__50995),
            .I(\uart_drone.N_145 ));
    InMux I__8689 (
            .O(N__50992),
            .I(N__50989));
    LocalMux I__8688 (
            .O(N__50989),
            .I(\ppm_encoder_1.N_436 ));
    InMux I__8687 (
            .O(N__50986),
            .I(N__50970));
    InMux I__8686 (
            .O(N__50985),
            .I(N__50970));
    InMux I__8685 (
            .O(N__50984),
            .I(N__50970));
    InMux I__8684 (
            .O(N__50983),
            .I(N__50970));
    InMux I__8683 (
            .O(N__50982),
            .I(N__50961));
    InMux I__8682 (
            .O(N__50981),
            .I(N__50961));
    InMux I__8681 (
            .O(N__50980),
            .I(N__50961));
    InMux I__8680 (
            .O(N__50979),
            .I(N__50961));
    LocalMux I__8679 (
            .O(N__50970),
            .I(N__50951));
    LocalMux I__8678 (
            .O(N__50961),
            .I(N__50951));
    InMux I__8677 (
            .O(N__50960),
            .I(N__50944));
    InMux I__8676 (
            .O(N__50959),
            .I(N__50944));
    InMux I__8675 (
            .O(N__50958),
            .I(N__50941));
    InMux I__8674 (
            .O(N__50957),
            .I(N__50938));
    InMux I__8673 (
            .O(N__50956),
            .I(N__50935));
    Span4Mux_s3_v I__8672 (
            .O(N__50951),
            .I(N__50931));
    InMux I__8671 (
            .O(N__50950),
            .I(N__50928));
    InMux I__8670 (
            .O(N__50949),
            .I(N__50925));
    LocalMux I__8669 (
            .O(N__50944),
            .I(N__50922));
    LocalMux I__8668 (
            .O(N__50941),
            .I(N__50915));
    LocalMux I__8667 (
            .O(N__50938),
            .I(N__50915));
    LocalMux I__8666 (
            .O(N__50935),
            .I(N__50912));
    InMux I__8665 (
            .O(N__50934),
            .I(N__50909));
    Span4Mux_h I__8664 (
            .O(N__50931),
            .I(N__50904));
    LocalMux I__8663 (
            .O(N__50928),
            .I(N__50904));
    LocalMux I__8662 (
            .O(N__50925),
            .I(N__50899));
    Span4Mux_s3_v I__8661 (
            .O(N__50922),
            .I(N__50899));
    InMux I__8660 (
            .O(N__50921),
            .I(N__50896));
    InMux I__8659 (
            .O(N__50920),
            .I(N__50893));
    Span4Mux_h I__8658 (
            .O(N__50915),
            .I(N__50886));
    Span4Mux_h I__8657 (
            .O(N__50912),
            .I(N__50886));
    LocalMux I__8656 (
            .O(N__50909),
            .I(N__50886));
    Span4Mux_h I__8655 (
            .O(N__50904),
            .I(N__50881));
    Span4Mux_h I__8654 (
            .O(N__50899),
            .I(N__50881));
    LocalMux I__8653 (
            .O(N__50896),
            .I(N__50878));
    LocalMux I__8652 (
            .O(N__50893),
            .I(\ppm_encoder_1.N_508 ));
    Odrv4 I__8651 (
            .O(N__50886),
            .I(\ppm_encoder_1.N_508 ));
    Odrv4 I__8650 (
            .O(N__50881),
            .I(\ppm_encoder_1.N_508 ));
    Odrv12 I__8649 (
            .O(N__50878),
            .I(\ppm_encoder_1.N_508 ));
    CascadeMux I__8648 (
            .O(N__50869),
            .I(N__50866));
    InMux I__8647 (
            .O(N__50866),
            .I(N__50863));
    LocalMux I__8646 (
            .O(N__50863),
            .I(N__50860));
    Span4Mux_h I__8645 (
            .O(N__50860),
            .I(N__50857));
    Span4Mux_v I__8644 (
            .O(N__50857),
            .I(N__50854));
    Odrv4 I__8643 (
            .O(N__50854),
            .I(\ppm_encoder_1.pulses2count_9_0_0_12 ));
    InMux I__8642 (
            .O(N__50851),
            .I(N__50845));
    InMux I__8641 (
            .O(N__50850),
            .I(N__50842));
    CascadeMux I__8640 (
            .O(N__50849),
            .I(N__50839));
    CascadeMux I__8639 (
            .O(N__50848),
            .I(N__50836));
    LocalMux I__8638 (
            .O(N__50845),
            .I(N__50833));
    LocalMux I__8637 (
            .O(N__50842),
            .I(N__50830));
    InMux I__8636 (
            .O(N__50839),
            .I(N__50825));
    InMux I__8635 (
            .O(N__50836),
            .I(N__50825));
    Span4Mux_v I__8634 (
            .O(N__50833),
            .I(N__50818));
    Span4Mux_v I__8633 (
            .O(N__50830),
            .I(N__50818));
    LocalMux I__8632 (
            .O(N__50825),
            .I(N__50818));
    Span4Mux_h I__8631 (
            .O(N__50818),
            .I(N__50815));
    Odrv4 I__8630 (
            .O(N__50815),
            .I(\ppm_encoder_1.init_pulsesZ0Z_12 ));
    InMux I__8629 (
            .O(N__50812),
            .I(N__50809));
    LocalMux I__8628 (
            .O(N__50809),
            .I(N__50806));
    Odrv12 I__8627 (
            .O(N__50806),
            .I(\ppm_encoder_1.pulses2count_9_0_3_12 ));
    InMux I__8626 (
            .O(N__50803),
            .I(N__50800));
    LocalMux I__8625 (
            .O(N__50800),
            .I(\uart_drone.N_144_1 ));
    CascadeMux I__8624 (
            .O(N__50797),
            .I(N__50793));
    InMux I__8623 (
            .O(N__50796),
            .I(N__50790));
    InMux I__8622 (
            .O(N__50793),
            .I(N__50787));
    LocalMux I__8621 (
            .O(N__50790),
            .I(N__50784));
    LocalMux I__8620 (
            .O(N__50787),
            .I(N__50779));
    Span4Mux_v I__8619 (
            .O(N__50784),
            .I(N__50775));
    InMux I__8618 (
            .O(N__50783),
            .I(N__50770));
    InMux I__8617 (
            .O(N__50782),
            .I(N__50770));
    Span4Mux_h I__8616 (
            .O(N__50779),
            .I(N__50767));
    InMux I__8615 (
            .O(N__50778),
            .I(N__50764));
    Odrv4 I__8614 (
            .O(N__50775),
            .I(\uart_drone.N_143 ));
    LocalMux I__8613 (
            .O(N__50770),
            .I(\uart_drone.N_143 ));
    Odrv4 I__8612 (
            .O(N__50767),
            .I(\uart_drone.N_143 ));
    LocalMux I__8611 (
            .O(N__50764),
            .I(\uart_drone.N_143 ));
    InMux I__8610 (
            .O(N__50755),
            .I(N__50752));
    LocalMux I__8609 (
            .O(N__50752),
            .I(N__50749));
    Span4Mux_h I__8608 (
            .O(N__50749),
            .I(N__50746));
    Odrv4 I__8607 (
            .O(N__50746),
            .I(\ppm_encoder_1.pulses2count_9_0_1_13 ));
    InMux I__8606 (
            .O(N__50743),
            .I(N__50740));
    LocalMux I__8605 (
            .O(N__50740),
            .I(N__50736));
    InMux I__8604 (
            .O(N__50739),
            .I(N__50733));
    Span4Mux_h I__8603 (
            .O(N__50736),
            .I(N__50730));
    LocalMux I__8602 (
            .O(N__50733),
            .I(N__50727));
    Span4Mux_h I__8601 (
            .O(N__50730),
            .I(N__50724));
    Span12Mux_s7_v I__8600 (
            .O(N__50727),
            .I(N__50721));
    Odrv4 I__8599 (
            .O(N__50724),
            .I(\ppm_encoder_1.un2_throttle_0_2_13 ));
    Odrv12 I__8598 (
            .O(N__50721),
            .I(\ppm_encoder_1.un2_throttle_0_2_13 ));
    CascadeMux I__8597 (
            .O(N__50716),
            .I(N__50713));
    InMux I__8596 (
            .O(N__50713),
            .I(N__50710));
    LocalMux I__8595 (
            .O(N__50710),
            .I(N__50707));
    Span4Mux_s1_v I__8594 (
            .O(N__50707),
            .I(N__50704));
    Odrv4 I__8593 (
            .O(N__50704),
            .I(\ppm_encoder_1.pulses2countZ0Z_13 ));
    InMux I__8592 (
            .O(N__50701),
            .I(N__50697));
    CascadeMux I__8591 (
            .O(N__50700),
            .I(N__50693));
    LocalMux I__8590 (
            .O(N__50697),
            .I(N__50690));
    CascadeMux I__8589 (
            .O(N__50696),
            .I(N__50687));
    InMux I__8588 (
            .O(N__50693),
            .I(N__50684));
    Span4Mux_h I__8587 (
            .O(N__50690),
            .I(N__50681));
    InMux I__8586 (
            .O(N__50687),
            .I(N__50678));
    LocalMux I__8585 (
            .O(N__50684),
            .I(\ppm_encoder_1.aileronZ0Z_12 ));
    Odrv4 I__8584 (
            .O(N__50681),
            .I(\ppm_encoder_1.aileronZ0Z_12 ));
    LocalMux I__8583 (
            .O(N__50678),
            .I(\ppm_encoder_1.aileronZ0Z_12 ));
    InMux I__8582 (
            .O(N__50671),
            .I(N__50668));
    LocalMux I__8581 (
            .O(N__50668),
            .I(N__50665));
    Span4Mux_s2_v I__8580 (
            .O(N__50665),
            .I(N__50662));
    Odrv4 I__8579 (
            .O(N__50662),
            .I(\ppm_encoder_1.pulses2countZ0Z_12 ));
    InMux I__8578 (
            .O(N__50659),
            .I(N__50656));
    LocalMux I__8577 (
            .O(N__50656),
            .I(N__50653));
    Span4Mux_v I__8576 (
            .O(N__50653),
            .I(N__50650));
    Span4Mux_h I__8575 (
            .O(N__50650),
            .I(N__50647));
    Odrv4 I__8574 (
            .O(N__50647),
            .I(\ppm_encoder_1.pulses2count_9_i_3_2 ));
    CascadeMux I__8573 (
            .O(N__50644),
            .I(N__50641));
    InMux I__8572 (
            .O(N__50641),
            .I(N__50638));
    LocalMux I__8571 (
            .O(N__50638),
            .I(N__50634));
    InMux I__8570 (
            .O(N__50637),
            .I(N__50631));
    Span4Mux_v I__8569 (
            .O(N__50634),
            .I(N__50627));
    LocalMux I__8568 (
            .O(N__50631),
            .I(N__50624));
    InMux I__8567 (
            .O(N__50630),
            .I(N__50621));
    Span4Mux_h I__8566 (
            .O(N__50627),
            .I(N__50616));
    Span4Mux_h I__8565 (
            .O(N__50624),
            .I(N__50616));
    LocalMux I__8564 (
            .O(N__50621),
            .I(\ppm_encoder_1.aileronZ0Z_2 ));
    Odrv4 I__8563 (
            .O(N__50616),
            .I(\ppm_encoder_1.aileronZ0Z_2 ));
    InMux I__8562 (
            .O(N__50611),
            .I(N__50608));
    LocalMux I__8561 (
            .O(N__50608),
            .I(N__50605));
    Span4Mux_h I__8560 (
            .O(N__50605),
            .I(N__50602));
    Odrv4 I__8559 (
            .O(N__50602),
            .I(\ppm_encoder_1.pulses2count_9_0_0_1_3 ));
    CascadeMux I__8558 (
            .O(N__50599),
            .I(N__50595));
    CascadeMux I__8557 (
            .O(N__50598),
            .I(N__50591));
    InMux I__8556 (
            .O(N__50595),
            .I(N__50588));
    CascadeMux I__8555 (
            .O(N__50594),
            .I(N__50585));
    InMux I__8554 (
            .O(N__50591),
            .I(N__50580));
    LocalMux I__8553 (
            .O(N__50588),
            .I(N__50577));
    InMux I__8552 (
            .O(N__50585),
            .I(N__50574));
    InMux I__8551 (
            .O(N__50584),
            .I(N__50571));
    InMux I__8550 (
            .O(N__50583),
            .I(N__50568));
    LocalMux I__8549 (
            .O(N__50580),
            .I(N__50565));
    Span4Mux_v I__8548 (
            .O(N__50577),
            .I(N__50560));
    LocalMux I__8547 (
            .O(N__50574),
            .I(N__50560));
    LocalMux I__8546 (
            .O(N__50571),
            .I(N__50556));
    LocalMux I__8545 (
            .O(N__50568),
            .I(N__50553));
    Span4Mux_h I__8544 (
            .O(N__50565),
            .I(N__50550));
    Span4Mux_h I__8543 (
            .O(N__50560),
            .I(N__50547));
    InMux I__8542 (
            .O(N__50559),
            .I(N__50544));
    Span4Mux_h I__8541 (
            .O(N__50556),
            .I(N__50539));
    Span4Mux_v I__8540 (
            .O(N__50553),
            .I(N__50539));
    Odrv4 I__8539 (
            .O(N__50550),
            .I(\ppm_encoder_1.N_514 ));
    Odrv4 I__8538 (
            .O(N__50547),
            .I(\ppm_encoder_1.N_514 ));
    LocalMux I__8537 (
            .O(N__50544),
            .I(\ppm_encoder_1.N_514 ));
    Odrv4 I__8536 (
            .O(N__50539),
            .I(\ppm_encoder_1.N_514 ));
    InMux I__8535 (
            .O(N__50530),
            .I(N__50525));
    CascadeMux I__8534 (
            .O(N__50529),
            .I(N__50522));
    CascadeMux I__8533 (
            .O(N__50528),
            .I(N__50519));
    LocalMux I__8532 (
            .O(N__50525),
            .I(N__50516));
    InMux I__8531 (
            .O(N__50522),
            .I(N__50513));
    InMux I__8530 (
            .O(N__50519),
            .I(N__50510));
    Span12Mux_h I__8529 (
            .O(N__50516),
            .I(N__50507));
    LocalMux I__8528 (
            .O(N__50513),
            .I(N__50504));
    LocalMux I__8527 (
            .O(N__50510),
            .I(\ppm_encoder_1.throttleZ0Z_3 ));
    Odrv12 I__8526 (
            .O(N__50507),
            .I(\ppm_encoder_1.throttleZ0Z_3 ));
    Odrv4 I__8525 (
            .O(N__50504),
            .I(\ppm_encoder_1.throttleZ0Z_3 ));
    CascadeMux I__8524 (
            .O(N__50497),
            .I(N__50492));
    InMux I__8523 (
            .O(N__50496),
            .I(N__50486));
    InMux I__8522 (
            .O(N__50495),
            .I(N__50486));
    InMux I__8521 (
            .O(N__50492),
            .I(N__50483));
    CascadeMux I__8520 (
            .O(N__50491),
            .I(N__50479));
    LocalMux I__8519 (
            .O(N__50486),
            .I(N__50474));
    LocalMux I__8518 (
            .O(N__50483),
            .I(N__50474));
    InMux I__8517 (
            .O(N__50482),
            .I(N__50469));
    InMux I__8516 (
            .O(N__50479),
            .I(N__50469));
    Span4Mux_h I__8515 (
            .O(N__50474),
            .I(N__50466));
    LocalMux I__8514 (
            .O(N__50469),
            .I(N__50463));
    Span4Mux_h I__8513 (
            .O(N__50466),
            .I(N__50460));
    Sp12to4 I__8512 (
            .O(N__50463),
            .I(N__50457));
    Odrv4 I__8511 (
            .O(N__50460),
            .I(\ppm_encoder_1.N_529 ));
    Odrv12 I__8510 (
            .O(N__50457),
            .I(\ppm_encoder_1.N_529 ));
    InMux I__8509 (
            .O(N__50452),
            .I(N__50448));
    InMux I__8508 (
            .O(N__50451),
            .I(N__50445));
    LocalMux I__8507 (
            .O(N__50448),
            .I(N__50440));
    LocalMux I__8506 (
            .O(N__50445),
            .I(N__50440));
    Span4Mux_h I__8505 (
            .O(N__50440),
            .I(N__50434));
    InMux I__8504 (
            .O(N__50439),
            .I(N__50427));
    InMux I__8503 (
            .O(N__50438),
            .I(N__50427));
    InMux I__8502 (
            .O(N__50437),
            .I(N__50427));
    Odrv4 I__8501 (
            .O(N__50434),
            .I(\ppm_encoder_1.N_304 ));
    LocalMux I__8500 (
            .O(N__50427),
            .I(\ppm_encoder_1.N_304 ));
    CascadeMux I__8499 (
            .O(N__50422),
            .I(\ppm_encoder_1.pulses2count_9_0_0_3_3_cascade_ ));
    InMux I__8498 (
            .O(N__50419),
            .I(N__50415));
    InMux I__8497 (
            .O(N__50418),
            .I(N__50411));
    LocalMux I__8496 (
            .O(N__50415),
            .I(N__50408));
    CascadeMux I__8495 (
            .O(N__50414),
            .I(N__50405));
    LocalMux I__8494 (
            .O(N__50411),
            .I(N__50402));
    Span4Mux_h I__8493 (
            .O(N__50408),
            .I(N__50399));
    InMux I__8492 (
            .O(N__50405),
            .I(N__50396));
    Span4Mux_v I__8491 (
            .O(N__50402),
            .I(N__50391));
    Span4Mux_v I__8490 (
            .O(N__50399),
            .I(N__50391));
    LocalMux I__8489 (
            .O(N__50396),
            .I(\ppm_encoder_1.aileronZ0Z_3 ));
    Odrv4 I__8488 (
            .O(N__50391),
            .I(\ppm_encoder_1.aileronZ0Z_3 ));
    CEMux I__8487 (
            .O(N__50386),
            .I(N__50380));
    CEMux I__8486 (
            .O(N__50385),
            .I(N__50376));
    CEMux I__8485 (
            .O(N__50384),
            .I(N__50373));
    CEMux I__8484 (
            .O(N__50383),
            .I(N__50370));
    LocalMux I__8483 (
            .O(N__50380),
            .I(N__50367));
    CEMux I__8482 (
            .O(N__50379),
            .I(N__50364));
    LocalMux I__8481 (
            .O(N__50376),
            .I(N__50361));
    LocalMux I__8480 (
            .O(N__50373),
            .I(N__50358));
    LocalMux I__8479 (
            .O(N__50370),
            .I(N__50355));
    Span4Mux_v I__8478 (
            .O(N__50367),
            .I(N__50350));
    LocalMux I__8477 (
            .O(N__50364),
            .I(N__50350));
    Span4Mux_h I__8476 (
            .O(N__50361),
            .I(N__50344));
    Span4Mux_h I__8475 (
            .O(N__50358),
            .I(N__50344));
    Span4Mux_v I__8474 (
            .O(N__50355),
            .I(N__50341));
    Span4Mux_h I__8473 (
            .O(N__50350),
            .I(N__50338));
    CEMux I__8472 (
            .O(N__50349),
            .I(N__50335));
    IoSpan4Mux I__8471 (
            .O(N__50344),
            .I(N__50332));
    Span4Mux_h I__8470 (
            .O(N__50341),
            .I(N__50327));
    Span4Mux_h I__8469 (
            .O(N__50338),
            .I(N__50327));
    LocalMux I__8468 (
            .O(N__50335),
            .I(N__50324));
    Odrv4 I__8467 (
            .O(N__50332),
            .I(\ppm_encoder_1.N_295_i_0 ));
    Odrv4 I__8466 (
            .O(N__50327),
            .I(\ppm_encoder_1.N_295_i_0 ));
    Odrv12 I__8465 (
            .O(N__50324),
            .I(\ppm_encoder_1.N_295_i_0 ));
    InMux I__8464 (
            .O(N__50317),
            .I(N__50314));
    LocalMux I__8463 (
            .O(N__50314),
            .I(\ppm_encoder_1.pulses2countZ0Z_2 ));
    CascadeMux I__8462 (
            .O(N__50311),
            .I(N__50308));
    InMux I__8461 (
            .O(N__50308),
            .I(N__50305));
    LocalMux I__8460 (
            .O(N__50305),
            .I(\ppm_encoder_1.pulses2countZ0Z_3 ));
    InMux I__8459 (
            .O(N__50302),
            .I(N__50299));
    LocalMux I__8458 (
            .O(N__50299),
            .I(N__50296));
    Span4Mux_s2_v I__8457 (
            .O(N__50296),
            .I(N__50293));
    Odrv4 I__8456 (
            .O(N__50293),
            .I(\ppm_encoder_1.counter24_0_I_9_c_RNOZ0 ));
    InMux I__8455 (
            .O(N__50290),
            .I(N__50287));
    LocalMux I__8454 (
            .O(N__50287),
            .I(\ppm_encoder_1.un1_elevator_cry_6_THRU_CO ));
    InMux I__8453 (
            .O(N__50284),
            .I(N__50281));
    LocalMux I__8452 (
            .O(N__50281),
            .I(N__50277));
    InMux I__8451 (
            .O(N__50280),
            .I(N__50274));
    Span4Mux_h I__8450 (
            .O(N__50277),
            .I(N__50271));
    LocalMux I__8449 (
            .O(N__50274),
            .I(\ppm_encoder_1.elevatorZ0Z_7 ));
    Odrv4 I__8448 (
            .O(N__50271),
            .I(\ppm_encoder_1.elevatorZ0Z_7 ));
    InMux I__8447 (
            .O(N__50266),
            .I(N__50263));
    LocalMux I__8446 (
            .O(N__50263),
            .I(N__50260));
    Odrv4 I__8445 (
            .O(N__50260),
            .I(\ppm_encoder_1.counter24_0_I_1_c_RNOZ0 ));
    InMux I__8444 (
            .O(N__50257),
            .I(N__50254));
    LocalMux I__8443 (
            .O(N__50254),
            .I(N__50251));
    Span4Mux_h I__8442 (
            .O(N__50251),
            .I(N__50248));
    Odrv4 I__8441 (
            .O(N__50248),
            .I(\ppm_encoder_1.pulses2count_9_0_3_1 ));
    CascadeMux I__8440 (
            .O(N__50245),
            .I(N__50242));
    InMux I__8439 (
            .O(N__50242),
            .I(N__50238));
    InMux I__8438 (
            .O(N__50241),
            .I(N__50235));
    LocalMux I__8437 (
            .O(N__50238),
            .I(N__50231));
    LocalMux I__8436 (
            .O(N__50235),
            .I(N__50228));
    CascadeMux I__8435 (
            .O(N__50234),
            .I(N__50225));
    Span4Mux_h I__8434 (
            .O(N__50231),
            .I(N__50222));
    Span4Mux_s2_v I__8433 (
            .O(N__50228),
            .I(N__50219));
    InMux I__8432 (
            .O(N__50225),
            .I(N__50216));
    Span4Mux_h I__8431 (
            .O(N__50222),
            .I(N__50213));
    Span4Mux_v I__8430 (
            .O(N__50219),
            .I(N__50210));
    LocalMux I__8429 (
            .O(N__50216),
            .I(\ppm_encoder_1.aileronZ0Z_1 ));
    Odrv4 I__8428 (
            .O(N__50213),
            .I(\ppm_encoder_1.aileronZ0Z_1 ));
    Odrv4 I__8427 (
            .O(N__50210),
            .I(\ppm_encoder_1.aileronZ0Z_1 ));
    InMux I__8426 (
            .O(N__50203),
            .I(N__50200));
    LocalMux I__8425 (
            .O(N__50200),
            .I(\ppm_encoder_1.pulses2countZ0Z_1 ));
    InMux I__8424 (
            .O(N__50197),
            .I(N__50194));
    LocalMux I__8423 (
            .O(N__50194),
            .I(N__50191));
    Span4Mux_h I__8422 (
            .O(N__50191),
            .I(N__50188));
    Odrv4 I__8421 (
            .O(N__50188),
            .I(\ppm_encoder_1.pulses2count_9_0_3_11 ));
    InMux I__8420 (
            .O(N__50185),
            .I(N__50181));
    CascadeMux I__8419 (
            .O(N__50184),
            .I(N__50178));
    LocalMux I__8418 (
            .O(N__50181),
            .I(N__50175));
    InMux I__8417 (
            .O(N__50178),
            .I(N__50171));
    Span4Mux_v I__8416 (
            .O(N__50175),
            .I(N__50168));
    InMux I__8415 (
            .O(N__50174),
            .I(N__50165));
    LocalMux I__8414 (
            .O(N__50171),
            .I(N__50160));
    Span4Mux_h I__8413 (
            .O(N__50168),
            .I(N__50160));
    LocalMux I__8412 (
            .O(N__50165),
            .I(N__50157));
    Odrv4 I__8411 (
            .O(N__50160),
            .I(\ppm_encoder_1.aileronZ0Z_11 ));
    Odrv4 I__8410 (
            .O(N__50157),
            .I(\ppm_encoder_1.aileronZ0Z_11 ));
    CascadeMux I__8409 (
            .O(N__50152),
            .I(N__50149));
    InMux I__8408 (
            .O(N__50149),
            .I(N__50146));
    LocalMux I__8407 (
            .O(N__50146),
            .I(\ppm_encoder_1.pulses2countZ0Z_11 ));
    InMux I__8406 (
            .O(N__50143),
            .I(N__50140));
    LocalMux I__8405 (
            .O(N__50140),
            .I(N__50137));
    Odrv4 I__8404 (
            .O(N__50137),
            .I(\ppm_encoder_1.counter24_0_I_33_c_RNOZ0 ));
    InMux I__8403 (
            .O(N__50134),
            .I(N__50131));
    LocalMux I__8402 (
            .O(N__50131),
            .I(N__50128));
    Span4Mux_h I__8401 (
            .O(N__50128),
            .I(N__50125));
    Odrv4 I__8400 (
            .O(N__50125),
            .I(\ppm_encoder_1.pulses2count_9_i_0_2_10 ));
    CascadeMux I__8399 (
            .O(N__50122),
            .I(N__50119));
    InMux I__8398 (
            .O(N__50119),
            .I(N__50114));
    CascadeMux I__8397 (
            .O(N__50118),
            .I(N__50111));
    CascadeMux I__8396 (
            .O(N__50117),
            .I(N__50107));
    LocalMux I__8395 (
            .O(N__50114),
            .I(N__50104));
    InMux I__8394 (
            .O(N__50111),
            .I(N__50101));
    InMux I__8393 (
            .O(N__50110),
            .I(N__50098));
    InMux I__8392 (
            .O(N__50107),
            .I(N__50095));
    Span4Mux_s3_v I__8391 (
            .O(N__50104),
            .I(N__50092));
    LocalMux I__8390 (
            .O(N__50101),
            .I(N__50089));
    LocalMux I__8389 (
            .O(N__50098),
            .I(N__50084));
    LocalMux I__8388 (
            .O(N__50095),
            .I(N__50084));
    Odrv4 I__8387 (
            .O(N__50092),
            .I(\ppm_encoder_1.init_pulsesZ0Z_10 ));
    Odrv4 I__8386 (
            .O(N__50089),
            .I(\ppm_encoder_1.init_pulsesZ0Z_10 ));
    Odrv4 I__8385 (
            .O(N__50084),
            .I(\ppm_encoder_1.init_pulsesZ0Z_10 ));
    InMux I__8384 (
            .O(N__50077),
            .I(N__50074));
    LocalMux I__8383 (
            .O(N__50074),
            .I(N__50071));
    Span12Mux_s5_v I__8382 (
            .O(N__50071),
            .I(N__50068));
    Odrv12 I__8381 (
            .O(N__50068),
            .I(\ppm_encoder_1.pulses2count_9_i_0_1_10 ));
    InMux I__8380 (
            .O(N__50065),
            .I(N__50062));
    LocalMux I__8379 (
            .O(N__50062),
            .I(\ppm_encoder_1.pulses2countZ0Z_10 ));
    InMux I__8378 (
            .O(N__50059),
            .I(N__50056));
    LocalMux I__8377 (
            .O(N__50056),
            .I(N__50053));
    Span4Mux_v I__8376 (
            .O(N__50053),
            .I(N__50050));
    Odrv4 I__8375 (
            .O(N__50050),
            .I(\ppm_encoder_1.pulses2count_9_0_0_0 ));
    InMux I__8374 (
            .O(N__50047),
            .I(N__50044));
    LocalMux I__8373 (
            .O(N__50044),
            .I(\ppm_encoder_1.pulses2count_9_0_2_0 ));
    InMux I__8372 (
            .O(N__50041),
            .I(N__50038));
    LocalMux I__8371 (
            .O(N__50038),
            .I(\ppm_encoder_1.pulses2countZ0Z_0 ));
    InMux I__8370 (
            .O(N__50035),
            .I(N__50032));
    LocalMux I__8369 (
            .O(N__50032),
            .I(N__50029));
    Odrv4 I__8368 (
            .O(N__50029),
            .I(\ppm_encoder_1.pulses2count_9_i_2_4 ));
    CascadeMux I__8367 (
            .O(N__50026),
            .I(N__50023));
    InMux I__8366 (
            .O(N__50023),
            .I(N__50020));
    LocalMux I__8365 (
            .O(N__50020),
            .I(\ppm_encoder_1.pulses2count_9_i_1_4 ));
    InMux I__8364 (
            .O(N__50017),
            .I(N__50014));
    LocalMux I__8363 (
            .O(N__50014),
            .I(N__50010));
    CascadeMux I__8362 (
            .O(N__50013),
            .I(N__50005));
    Span4Mux_v I__8361 (
            .O(N__50010),
            .I(N__50002));
    InMux I__8360 (
            .O(N__50009),
            .I(N__49999));
    InMux I__8359 (
            .O(N__50008),
            .I(N__49994));
    InMux I__8358 (
            .O(N__50005),
            .I(N__49994));
    Span4Mux_h I__8357 (
            .O(N__50002),
            .I(N__49989));
    LocalMux I__8356 (
            .O(N__49999),
            .I(N__49989));
    LocalMux I__8355 (
            .O(N__49994),
            .I(N__49986));
    Odrv4 I__8354 (
            .O(N__49989),
            .I(\ppm_encoder_1.init_pulsesZ0Z_4 ));
    Odrv12 I__8353 (
            .O(N__49986),
            .I(\ppm_encoder_1.init_pulsesZ0Z_4 ));
    InMux I__8352 (
            .O(N__49981),
            .I(N__49978));
    LocalMux I__8351 (
            .O(N__49978),
            .I(N__49975));
    Span4Mux_s1_v I__8350 (
            .O(N__49975),
            .I(N__49972));
    Odrv4 I__8349 (
            .O(N__49972),
            .I(\ppm_encoder_1.pulses2countZ0Z_4 ));
    CascadeMux I__8348 (
            .O(N__49969),
            .I(N__49964));
    CascadeMux I__8347 (
            .O(N__49968),
            .I(N__49961));
    InMux I__8346 (
            .O(N__49967),
            .I(N__49957));
    InMux I__8345 (
            .O(N__49964),
            .I(N__49954));
    InMux I__8344 (
            .O(N__49961),
            .I(N__49951));
    InMux I__8343 (
            .O(N__49960),
            .I(N__49948));
    LocalMux I__8342 (
            .O(N__49957),
            .I(N__49945));
    LocalMux I__8341 (
            .O(N__49954),
            .I(N__49942));
    LocalMux I__8340 (
            .O(N__49951),
            .I(N__49939));
    LocalMux I__8339 (
            .O(N__49948),
            .I(N__49936));
    Span12Mux_s2_v I__8338 (
            .O(N__49945),
            .I(N__49933));
    Span4Mux_s2_v I__8337 (
            .O(N__49942),
            .I(N__49928));
    Span4Mux_h I__8336 (
            .O(N__49939),
            .I(N__49928));
    Odrv4 I__8335 (
            .O(N__49936),
            .I(\ppm_encoder_1.init_pulsesZ0Z_5 ));
    Odrv12 I__8334 (
            .O(N__49933),
            .I(\ppm_encoder_1.init_pulsesZ0Z_5 ));
    Odrv4 I__8333 (
            .O(N__49928),
            .I(\ppm_encoder_1.init_pulsesZ0Z_5 ));
    InMux I__8332 (
            .O(N__49921),
            .I(N__49918));
    LocalMux I__8331 (
            .O(N__49918),
            .I(N__49915));
    Span4Mux_h I__8330 (
            .O(N__49915),
            .I(N__49912));
    Span4Mux_h I__8329 (
            .O(N__49912),
            .I(N__49908));
    InMux I__8328 (
            .O(N__49911),
            .I(N__49905));
    Odrv4 I__8327 (
            .O(N__49908),
            .I(\ppm_encoder_1.N_307 ));
    LocalMux I__8326 (
            .O(N__49905),
            .I(\ppm_encoder_1.N_307 ));
    CascadeMux I__8325 (
            .O(N__49900),
            .I(N__49897));
    InMux I__8324 (
            .O(N__49897),
            .I(N__49894));
    LocalMux I__8323 (
            .O(N__49894),
            .I(N__49891));
    Span4Mux_s1_v I__8322 (
            .O(N__49891),
            .I(N__49888));
    Odrv4 I__8321 (
            .O(N__49888),
            .I(\ppm_encoder_1.pulses2countZ0Z_5 ));
    InMux I__8320 (
            .O(N__49885),
            .I(N__49882));
    LocalMux I__8319 (
            .O(N__49882),
            .I(\ppm_encoder_1.pulses2countZ0Z_8 ));
    CascadeMux I__8318 (
            .O(N__49879),
            .I(N__49876));
    InMux I__8317 (
            .O(N__49876),
            .I(N__49873));
    LocalMux I__8316 (
            .O(N__49873),
            .I(N__49870));
    Span4Mux_h I__8315 (
            .O(N__49870),
            .I(N__49867));
    Span4Mux_h I__8314 (
            .O(N__49867),
            .I(N__49864));
    Odrv4 I__8313 (
            .O(N__49864),
            .I(\ppm_encoder_1.pulses2countZ0Z_9 ));
    InMux I__8312 (
            .O(N__49861),
            .I(N__49858));
    LocalMux I__8311 (
            .O(N__49858),
            .I(\ppm_encoder_1.counter24_0_I_27_c_RNOZ0 ));
    InMux I__8310 (
            .O(N__49855),
            .I(N__49851));
    InMux I__8309 (
            .O(N__49854),
            .I(N__49848));
    LocalMux I__8308 (
            .O(N__49851),
            .I(N__49845));
    LocalMux I__8307 (
            .O(N__49848),
            .I(N__49842));
    Span12Mux_s11_h I__8306 (
            .O(N__49845),
            .I(N__49839));
    Span12Mux_s2_v I__8305 (
            .O(N__49842),
            .I(N__49836));
    Odrv12 I__8304 (
            .O(N__49839),
            .I(\ppm_encoder_1.counter24_0_I_57_c_RNIJMMDZ0 ));
    Odrv12 I__8303 (
            .O(N__49836),
            .I(\ppm_encoder_1.counter24_0_I_57_c_RNIJMMDZ0 ));
    CascadeMux I__8302 (
            .O(N__49831),
            .I(\ppm_encoder_1.counter24_0_I_57_c_RNIJMMDZ0_cascade_ ));
    InMux I__8301 (
            .O(N__49828),
            .I(N__49825));
    LocalMux I__8300 (
            .O(N__49825),
            .I(\ppm_encoder_1.N_500 ));
    IoInMux I__8299 (
            .O(N__49822),
            .I(N__49819));
    LocalMux I__8298 (
            .O(N__49819),
            .I(N__49816));
    IoSpan4Mux I__8297 (
            .O(N__49816),
            .I(N__49813));
    Span4Mux_s2_v I__8296 (
            .O(N__49813),
            .I(N__49810));
    Span4Mux_v I__8295 (
            .O(N__49810),
            .I(N__49806));
    InMux I__8294 (
            .O(N__49809),
            .I(N__49803));
    Odrv4 I__8293 (
            .O(N__49806),
            .I(ppm_output_c));
    LocalMux I__8292 (
            .O(N__49803),
            .I(ppm_output_c));
    CascadeMux I__8291 (
            .O(N__49798),
            .I(N__49794));
    CascadeMux I__8290 (
            .O(N__49797),
            .I(N__49791));
    InMux I__8289 (
            .O(N__49794),
            .I(N__49786));
    InMux I__8288 (
            .O(N__49791),
            .I(N__49786));
    LocalMux I__8287 (
            .O(N__49786),
            .I(\ppm_encoder_1.N_486_9 ));
    InMux I__8286 (
            .O(N__49783),
            .I(N__49776));
    InMux I__8285 (
            .O(N__49782),
            .I(N__49771));
    InMux I__8284 (
            .O(N__49781),
            .I(N__49771));
    InMux I__8283 (
            .O(N__49780),
            .I(N__49766));
    InMux I__8282 (
            .O(N__49779),
            .I(N__49766));
    LocalMux I__8281 (
            .O(N__49776),
            .I(N__49761));
    LocalMux I__8280 (
            .O(N__49771),
            .I(N__49758));
    LocalMux I__8279 (
            .O(N__49766),
            .I(N__49755));
    InMux I__8278 (
            .O(N__49765),
            .I(N__49750));
    InMux I__8277 (
            .O(N__49764),
            .I(N__49750));
    Odrv4 I__8276 (
            .O(N__49761),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_1 ));
    Odrv12 I__8275 (
            .O(N__49758),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_1 ));
    Odrv4 I__8274 (
            .O(N__49755),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_1 ));
    LocalMux I__8273 (
            .O(N__49750),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_1 ));
    InMux I__8272 (
            .O(N__49741),
            .I(N__49737));
    InMux I__8271 (
            .O(N__49740),
            .I(N__49734));
    LocalMux I__8270 (
            .O(N__49737),
            .I(N__49730));
    LocalMux I__8269 (
            .O(N__49734),
            .I(N__49727));
    InMux I__8268 (
            .O(N__49733),
            .I(N__49724));
    Span4Mux_h I__8267 (
            .O(N__49730),
            .I(N__49721));
    Span4Mux_v I__8266 (
            .O(N__49727),
            .I(N__49716));
    LocalMux I__8265 (
            .O(N__49724),
            .I(N__49716));
    Span4Mux_h I__8264 (
            .O(N__49721),
            .I(N__49713));
    Span4Mux_h I__8263 (
            .O(N__49716),
            .I(N__49710));
    Odrv4 I__8262 (
            .O(N__49713),
            .I(\ppm_encoder_1.N_486 ));
    Odrv4 I__8261 (
            .O(N__49710),
            .I(\ppm_encoder_1.N_486 ));
    CascadeMux I__8260 (
            .O(N__49705),
            .I(\ppm_encoder_1.N_486_cascade_ ));
    InMux I__8259 (
            .O(N__49702),
            .I(N__49693));
    CascadeMux I__8258 (
            .O(N__49701),
            .I(N__49687));
    InMux I__8257 (
            .O(N__49700),
            .I(N__49680));
    InMux I__8256 (
            .O(N__49699),
            .I(N__49680));
    InMux I__8255 (
            .O(N__49698),
            .I(N__49680));
    InMux I__8254 (
            .O(N__49697),
            .I(N__49677));
    CascadeMux I__8253 (
            .O(N__49696),
            .I(N__49673));
    LocalMux I__8252 (
            .O(N__49693),
            .I(N__49669));
    InMux I__8251 (
            .O(N__49692),
            .I(N__49664));
    InMux I__8250 (
            .O(N__49691),
            .I(N__49664));
    InMux I__8249 (
            .O(N__49690),
            .I(N__49659));
    InMux I__8248 (
            .O(N__49687),
            .I(N__49659));
    LocalMux I__8247 (
            .O(N__49680),
            .I(N__49652));
    LocalMux I__8246 (
            .O(N__49677),
            .I(N__49652));
    CascadeMux I__8245 (
            .O(N__49676),
            .I(N__49649));
    InMux I__8244 (
            .O(N__49673),
            .I(N__49636));
    InMux I__8243 (
            .O(N__49672),
            .I(N__49636));
    Span4Mux_s1_v I__8242 (
            .O(N__49669),
            .I(N__49629));
    LocalMux I__8241 (
            .O(N__49664),
            .I(N__49629));
    LocalMux I__8240 (
            .O(N__49659),
            .I(N__49629));
    InMux I__8239 (
            .O(N__49658),
            .I(N__49624));
    InMux I__8238 (
            .O(N__49657),
            .I(N__49624));
    Span4Mux_s3_v I__8237 (
            .O(N__49652),
            .I(N__49620));
    InMux I__8236 (
            .O(N__49649),
            .I(N__49615));
    InMux I__8235 (
            .O(N__49648),
            .I(N__49615));
    InMux I__8234 (
            .O(N__49647),
            .I(N__49608));
    InMux I__8233 (
            .O(N__49646),
            .I(N__49608));
    InMux I__8232 (
            .O(N__49645),
            .I(N__49608));
    InMux I__8231 (
            .O(N__49644),
            .I(N__49599));
    InMux I__8230 (
            .O(N__49643),
            .I(N__49599));
    InMux I__8229 (
            .O(N__49642),
            .I(N__49599));
    InMux I__8228 (
            .O(N__49641),
            .I(N__49599));
    LocalMux I__8227 (
            .O(N__49636),
            .I(N__49592));
    Span4Mux_v I__8226 (
            .O(N__49629),
            .I(N__49592));
    LocalMux I__8225 (
            .O(N__49624),
            .I(N__49592));
    InMux I__8224 (
            .O(N__49623),
            .I(N__49589));
    Span4Mux_h I__8223 (
            .O(N__49620),
            .I(N__49586));
    LocalMux I__8222 (
            .O(N__49615),
            .I(N__49583));
    LocalMux I__8221 (
            .O(N__49608),
            .I(N__49580));
    LocalMux I__8220 (
            .O(N__49599),
            .I(N__49575));
    Span4Mux_h I__8219 (
            .O(N__49592),
            .I(N__49575));
    LocalMux I__8218 (
            .O(N__49589),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ));
    Odrv4 I__8217 (
            .O(N__49586),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ));
    Odrv4 I__8216 (
            .O(N__49583),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ));
    Odrv4 I__8215 (
            .O(N__49580),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ));
    Odrv4 I__8214 (
            .O(N__49575),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ));
    InMux I__8213 (
            .O(N__49564),
            .I(N__49555));
    InMux I__8212 (
            .O(N__49563),
            .I(N__49555));
    InMux I__8211 (
            .O(N__49562),
            .I(N__49555));
    LocalMux I__8210 (
            .O(N__49555),
            .I(\ppm_encoder_1.counter24_0_N_2_THRU_CO ));
    InMux I__8209 (
            .O(N__49552),
            .I(N__49546));
    InMux I__8208 (
            .O(N__49551),
            .I(N__49539));
    InMux I__8207 (
            .O(N__49550),
            .I(N__49539));
    InMux I__8206 (
            .O(N__49549),
            .I(N__49539));
    LocalMux I__8205 (
            .O(N__49546),
            .I(N__49534));
    LocalMux I__8204 (
            .O(N__49539),
            .I(N__49534));
    Span4Mux_h I__8203 (
            .O(N__49534),
            .I(N__49528));
    InMux I__8202 (
            .O(N__49533),
            .I(N__49523));
    InMux I__8201 (
            .O(N__49532),
            .I(N__49523));
    CascadeMux I__8200 (
            .O(N__49531),
            .I(N__49520));
    Span4Mux_h I__8199 (
            .O(N__49528),
            .I(N__49517));
    LocalMux I__8198 (
            .O(N__49523),
            .I(N__49514));
    InMux I__8197 (
            .O(N__49520),
            .I(N__49511));
    Odrv4 I__8196 (
            .O(N__49517),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_0 ));
    Odrv4 I__8195 (
            .O(N__49514),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_0 ));
    LocalMux I__8194 (
            .O(N__49511),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_0 ));
    CascadeMux I__8193 (
            .O(N__49504),
            .I(N__49496));
    CascadeMux I__8192 (
            .O(N__49503),
            .I(N__49492));
    CascadeMux I__8191 (
            .O(N__49502),
            .I(N__49489));
    CascadeMux I__8190 (
            .O(N__49501),
            .I(N__49486));
    CascadeMux I__8189 (
            .O(N__49500),
            .I(N__49483));
    InMux I__8188 (
            .O(N__49499),
            .I(N__49477));
    InMux I__8187 (
            .O(N__49496),
            .I(N__49472));
    InMux I__8186 (
            .O(N__49495),
            .I(N__49472));
    InMux I__8185 (
            .O(N__49492),
            .I(N__49465));
    InMux I__8184 (
            .O(N__49489),
            .I(N__49465));
    InMux I__8183 (
            .O(N__49486),
            .I(N__49465));
    InMux I__8182 (
            .O(N__49483),
            .I(N__49456));
    InMux I__8181 (
            .O(N__49482),
            .I(N__49456));
    InMux I__8180 (
            .O(N__49481),
            .I(N__49456));
    InMux I__8179 (
            .O(N__49480),
            .I(N__49456));
    LocalMux I__8178 (
            .O(N__49477),
            .I(N__49448));
    LocalMux I__8177 (
            .O(N__49472),
            .I(N__49445));
    LocalMux I__8176 (
            .O(N__49465),
            .I(N__49437));
    LocalMux I__8175 (
            .O(N__49456),
            .I(N__49437));
    InMux I__8174 (
            .O(N__49455),
            .I(N__49426));
    InMux I__8173 (
            .O(N__49454),
            .I(N__49426));
    InMux I__8172 (
            .O(N__49453),
            .I(N__49426));
    InMux I__8171 (
            .O(N__49452),
            .I(N__49426));
    InMux I__8170 (
            .O(N__49451),
            .I(N__49426));
    Span4Mux_s2_v I__8169 (
            .O(N__49448),
            .I(N__49421));
    Span4Mux_s2_v I__8168 (
            .O(N__49445),
            .I(N__49421));
    InMux I__8167 (
            .O(N__49444),
            .I(N__49416));
    InMux I__8166 (
            .O(N__49443),
            .I(N__49416));
    InMux I__8165 (
            .O(N__49442),
            .I(N__49413));
    Span4Mux_h I__8164 (
            .O(N__49437),
            .I(N__49410));
    LocalMux I__8163 (
            .O(N__49426),
            .I(N__49405));
    Span4Mux_h I__8162 (
            .O(N__49421),
            .I(N__49405));
    LocalMux I__8161 (
            .O(N__49416),
            .I(\ppm_encoder_1.N_374 ));
    LocalMux I__8160 (
            .O(N__49413),
            .I(\ppm_encoder_1.N_374 ));
    Odrv4 I__8159 (
            .O(N__49410),
            .I(\ppm_encoder_1.N_374 ));
    Odrv4 I__8158 (
            .O(N__49405),
            .I(\ppm_encoder_1.N_374 ));
    CascadeMux I__8157 (
            .O(N__49396),
            .I(N__49391));
    CascadeMux I__8156 (
            .O(N__49395),
            .I(N__49387));
    InMux I__8155 (
            .O(N__49394),
            .I(N__49378));
    InMux I__8154 (
            .O(N__49391),
            .I(N__49371));
    InMux I__8153 (
            .O(N__49390),
            .I(N__49371));
    InMux I__8152 (
            .O(N__49387),
            .I(N__49371));
    CascadeMux I__8151 (
            .O(N__49386),
            .I(N__49366));
    CascadeMux I__8150 (
            .O(N__49385),
            .I(N__49363));
    CascadeMux I__8149 (
            .O(N__49384),
            .I(N__49360));
    CascadeMux I__8148 (
            .O(N__49383),
            .I(N__49357));
    CascadeMux I__8147 (
            .O(N__49382),
            .I(N__49354));
    CascadeMux I__8146 (
            .O(N__49381),
            .I(N__49351));
    LocalMux I__8145 (
            .O(N__49378),
            .I(N__49348));
    LocalMux I__8144 (
            .O(N__49371),
            .I(N__49345));
    InMux I__8143 (
            .O(N__49370),
            .I(N__49340));
    InMux I__8142 (
            .O(N__49369),
            .I(N__49340));
    InMux I__8141 (
            .O(N__49366),
            .I(N__49333));
    InMux I__8140 (
            .O(N__49363),
            .I(N__49333));
    InMux I__8139 (
            .O(N__49360),
            .I(N__49333));
    InMux I__8138 (
            .O(N__49357),
            .I(N__49328));
    InMux I__8137 (
            .O(N__49354),
            .I(N__49328));
    InMux I__8136 (
            .O(N__49351),
            .I(N__49325));
    Span4Mux_v I__8135 (
            .O(N__49348),
            .I(N__49322));
    Span4Mux_s3_v I__8134 (
            .O(N__49345),
            .I(N__49319));
    LocalMux I__8133 (
            .O(N__49340),
            .I(N__49314));
    LocalMux I__8132 (
            .O(N__49333),
            .I(N__49314));
    LocalMux I__8131 (
            .O(N__49328),
            .I(N__49309));
    LocalMux I__8130 (
            .O(N__49325),
            .I(N__49309));
    Span4Mux_h I__8129 (
            .O(N__49322),
            .I(N__49300));
    Span4Mux_h I__8128 (
            .O(N__49319),
            .I(N__49293));
    Span4Mux_s3_v I__8127 (
            .O(N__49314),
            .I(N__49293));
    Span4Mux_h I__8126 (
            .O(N__49309),
            .I(N__49293));
    InMux I__8125 (
            .O(N__49308),
            .I(N__49280));
    InMux I__8124 (
            .O(N__49307),
            .I(N__49280));
    InMux I__8123 (
            .O(N__49306),
            .I(N__49280));
    InMux I__8122 (
            .O(N__49305),
            .I(N__49280));
    InMux I__8121 (
            .O(N__49304),
            .I(N__49280));
    InMux I__8120 (
            .O(N__49303),
            .I(N__49280));
    Odrv4 I__8119 (
            .O(N__49300),
            .I(\ppm_encoder_1.N_298 ));
    Odrv4 I__8118 (
            .O(N__49293),
            .I(\ppm_encoder_1.N_298 ));
    LocalMux I__8117 (
            .O(N__49280),
            .I(\ppm_encoder_1.N_298 ));
    InMux I__8116 (
            .O(N__49273),
            .I(N__49270));
    LocalMux I__8115 (
            .O(N__49270),
            .I(N__49267));
    Span4Mux_h I__8114 (
            .O(N__49267),
            .I(N__49264));
    Odrv4 I__8113 (
            .O(N__49264),
            .I(\ppm_encoder_1.un1_init_pulses_11_0 ));
    CascadeMux I__8112 (
            .O(N__49261),
            .I(\ppm_encoder_1.N_374_cascade_ ));
    InMux I__8111 (
            .O(N__49258),
            .I(N__49255));
    LocalMux I__8110 (
            .O(N__49255),
            .I(N__49252));
    Span4Mux_v I__8109 (
            .O(N__49252),
            .I(N__49249));
    Odrv4 I__8108 (
            .O(N__49249),
            .I(\ppm_encoder_1.un1_init_pulses_10_0 ));
    CascadeMux I__8107 (
            .O(N__49246),
            .I(N__49242));
    InMux I__8106 (
            .O(N__49245),
            .I(N__49239));
    InMux I__8105 (
            .O(N__49242),
            .I(N__49236));
    LocalMux I__8104 (
            .O(N__49239),
            .I(N__49233));
    LocalMux I__8103 (
            .O(N__49236),
            .I(N__49230));
    Span4Mux_h I__8102 (
            .O(N__49233),
            .I(N__49227));
    Span4Mux_h I__8101 (
            .O(N__49230),
            .I(N__49224));
    Odrv4 I__8100 (
            .O(N__49227),
            .I(\ppm_encoder_1.init_pulsesZ0Z_0 ));
    Odrv4 I__8099 (
            .O(N__49224),
            .I(\ppm_encoder_1.init_pulsesZ0Z_0 ));
    CascadeMux I__8098 (
            .O(N__49219),
            .I(N__49214));
    InMux I__8097 (
            .O(N__49218),
            .I(N__49211));
    InMux I__8096 (
            .O(N__49217),
            .I(N__49206));
    InMux I__8095 (
            .O(N__49214),
            .I(N__49206));
    LocalMux I__8094 (
            .O(N__49211),
            .I(N__49203));
    LocalMux I__8093 (
            .O(N__49206),
            .I(N__49200));
    Span4Mux_h I__8092 (
            .O(N__49203),
            .I(N__49197));
    Span4Mux_h I__8091 (
            .O(N__49200),
            .I(N__49194));
    Odrv4 I__8090 (
            .O(N__49197),
            .I(\ppm_encoder_1.init_pulsesZ0Z_16 ));
    Odrv4 I__8089 (
            .O(N__49194),
            .I(\ppm_encoder_1.init_pulsesZ0Z_16 ));
    InMux I__8088 (
            .O(N__49189),
            .I(N__49186));
    LocalMux I__8087 (
            .O(N__49186),
            .I(\ppm_encoder_1.pulses2countZ0Z_16 ));
    InMux I__8086 (
            .O(N__49183),
            .I(N__49180));
    LocalMux I__8085 (
            .O(N__49180),
            .I(N__49176));
    CascadeMux I__8084 (
            .O(N__49179),
            .I(N__49173));
    Span4Mux_s3_v I__8083 (
            .O(N__49176),
            .I(N__49169));
    InMux I__8082 (
            .O(N__49173),
            .I(N__49166));
    InMux I__8081 (
            .O(N__49172),
            .I(N__49163));
    Odrv4 I__8080 (
            .O(N__49169),
            .I(\ppm_encoder_1.init_pulsesZ0Z_17 ));
    LocalMux I__8079 (
            .O(N__49166),
            .I(\ppm_encoder_1.init_pulsesZ0Z_17 ));
    LocalMux I__8078 (
            .O(N__49163),
            .I(\ppm_encoder_1.init_pulsesZ0Z_17 ));
    CascadeMux I__8077 (
            .O(N__49156),
            .I(N__49153));
    InMux I__8076 (
            .O(N__49153),
            .I(N__49150));
    LocalMux I__8075 (
            .O(N__49150),
            .I(\ppm_encoder_1.pulses2countZ0Z_17 ));
    InMux I__8074 (
            .O(N__49147),
            .I(N__49144));
    LocalMux I__8073 (
            .O(N__49144),
            .I(\ppm_encoder_1.counter24_0_I_21_c_RNOZ0 ));
    CascadeMux I__8072 (
            .O(N__49141),
            .I(N__49138));
    InMux I__8071 (
            .O(N__49138),
            .I(N__49133));
    CascadeMux I__8070 (
            .O(N__49137),
            .I(N__49130));
    CascadeMux I__8069 (
            .O(N__49136),
            .I(N__49127));
    LocalMux I__8068 (
            .O(N__49133),
            .I(N__49123));
    InMux I__8067 (
            .O(N__49130),
            .I(N__49118));
    InMux I__8066 (
            .O(N__49127),
            .I(N__49118));
    InMux I__8065 (
            .O(N__49126),
            .I(N__49115));
    Span4Mux_s2_v I__8064 (
            .O(N__49123),
            .I(N__49112));
    LocalMux I__8063 (
            .O(N__49118),
            .I(N__49109));
    LocalMux I__8062 (
            .O(N__49115),
            .I(N__49106));
    Odrv4 I__8061 (
            .O(N__49112),
            .I(\ppm_encoder_1.init_pulsesZ0Z_6 ));
    Odrv4 I__8060 (
            .O(N__49109),
            .I(\ppm_encoder_1.init_pulsesZ0Z_6 ));
    Odrv12 I__8059 (
            .O(N__49106),
            .I(\ppm_encoder_1.init_pulsesZ0Z_6 ));
    InMux I__8058 (
            .O(N__49099),
            .I(N__49096));
    LocalMux I__8057 (
            .O(N__49096),
            .I(N__49093));
    Span4Mux_h I__8056 (
            .O(N__49093),
            .I(N__49089));
    InMux I__8055 (
            .O(N__49092),
            .I(N__49086));
    Odrv4 I__8054 (
            .O(N__49089),
            .I(\ppm_encoder_1.N_306 ));
    LocalMux I__8053 (
            .O(N__49086),
            .I(\ppm_encoder_1.N_306 ));
    InMux I__8052 (
            .O(N__49081),
            .I(N__49078));
    LocalMux I__8051 (
            .O(N__49078),
            .I(\ppm_encoder_1.pulses2countZ0Z_6 ));
    CascadeMux I__8050 (
            .O(N__49075),
            .I(N__49072));
    InMux I__8049 (
            .O(N__49072),
            .I(N__49068));
    CascadeMux I__8048 (
            .O(N__49071),
            .I(N__49065));
    LocalMux I__8047 (
            .O(N__49068),
            .I(N__49060));
    InMux I__8046 (
            .O(N__49065),
            .I(N__49055));
    InMux I__8045 (
            .O(N__49064),
            .I(N__49055));
    InMux I__8044 (
            .O(N__49063),
            .I(N__49052));
    Span4Mux_h I__8043 (
            .O(N__49060),
            .I(N__49047));
    LocalMux I__8042 (
            .O(N__49055),
            .I(N__49047));
    LocalMux I__8041 (
            .O(N__49052),
            .I(\ppm_encoder_1.init_pulsesZ0Z_7 ));
    Odrv4 I__8040 (
            .O(N__49047),
            .I(\ppm_encoder_1.init_pulsesZ0Z_7 ));
    InMux I__8039 (
            .O(N__49042),
            .I(N__49039));
    LocalMux I__8038 (
            .O(N__49039),
            .I(N__49036));
    Span4Mux_v I__8037 (
            .O(N__49036),
            .I(N__49032));
    InMux I__8036 (
            .O(N__49035),
            .I(N__49029));
    Odrv4 I__8035 (
            .O(N__49032),
            .I(\ppm_encoder_1.N_310 ));
    LocalMux I__8034 (
            .O(N__49029),
            .I(\ppm_encoder_1.N_310 ));
    CascadeMux I__8033 (
            .O(N__49024),
            .I(N__49021));
    InMux I__8032 (
            .O(N__49021),
            .I(N__49018));
    LocalMux I__8031 (
            .O(N__49018),
            .I(\ppm_encoder_1.pulses2countZ0Z_7 ));
    InMux I__8030 (
            .O(N__49015),
            .I(N__49012));
    LocalMux I__8029 (
            .O(N__49012),
            .I(N__49009));
    Span4Mux_h I__8028 (
            .O(N__49009),
            .I(N__49006));
    Span4Mux_s1_v I__8027 (
            .O(N__49006),
            .I(N__49001));
    InMux I__8026 (
            .O(N__49005),
            .I(N__48998));
    InMux I__8025 (
            .O(N__49004),
            .I(N__48995));
    Odrv4 I__8024 (
            .O(N__49001),
            .I(\ppm_encoder_1.init_pulsesZ0Z_18 ));
    LocalMux I__8023 (
            .O(N__48998),
            .I(\ppm_encoder_1.init_pulsesZ0Z_18 ));
    LocalMux I__8022 (
            .O(N__48995),
            .I(\ppm_encoder_1.init_pulsesZ0Z_18 ));
    InMux I__8021 (
            .O(N__48988),
            .I(N__48985));
    LocalMux I__8020 (
            .O(N__48985),
            .I(\ppm_encoder_1.pulses2countZ0Z_18 ));
    InMux I__8019 (
            .O(N__48982),
            .I(N__48979));
    LocalMux I__8018 (
            .O(N__48979),
            .I(\ppm_encoder_1.counter24_0_I_57_c_RNOZ0 ));
    InMux I__8017 (
            .O(N__48976),
            .I(N__48973));
    LocalMux I__8016 (
            .O(N__48973),
            .I(N__48970));
    Span4Mux_s1_v I__8015 (
            .O(N__48970),
            .I(N__48967));
    Odrv4 I__8014 (
            .O(N__48967),
            .I(\ppm_encoder_1.pulses2count_9_i_2_8 ));
    CascadeMux I__8013 (
            .O(N__48964),
            .I(N__48958));
    InMux I__8012 (
            .O(N__48963),
            .I(N__48955));
    InMux I__8011 (
            .O(N__48962),
            .I(N__48952));
    InMux I__8010 (
            .O(N__48961),
            .I(N__48949));
    InMux I__8009 (
            .O(N__48958),
            .I(N__48946));
    LocalMux I__8008 (
            .O(N__48955),
            .I(N__48943));
    LocalMux I__8007 (
            .O(N__48952),
            .I(N__48940));
    LocalMux I__8006 (
            .O(N__48949),
            .I(N__48937));
    LocalMux I__8005 (
            .O(N__48946),
            .I(N__48934));
    Span4Mux_h I__8004 (
            .O(N__48943),
            .I(N__48929));
    Span4Mux_h I__8003 (
            .O(N__48940),
            .I(N__48929));
    Span4Mux_h I__8002 (
            .O(N__48937),
            .I(N__48926));
    Span4Mux_h I__8001 (
            .O(N__48934),
            .I(N__48921));
    Span4Mux_h I__8000 (
            .O(N__48929),
            .I(N__48921));
    Odrv4 I__7999 (
            .O(N__48926),
            .I(\ppm_encoder_1.init_pulsesZ0Z_8 ));
    Odrv4 I__7998 (
            .O(N__48921),
            .I(\ppm_encoder_1.init_pulsesZ0Z_8 ));
    InMux I__7997 (
            .O(N__48916),
            .I(N__48913));
    LocalMux I__7996 (
            .O(N__48913),
            .I(N__48910));
    Span4Mux_s3_v I__7995 (
            .O(N__48910),
            .I(N__48907));
    Span4Mux_v I__7994 (
            .O(N__48907),
            .I(N__48904));
    Odrv4 I__7993 (
            .O(N__48904),
            .I(\ppm_encoder_1.pulses2count_9_i_1_8 ));
    InMux I__7992 (
            .O(N__48901),
            .I(N__48898));
    LocalMux I__7991 (
            .O(N__48898),
            .I(\dron_frame_decoder_1.state_ns_i_a2_0_1_0 ));
    CascadeMux I__7990 (
            .O(N__48895),
            .I(\dron_frame_decoder_1.N_224_cascade_ ));
    CascadeMux I__7989 (
            .O(N__48892),
            .I(\dron_frame_decoder_1.state_ns_i_a2_1_1Z0Z_0_cascade_ ));
    InMux I__7988 (
            .O(N__48889),
            .I(N__48886));
    LocalMux I__7987 (
            .O(N__48886),
            .I(\dron_frame_decoder_1.N_220 ));
    InMux I__7986 (
            .O(N__48883),
            .I(N__48880));
    LocalMux I__7985 (
            .O(N__48880),
            .I(N__48877));
    Odrv4 I__7984 (
            .O(N__48877),
            .I(\dron_frame_decoder_1.N_224 ));
    CascadeMux I__7983 (
            .O(N__48874),
            .I(\dron_frame_decoder_1.N_220_cascade_ ));
    InMux I__7982 (
            .O(N__48871),
            .I(N__48866));
    InMux I__7981 (
            .O(N__48870),
            .I(N__48861));
    InMux I__7980 (
            .O(N__48869),
            .I(N__48861));
    LocalMux I__7979 (
            .O(N__48866),
            .I(\dron_frame_decoder_1.stateZ0Z_1 ));
    LocalMux I__7978 (
            .O(N__48861),
            .I(\dron_frame_decoder_1.stateZ0Z_1 ));
    CascadeMux I__7977 (
            .O(N__48856),
            .I(N__48853));
    InMux I__7976 (
            .O(N__48853),
            .I(N__48850));
    LocalMux I__7975 (
            .O(N__48850),
            .I(\dron_frame_decoder_1.N_200 ));
    InMux I__7974 (
            .O(N__48847),
            .I(N__48844));
    LocalMux I__7973 (
            .O(N__48844),
            .I(\dron_frame_decoder_1.N_198 ));
    CascadeMux I__7972 (
            .O(N__48841),
            .I(N__48838));
    InMux I__7971 (
            .O(N__48838),
            .I(N__48830));
    InMux I__7970 (
            .O(N__48837),
            .I(N__48830));
    InMux I__7969 (
            .O(N__48836),
            .I(N__48825));
    InMux I__7968 (
            .O(N__48835),
            .I(N__48825));
    LocalMux I__7967 (
            .O(N__48830),
            .I(\dron_frame_decoder_1.stateZ0Z_0 ));
    LocalMux I__7966 (
            .O(N__48825),
            .I(\dron_frame_decoder_1.stateZ0Z_0 ));
    InMux I__7965 (
            .O(N__48820),
            .I(N__48817));
    LocalMux I__7964 (
            .O(N__48817),
            .I(N__48814));
    Odrv4 I__7963 (
            .O(N__48814),
            .I(\dron_frame_decoder_1.state_ns_i_a2_0_2_0 ));
    InMux I__7962 (
            .O(N__48811),
            .I(N__48808));
    LocalMux I__7961 (
            .O(N__48808),
            .I(\ppm_encoder_1.counter24_0_I_15_c_RNOZ0 ));
    InMux I__7960 (
            .O(N__48805),
            .I(N__48801));
    CascadeMux I__7959 (
            .O(N__48804),
            .I(N__48796));
    LocalMux I__7958 (
            .O(N__48801),
            .I(N__48793));
    InMux I__7957 (
            .O(N__48800),
            .I(N__48790));
    InMux I__7956 (
            .O(N__48799),
            .I(N__48785));
    InMux I__7955 (
            .O(N__48796),
            .I(N__48785));
    Span4Mux_h I__7954 (
            .O(N__48793),
            .I(N__48780));
    LocalMux I__7953 (
            .O(N__48790),
            .I(N__48780));
    LocalMux I__7952 (
            .O(N__48785),
            .I(N__48777));
    Odrv4 I__7951 (
            .O(N__48780),
            .I(\ppm_encoder_1.init_pulsesZ0Z_15 ));
    Odrv4 I__7950 (
            .O(N__48777),
            .I(\ppm_encoder_1.init_pulsesZ0Z_15 ));
    InMux I__7949 (
            .O(N__48772),
            .I(N__48767));
    CascadeMux I__7948 (
            .O(N__48771),
            .I(N__48764));
    CascadeMux I__7947 (
            .O(N__48770),
            .I(N__48760));
    LocalMux I__7946 (
            .O(N__48767),
            .I(N__48757));
    InMux I__7945 (
            .O(N__48764),
            .I(N__48754));
    InMux I__7944 (
            .O(N__48763),
            .I(N__48749));
    InMux I__7943 (
            .O(N__48760),
            .I(N__48749));
    Span4Mux_h I__7942 (
            .O(N__48757),
            .I(N__48744));
    LocalMux I__7941 (
            .O(N__48754),
            .I(N__48744));
    LocalMux I__7940 (
            .O(N__48749),
            .I(N__48741));
    Odrv4 I__7939 (
            .O(N__48744),
            .I(\ppm_encoder_1.init_pulsesZ0Z_14 ));
    Odrv4 I__7938 (
            .O(N__48741),
            .I(\ppm_encoder_1.init_pulsesZ0Z_14 ));
    InMux I__7937 (
            .O(N__48736),
            .I(N__48733));
    LocalMux I__7936 (
            .O(N__48733),
            .I(N__48730));
    Span4Mux_s1_v I__7935 (
            .O(N__48730),
            .I(N__48727));
    Span4Mux_v I__7934 (
            .O(N__48727),
            .I(N__48723));
    InMux I__7933 (
            .O(N__48726),
            .I(N__48720));
    Odrv4 I__7932 (
            .O(N__48723),
            .I(\ppm_encoder_1.N_309 ));
    LocalMux I__7931 (
            .O(N__48720),
            .I(\ppm_encoder_1.N_309 ));
    InMux I__7930 (
            .O(N__48715),
            .I(N__48712));
    LocalMux I__7929 (
            .O(N__48712),
            .I(\dron_frame_decoder_1.drone_altitude_9 ));
    CEMux I__7928 (
            .O(N__48709),
            .I(N__48705));
    CEMux I__7927 (
            .O(N__48708),
            .I(N__48702));
    LocalMux I__7926 (
            .O(N__48705),
            .I(N__48696));
    LocalMux I__7925 (
            .O(N__48702),
            .I(N__48696));
    CEMux I__7924 (
            .O(N__48701),
            .I(N__48693));
    Span4Mux_v I__7923 (
            .O(N__48696),
            .I(N__48686));
    LocalMux I__7922 (
            .O(N__48693),
            .I(N__48686));
    CEMux I__7921 (
            .O(N__48692),
            .I(N__48683));
    CEMux I__7920 (
            .O(N__48691),
            .I(N__48680));
    Span4Mux_s3_h I__7919 (
            .O(N__48686),
            .I(N__48677));
    LocalMux I__7918 (
            .O(N__48683),
            .I(N__48674));
    LocalMux I__7917 (
            .O(N__48680),
            .I(N__48671));
    Span4Mux_h I__7916 (
            .O(N__48677),
            .I(N__48666));
    Span4Mux_h I__7915 (
            .O(N__48674),
            .I(N__48666));
    Span4Mux_v I__7914 (
            .O(N__48671),
            .I(N__48663));
    Span4Mux_h I__7913 (
            .O(N__48666),
            .I(N__48660));
    Span4Mux_h I__7912 (
            .O(N__48663),
            .I(N__48657));
    Odrv4 I__7911 (
            .O(N__48660),
            .I(\Commands_frame_decoder.state_RNIF38SZ0Z_6 ));
    Odrv4 I__7910 (
            .O(N__48657),
            .I(\Commands_frame_decoder.state_RNIF38SZ0Z_6 ));
    InMux I__7909 (
            .O(N__48652),
            .I(N__48649));
    LocalMux I__7908 (
            .O(N__48649),
            .I(\dron_frame_decoder_1.state_RNI3T3K1Z0Z_7 ));
    InMux I__7907 (
            .O(N__48646),
            .I(N__48643));
    LocalMux I__7906 (
            .O(N__48643),
            .I(\dron_frame_decoder_1.drone_altitude_10 ));
    InMux I__7905 (
            .O(N__48640),
            .I(N__48637));
    LocalMux I__7904 (
            .O(N__48637),
            .I(N__48634));
    Span4Mux_h I__7903 (
            .O(N__48634),
            .I(N__48631));
    Span4Mux_h I__7902 (
            .O(N__48631),
            .I(N__48628));
    Odrv4 I__7901 (
            .O(N__48628),
            .I(drone_altitude_i_10));
    InMux I__7900 (
            .O(N__48625),
            .I(N__48621));
    InMux I__7899 (
            .O(N__48624),
            .I(N__48618));
    LocalMux I__7898 (
            .O(N__48621),
            .I(N__48614));
    LocalMux I__7897 (
            .O(N__48618),
            .I(N__48611));
    InMux I__7896 (
            .O(N__48617),
            .I(N__48608));
    Span4Mux_v I__7895 (
            .O(N__48614),
            .I(N__48603));
    Span4Mux_h I__7894 (
            .O(N__48611),
            .I(N__48603));
    LocalMux I__7893 (
            .O(N__48608),
            .I(\Commands_frame_decoder.stateZ0Z_13 ));
    Odrv4 I__7892 (
            .O(N__48603),
            .I(\Commands_frame_decoder.stateZ0Z_13 ));
    InMux I__7891 (
            .O(N__48598),
            .I(N__48594));
    InMux I__7890 (
            .O(N__48597),
            .I(N__48591));
    LocalMux I__7889 (
            .O(N__48594),
            .I(N__48588));
    LocalMux I__7888 (
            .O(N__48591),
            .I(\Commands_frame_decoder.stateZ0Z_12 ));
    Odrv12 I__7887 (
            .O(N__48588),
            .I(\Commands_frame_decoder.stateZ0Z_12 ));
    InMux I__7886 (
            .O(N__48583),
            .I(N__48580));
    LocalMux I__7885 (
            .O(N__48580),
            .I(N__48577));
    Span4Mux_h I__7884 (
            .O(N__48577),
            .I(N__48574));
    Odrv4 I__7883 (
            .O(N__48574),
            .I(\Commands_frame_decoder.source_xy_ki_1_sqmuxa ));
    CascadeMux I__7882 (
            .O(N__48571),
            .I(\Commands_frame_decoder.source_xy_ki_1_sqmuxa_cascade_ ));
    InMux I__7881 (
            .O(N__48568),
            .I(N__48565));
    LocalMux I__7880 (
            .O(N__48565),
            .I(\dron_frame_decoder_1.N_230_5 ));
    CascadeMux I__7879 (
            .O(N__48562),
            .I(\dron_frame_decoder_1.N_230_5_cascade_ ));
    CascadeMux I__7878 (
            .O(N__48559),
            .I(N__48545));
    InMux I__7877 (
            .O(N__48558),
            .I(N__48540));
    InMux I__7876 (
            .O(N__48557),
            .I(N__48535));
    InMux I__7875 (
            .O(N__48556),
            .I(N__48535));
    InMux I__7874 (
            .O(N__48555),
            .I(N__48526));
    InMux I__7873 (
            .O(N__48554),
            .I(N__48526));
    InMux I__7872 (
            .O(N__48553),
            .I(N__48526));
    InMux I__7871 (
            .O(N__48552),
            .I(N__48526));
    InMux I__7870 (
            .O(N__48551),
            .I(N__48523));
    InMux I__7869 (
            .O(N__48550),
            .I(N__48518));
    InMux I__7868 (
            .O(N__48549),
            .I(N__48518));
    InMux I__7867 (
            .O(N__48548),
            .I(N__48515));
    InMux I__7866 (
            .O(N__48545),
            .I(N__48508));
    InMux I__7865 (
            .O(N__48544),
            .I(N__48508));
    InMux I__7864 (
            .O(N__48543),
            .I(N__48508));
    LocalMux I__7863 (
            .O(N__48540),
            .I(N__48503));
    LocalMux I__7862 (
            .O(N__48535),
            .I(N__48503));
    LocalMux I__7861 (
            .O(N__48526),
            .I(uart_drone_data_rdy));
    LocalMux I__7860 (
            .O(N__48523),
            .I(uart_drone_data_rdy));
    LocalMux I__7859 (
            .O(N__48518),
            .I(uart_drone_data_rdy));
    LocalMux I__7858 (
            .O(N__48515),
            .I(uart_drone_data_rdy));
    LocalMux I__7857 (
            .O(N__48508),
            .I(uart_drone_data_rdy));
    Odrv12 I__7856 (
            .O(N__48503),
            .I(uart_drone_data_rdy));
    InMux I__7855 (
            .O(N__48490),
            .I(N__48487));
    LocalMux I__7854 (
            .O(N__48487),
            .I(\dron_frame_decoder_1.drone_altitude_5 ));
    InMux I__7853 (
            .O(N__48484),
            .I(N__48481));
    LocalMux I__7852 (
            .O(N__48481),
            .I(\dron_frame_decoder_1.drone_altitude_6 ));
    InMux I__7851 (
            .O(N__48478),
            .I(N__48475));
    LocalMux I__7850 (
            .O(N__48475),
            .I(\dron_frame_decoder_1.drone_altitude_7 ));
    CEMux I__7849 (
            .O(N__48472),
            .I(N__48469));
    LocalMux I__7848 (
            .O(N__48469),
            .I(N__48466));
    Span4Mux_v I__7847 (
            .O(N__48466),
            .I(N__48463));
    Odrv4 I__7846 (
            .O(N__48463),
            .I(\dron_frame_decoder_1.N_740_0 ));
    InMux I__7845 (
            .O(N__48460),
            .I(N__48457));
    LocalMux I__7844 (
            .O(N__48457),
            .I(N__48454));
    Odrv4 I__7843 (
            .O(N__48454),
            .I(drone_altitude_12));
    InMux I__7842 (
            .O(N__48451),
            .I(N__48448));
    LocalMux I__7841 (
            .O(N__48448),
            .I(N__48445));
    Odrv12 I__7840 (
            .O(N__48445),
            .I(drone_altitude_15));
    InMux I__7839 (
            .O(N__48442),
            .I(N__48439));
    LocalMux I__7838 (
            .O(N__48439),
            .I(N__48436));
    Span4Mux_h I__7837 (
            .O(N__48436),
            .I(N__48433));
    Odrv4 I__7836 (
            .O(N__48433),
            .I(\dron_frame_decoder_1.drone_altitude_8 ));
    InMux I__7835 (
            .O(N__48430),
            .I(N__48427));
    LocalMux I__7834 (
            .O(N__48427),
            .I(N__48424));
    Span4Mux_h I__7833 (
            .O(N__48424),
            .I(N__48421));
    Span4Mux_h I__7832 (
            .O(N__48421),
            .I(N__48418));
    Odrv4 I__7831 (
            .O(N__48418),
            .I(\pid_alt.error_axbZ0Z_1 ));
    InMux I__7830 (
            .O(N__48415),
            .I(N__48412));
    LocalMux I__7829 (
            .O(N__48412),
            .I(N__48409));
    Span4Mux_h I__7828 (
            .O(N__48409),
            .I(N__48406));
    Span4Mux_h I__7827 (
            .O(N__48406),
            .I(N__48403));
    Odrv4 I__7826 (
            .O(N__48403),
            .I(\pid_alt.error_axbZ0Z_12 ));
    InMux I__7825 (
            .O(N__48400),
            .I(N__48397));
    LocalMux I__7824 (
            .O(N__48397),
            .I(N__48393));
    InMux I__7823 (
            .O(N__48396),
            .I(N__48390));
    Span4Mux_v I__7822 (
            .O(N__48393),
            .I(N__48385));
    LocalMux I__7821 (
            .O(N__48390),
            .I(N__48385));
    Span4Mux_v I__7820 (
            .O(N__48385),
            .I(N__48381));
    InMux I__7819 (
            .O(N__48384),
            .I(N__48378));
    Sp12to4 I__7818 (
            .O(N__48381),
            .I(N__48375));
    LocalMux I__7817 (
            .O(N__48378),
            .I(N__48372));
    Span12Mux_s10_h I__7816 (
            .O(N__48375),
            .I(N__48366));
    Span12Mux_s10_h I__7815 (
            .O(N__48372),
            .I(N__48366));
    InMux I__7814 (
            .O(N__48371),
            .I(N__48363));
    Odrv12 I__7813 (
            .O(N__48366),
            .I(drone_altitude_0));
    LocalMux I__7812 (
            .O(N__48363),
            .I(drone_altitude_0));
    InMux I__7811 (
            .O(N__48358),
            .I(N__48355));
    LocalMux I__7810 (
            .O(N__48355),
            .I(drone_altitude_1));
    InMux I__7809 (
            .O(N__48352),
            .I(N__48349));
    LocalMux I__7808 (
            .O(N__48349),
            .I(\dron_frame_decoder_1.drone_altitude_4 ));
    InMux I__7807 (
            .O(N__48346),
            .I(N__48343));
    LocalMux I__7806 (
            .O(N__48343),
            .I(N__48340));
    Span4Mux_v I__7805 (
            .O(N__48340),
            .I(N__48337));
    Odrv4 I__7804 (
            .O(N__48337),
            .I(\Commands_frame_decoder.WDT8lt14_0 ));
    CascadeMux I__7803 (
            .O(N__48334),
            .I(N__48331));
    InMux I__7802 (
            .O(N__48331),
            .I(N__48328));
    LocalMux I__7801 (
            .O(N__48328),
            .I(N__48322));
    CascadeMux I__7800 (
            .O(N__48327),
            .I(N__48318));
    InMux I__7799 (
            .O(N__48326),
            .I(N__48315));
    InMux I__7798 (
            .O(N__48325),
            .I(N__48312));
    Span4Mux_h I__7797 (
            .O(N__48322),
            .I(N__48309));
    InMux I__7796 (
            .O(N__48321),
            .I(N__48304));
    InMux I__7795 (
            .O(N__48318),
            .I(N__48304));
    LocalMux I__7794 (
            .O(N__48315),
            .I(\Commands_frame_decoder.WDTZ0Z_15 ));
    LocalMux I__7793 (
            .O(N__48312),
            .I(\Commands_frame_decoder.WDTZ0Z_15 ));
    Odrv4 I__7792 (
            .O(N__48309),
            .I(\Commands_frame_decoder.WDTZ0Z_15 ));
    LocalMux I__7791 (
            .O(N__48304),
            .I(\Commands_frame_decoder.WDTZ0Z_15 ));
    InMux I__7790 (
            .O(N__48295),
            .I(N__48292));
    LocalMux I__7789 (
            .O(N__48292),
            .I(N__48288));
    InMux I__7788 (
            .O(N__48291),
            .I(N__48283));
    Span4Mux_h I__7787 (
            .O(N__48288),
            .I(N__48280));
    InMux I__7786 (
            .O(N__48287),
            .I(N__48277));
    InMux I__7785 (
            .O(N__48286),
            .I(N__48274));
    LocalMux I__7784 (
            .O(N__48283),
            .I(\Commands_frame_decoder.WDTZ0Z_14 ));
    Odrv4 I__7783 (
            .O(N__48280),
            .I(\Commands_frame_decoder.WDTZ0Z_14 ));
    LocalMux I__7782 (
            .O(N__48277),
            .I(\Commands_frame_decoder.WDTZ0Z_14 ));
    LocalMux I__7781 (
            .O(N__48274),
            .I(\Commands_frame_decoder.WDTZ0Z_14 ));
    InMux I__7780 (
            .O(N__48265),
            .I(N__48262));
    LocalMux I__7779 (
            .O(N__48262),
            .I(N__48258));
    InMux I__7778 (
            .O(N__48261),
            .I(N__48255));
    Span4Mux_h I__7777 (
            .O(N__48258),
            .I(N__48251));
    LocalMux I__7776 (
            .O(N__48255),
            .I(N__48248));
    InMux I__7775 (
            .O(N__48254),
            .I(N__48245));
    Span4Mux_v I__7774 (
            .O(N__48251),
            .I(N__48242));
    Span12Mux_v I__7773 (
            .O(N__48248),
            .I(N__48239));
    LocalMux I__7772 (
            .O(N__48245),
            .I(\Commands_frame_decoder.stateZ0Z_10 ));
    Odrv4 I__7771 (
            .O(N__48242),
            .I(\Commands_frame_decoder.stateZ0Z_10 ));
    Odrv12 I__7770 (
            .O(N__48239),
            .I(\Commands_frame_decoder.stateZ0Z_10 ));
    CascadeMux I__7769 (
            .O(N__48232),
            .I(\Commands_frame_decoder.N_403_cascade_ ));
    CascadeMux I__7768 (
            .O(N__48229),
            .I(N__48226));
    InMux I__7767 (
            .O(N__48226),
            .I(N__48220));
    InMux I__7766 (
            .O(N__48225),
            .I(N__48220));
    LocalMux I__7765 (
            .O(N__48220),
            .I(\Commands_frame_decoder.stateZ0Z_8 ));
    InMux I__7764 (
            .O(N__48217),
            .I(N__48213));
    InMux I__7763 (
            .O(N__48216),
            .I(N__48210));
    LocalMux I__7762 (
            .O(N__48213),
            .I(\Commands_frame_decoder.stateZ0Z_9 ));
    LocalMux I__7761 (
            .O(N__48210),
            .I(\Commands_frame_decoder.stateZ0Z_9 ));
    InMux I__7760 (
            .O(N__48205),
            .I(N__48202));
    LocalMux I__7759 (
            .O(N__48202),
            .I(N__48199));
    Span4Mux_v I__7758 (
            .O(N__48199),
            .I(N__48196));
    Span4Mux_v I__7757 (
            .O(N__48196),
            .I(N__48191));
    InMux I__7756 (
            .O(N__48195),
            .I(N__48186));
    InMux I__7755 (
            .O(N__48194),
            .I(N__48186));
    Odrv4 I__7754 (
            .O(N__48191),
            .I(\uart_drone.data_rdyc_1 ));
    LocalMux I__7753 (
            .O(N__48186),
            .I(\uart_drone.data_rdyc_1 ));
    CascadeMux I__7752 (
            .O(N__48181),
            .I(N__48178));
    InMux I__7751 (
            .O(N__48178),
            .I(N__48175));
    LocalMux I__7750 (
            .O(N__48175),
            .I(N__48172));
    Odrv4 I__7749 (
            .O(N__48172),
            .I(\uart_drone.timer_Count_RNO_0_0_4 ));
    InMux I__7748 (
            .O(N__48169),
            .I(N__48166));
    LocalMux I__7747 (
            .O(N__48166),
            .I(\uart_drone.timer_Count_RNO_0_0_3 ));
    InMux I__7746 (
            .O(N__48163),
            .I(N__48160));
    LocalMux I__7745 (
            .O(N__48160),
            .I(N__48157));
    Span4Mux_v I__7744 (
            .O(N__48157),
            .I(N__48154));
    Span4Mux_v I__7743 (
            .O(N__48154),
            .I(N__48151));
    Span4Mux_h I__7742 (
            .O(N__48151),
            .I(N__48148));
    Odrv4 I__7741 (
            .O(N__48148),
            .I(\uart_drone_sync.aux_1__0__0_0 ));
    InMux I__7740 (
            .O(N__48145),
            .I(N__48142));
    LocalMux I__7739 (
            .O(N__48142),
            .I(N__48139));
    Span4Mux_v I__7738 (
            .O(N__48139),
            .I(N__48136));
    Span4Mux_h I__7737 (
            .O(N__48136),
            .I(N__48133));
    Odrv4 I__7736 (
            .O(N__48133),
            .I(\uart_pc_sync.aux_1__0_Z0Z_0 ));
    InMux I__7735 (
            .O(N__48130),
            .I(N__48127));
    LocalMux I__7734 (
            .O(N__48127),
            .I(\uart_pc_sync.aux_2__0_Z0Z_0 ));
    InMux I__7733 (
            .O(N__48124),
            .I(N__48121));
    LocalMux I__7732 (
            .O(N__48121),
            .I(\uart_pc_sync.aux_3__0_Z0Z_0 ));
    IoInMux I__7731 (
            .O(N__48118),
            .I(N__48115));
    LocalMux I__7730 (
            .O(N__48115),
            .I(N__48112));
    Span4Mux_s3_v I__7729 (
            .O(N__48112),
            .I(N__48109));
    Span4Mux_v I__7728 (
            .O(N__48109),
            .I(N__48104));
    InMux I__7727 (
            .O(N__48108),
            .I(N__48100));
    InMux I__7726 (
            .O(N__48107),
            .I(N__48097));
    Sp12to4 I__7725 (
            .O(N__48104),
            .I(N__48094));
    CascadeMux I__7724 (
            .O(N__48103),
            .I(N__48091));
    LocalMux I__7723 (
            .O(N__48100),
            .I(N__48088));
    LocalMux I__7722 (
            .O(N__48097),
            .I(N__48085));
    Span12Mux_h I__7721 (
            .O(N__48094),
            .I(N__48082));
    InMux I__7720 (
            .O(N__48091),
            .I(N__48079));
    Span4Mux_h I__7719 (
            .O(N__48088),
            .I(N__48074));
    Span4Mux_h I__7718 (
            .O(N__48085),
            .I(N__48074));
    Odrv12 I__7717 (
            .O(N__48082),
            .I(debug_CH3_20A_c));
    LocalMux I__7716 (
            .O(N__48079),
            .I(debug_CH3_20A_c));
    Odrv4 I__7715 (
            .O(N__48074),
            .I(debug_CH3_20A_c));
    CEMux I__7714 (
            .O(N__48067),
            .I(N__48064));
    LocalMux I__7713 (
            .O(N__48064),
            .I(N__48059));
    CEMux I__7712 (
            .O(N__48063),
            .I(N__48056));
    CEMux I__7711 (
            .O(N__48062),
            .I(N__48053));
    Span4Mux_v I__7710 (
            .O(N__48059),
            .I(N__48050));
    LocalMux I__7709 (
            .O(N__48056),
            .I(N__48047));
    LocalMux I__7708 (
            .O(N__48053),
            .I(N__48044));
    Span4Mux_h I__7707 (
            .O(N__48050),
            .I(N__48039));
    Span4Mux_v I__7706 (
            .O(N__48047),
            .I(N__48039));
    Span4Mux_h I__7705 (
            .O(N__48044),
            .I(N__48036));
    Odrv4 I__7704 (
            .O(N__48039),
            .I(\scaler_4.debug_CH3_20A_c_0 ));
    Odrv4 I__7703 (
            .O(N__48036),
            .I(\scaler_4.debug_CH3_20A_c_0 ));
    CEMux I__7702 (
            .O(N__48031),
            .I(N__48028));
    LocalMux I__7701 (
            .O(N__48028),
            .I(N__48025));
    Odrv4 I__7700 (
            .O(N__48025),
            .I(\Commands_frame_decoder.state_RNIG48SZ0Z_7 ));
    InMux I__7699 (
            .O(N__48022),
            .I(N__48019));
    LocalMux I__7698 (
            .O(N__48019),
            .I(N__48016));
    Span4Mux_h I__7697 (
            .O(N__48016),
            .I(N__48013));
    Odrv4 I__7696 (
            .O(N__48013),
            .I(\ppm_encoder_1.un1_aileron_cry_10_THRU_CO ));
    InMux I__7695 (
            .O(N__48010),
            .I(\ppm_encoder_1.un1_aileron_cry_10 ));
    InMux I__7694 (
            .O(N__48007),
            .I(N__48004));
    LocalMux I__7693 (
            .O(N__48004),
            .I(N__48001));
    Span4Mux_h I__7692 (
            .O(N__48001),
            .I(N__47998));
    Odrv4 I__7691 (
            .O(N__47998),
            .I(\ppm_encoder_1.un1_aileron_cry_11_THRU_CO ));
    InMux I__7690 (
            .O(N__47995),
            .I(\ppm_encoder_1.un1_aileron_cry_11 ));
    InMux I__7689 (
            .O(N__47992),
            .I(\ppm_encoder_1.un1_aileron_cry_12 ));
    InMux I__7688 (
            .O(N__47989),
            .I(\ppm_encoder_1.un1_aileron_cry_13 ));
    CEMux I__7687 (
            .O(N__47986),
            .I(N__47981));
    CEMux I__7686 (
            .O(N__47985),
            .I(N__47977));
    CEMux I__7685 (
            .O(N__47984),
            .I(N__47974));
    LocalMux I__7684 (
            .O(N__47981),
            .I(N__47970));
    CEMux I__7683 (
            .O(N__47980),
            .I(N__47967));
    LocalMux I__7682 (
            .O(N__47977),
            .I(N__47964));
    LocalMux I__7681 (
            .O(N__47974),
            .I(N__47961));
    CEMux I__7680 (
            .O(N__47973),
            .I(N__47958));
    Span4Mux_v I__7679 (
            .O(N__47970),
            .I(N__47955));
    LocalMux I__7678 (
            .O(N__47967),
            .I(N__47951));
    Span4Mux_v I__7677 (
            .O(N__47964),
            .I(N__47948));
    Span4Mux_v I__7676 (
            .O(N__47961),
            .I(N__47945));
    LocalMux I__7675 (
            .O(N__47958),
            .I(N__47942));
    Sp12to4 I__7674 (
            .O(N__47955),
            .I(N__47939));
    CEMux I__7673 (
            .O(N__47954),
            .I(N__47936));
    Span4Mux_h I__7672 (
            .O(N__47951),
            .I(N__47933));
    Span4Mux_v I__7671 (
            .O(N__47948),
            .I(N__47928));
    Span4Mux_h I__7670 (
            .O(N__47945),
            .I(N__47928));
    Span12Mux_v I__7669 (
            .O(N__47942),
            .I(N__47923));
    Span12Mux_s10_h I__7668 (
            .O(N__47939),
            .I(N__47923));
    LocalMux I__7667 (
            .O(N__47936),
            .I(\ppm_encoder_1.pid_altitude_dv_0 ));
    Odrv4 I__7666 (
            .O(N__47933),
            .I(\ppm_encoder_1.pid_altitude_dv_0 ));
    Odrv4 I__7665 (
            .O(N__47928),
            .I(\ppm_encoder_1.pid_altitude_dv_0 ));
    Odrv12 I__7664 (
            .O(N__47923),
            .I(\ppm_encoder_1.pid_altitude_dv_0 ));
    InMux I__7663 (
            .O(N__47914),
            .I(N__47909));
    CascadeMux I__7662 (
            .O(N__47913),
            .I(N__47905));
    InMux I__7661 (
            .O(N__47912),
            .I(N__47902));
    LocalMux I__7660 (
            .O(N__47909),
            .I(N__47899));
    InMux I__7659 (
            .O(N__47908),
            .I(N__47894));
    InMux I__7658 (
            .O(N__47905),
            .I(N__47894));
    LocalMux I__7657 (
            .O(N__47902),
            .I(\uart_drone.timer_CountZ0Z_0 ));
    Odrv12 I__7656 (
            .O(N__47899),
            .I(\uart_drone.timer_CountZ0Z_0 ));
    LocalMux I__7655 (
            .O(N__47894),
            .I(\uart_drone.timer_CountZ0Z_0 ));
    CascadeMux I__7654 (
            .O(N__47887),
            .I(N__47882));
    InMux I__7653 (
            .O(N__47886),
            .I(N__47879));
    InMux I__7652 (
            .O(N__47885),
            .I(N__47874));
    InMux I__7651 (
            .O(N__47882),
            .I(N__47874));
    LocalMux I__7650 (
            .O(N__47879),
            .I(\uart_drone.timer_CountZ1Z_2 ));
    LocalMux I__7649 (
            .O(N__47874),
            .I(\uart_drone.timer_CountZ1Z_2 ));
    InMux I__7648 (
            .O(N__47869),
            .I(N__47866));
    LocalMux I__7647 (
            .O(N__47866),
            .I(\uart_drone.timer_Count_RNO_0_0_2 ));
    InMux I__7646 (
            .O(N__47863),
            .I(\uart_drone.un4_timer_Count_1_cry_1 ));
    InMux I__7645 (
            .O(N__47860),
            .I(\uart_drone.un4_timer_Count_1_cry_2 ));
    InMux I__7644 (
            .O(N__47857),
            .I(\uart_drone.un4_timer_Count_1_cry_3 ));
    InMux I__7643 (
            .O(N__47854),
            .I(N__47851));
    LocalMux I__7642 (
            .O(N__47851),
            .I(N__47848));
    Span4Mux_v I__7641 (
            .O(N__47848),
            .I(N__47845));
    Odrv4 I__7640 (
            .O(N__47845),
            .I(\ppm_encoder_1.un1_aileron_cry_2_THRU_CO ));
    InMux I__7639 (
            .O(N__47842),
            .I(\ppm_encoder_1.un1_aileron_cry_2 ));
    InMux I__7638 (
            .O(N__47839),
            .I(N__47836));
    LocalMux I__7637 (
            .O(N__47836),
            .I(\ppm_encoder_1.un1_aileron_cry_3_THRU_CO ));
    InMux I__7636 (
            .O(N__47833),
            .I(\ppm_encoder_1.un1_aileron_cry_3 ));
    InMux I__7635 (
            .O(N__47830),
            .I(N__47827));
    LocalMux I__7634 (
            .O(N__47827),
            .I(N__47824));
    Span4Mux_v I__7633 (
            .O(N__47824),
            .I(N__47821));
    Sp12to4 I__7632 (
            .O(N__47821),
            .I(N__47818));
    Odrv12 I__7631 (
            .O(N__47818),
            .I(\ppm_encoder_1.un1_aileron_cry_4_THRU_CO ));
    InMux I__7630 (
            .O(N__47815),
            .I(\ppm_encoder_1.un1_aileron_cry_4 ));
    InMux I__7629 (
            .O(N__47812),
            .I(N__47809));
    LocalMux I__7628 (
            .O(N__47809),
            .I(\ppm_encoder_1.un1_aileron_cry_5_THRU_CO ));
    InMux I__7627 (
            .O(N__47806),
            .I(\ppm_encoder_1.un1_aileron_cry_5 ));
    InMux I__7626 (
            .O(N__47803),
            .I(N__47800));
    LocalMux I__7625 (
            .O(N__47800),
            .I(N__47797));
    Span4Mux_h I__7624 (
            .O(N__47797),
            .I(N__47794));
    Odrv4 I__7623 (
            .O(N__47794),
            .I(\ppm_encoder_1.un1_aileron_cry_6_THRU_CO ));
    InMux I__7622 (
            .O(N__47791),
            .I(\ppm_encoder_1.un1_aileron_cry_6 ));
    InMux I__7621 (
            .O(N__47788),
            .I(N__47785));
    LocalMux I__7620 (
            .O(N__47785),
            .I(N__47782));
    Span12Mux_s10_h I__7619 (
            .O(N__47782),
            .I(N__47779));
    Odrv12 I__7618 (
            .O(N__47779),
            .I(\ppm_encoder_1.un1_aileron_cry_7_THRU_CO ));
    InMux I__7617 (
            .O(N__47776),
            .I(bfn_10_11_0_));
    InMux I__7616 (
            .O(N__47773),
            .I(N__47770));
    LocalMux I__7615 (
            .O(N__47770),
            .I(N__47767));
    Span4Mux_h I__7614 (
            .O(N__47767),
            .I(N__47764));
    Odrv4 I__7613 (
            .O(N__47764),
            .I(\ppm_encoder_1.un1_aileron_cry_8_THRU_CO ));
    InMux I__7612 (
            .O(N__47761),
            .I(\ppm_encoder_1.un1_aileron_cry_8 ));
    InMux I__7611 (
            .O(N__47758),
            .I(N__47755));
    LocalMux I__7610 (
            .O(N__47755),
            .I(N__47752));
    Span4Mux_h I__7609 (
            .O(N__47752),
            .I(N__47749));
    Odrv4 I__7608 (
            .O(N__47749),
            .I(\ppm_encoder_1.un1_aileron_cry_9_THRU_CO ));
    InMux I__7607 (
            .O(N__47746),
            .I(\ppm_encoder_1.un1_aileron_cry_9 ));
    CascadeMux I__7606 (
            .O(N__47743),
            .I(\uart_drone.N_152_cascade_ ));
    InMux I__7605 (
            .O(N__47740),
            .I(N__47734));
    InMux I__7604 (
            .O(N__47739),
            .I(N__47734));
    LocalMux I__7603 (
            .O(N__47734),
            .I(\uart_drone.un1_state_7_0 ));
    InMux I__7602 (
            .O(N__47731),
            .I(N__47728));
    LocalMux I__7601 (
            .O(N__47728),
            .I(\uart_drone.CO0 ));
    InMux I__7600 (
            .O(N__47725),
            .I(N__47722));
    LocalMux I__7599 (
            .O(N__47722),
            .I(N__47717));
    InMux I__7598 (
            .O(N__47721),
            .I(N__47714));
    InMux I__7597 (
            .O(N__47720),
            .I(N__47711));
    Span4Mux_v I__7596 (
            .O(N__47717),
            .I(N__47706));
    LocalMux I__7595 (
            .O(N__47714),
            .I(N__47706));
    LocalMux I__7594 (
            .O(N__47711),
            .I(\ppm_encoder_1.throttleZ0Z_12 ));
    Odrv4 I__7593 (
            .O(N__47706),
            .I(\ppm_encoder_1.throttleZ0Z_12 ));
    InMux I__7592 (
            .O(N__47701),
            .I(N__47698));
    LocalMux I__7591 (
            .O(N__47698),
            .I(N__47695));
    Span4Mux_h I__7590 (
            .O(N__47695),
            .I(N__47692));
    Odrv4 I__7589 (
            .O(N__47692),
            .I(\ppm_encoder_1.un1_aileron_cry_0_THRU_CO ));
    InMux I__7588 (
            .O(N__47689),
            .I(\ppm_encoder_1.un1_aileron_cry_0 ));
    InMux I__7587 (
            .O(N__47686),
            .I(N__47683));
    LocalMux I__7586 (
            .O(N__47683),
            .I(N__47680));
    Span4Mux_h I__7585 (
            .O(N__47680),
            .I(N__47677));
    Odrv4 I__7584 (
            .O(N__47677),
            .I(\ppm_encoder_1.un1_aileron_cry_1_THRU_CO ));
    InMux I__7583 (
            .O(N__47674),
            .I(\ppm_encoder_1.un1_aileron_cry_1 ));
    InMux I__7582 (
            .O(N__47671),
            .I(N__47668));
    LocalMux I__7581 (
            .O(N__47668),
            .I(N__47665));
    Span4Mux_s3_v I__7580 (
            .O(N__47665),
            .I(N__47662));
    Odrv4 I__7579 (
            .O(N__47662),
            .I(\ppm_encoder_1.un1_elevator_cry_5_THRU_CO ));
    InMux I__7578 (
            .O(N__47659),
            .I(\ppm_encoder_1.un1_elevator_cry_5 ));
    InMux I__7577 (
            .O(N__47656),
            .I(\ppm_encoder_1.un1_elevator_cry_6 ));
    InMux I__7576 (
            .O(N__47653),
            .I(N__47650));
    LocalMux I__7575 (
            .O(N__47650),
            .I(N__47647));
    Span4Mux_v I__7574 (
            .O(N__47647),
            .I(N__47644));
    Span4Mux_h I__7573 (
            .O(N__47644),
            .I(N__47641));
    Odrv4 I__7572 (
            .O(N__47641),
            .I(\ppm_encoder_1.un1_elevator_cry_7_THRU_CO ));
    InMux I__7571 (
            .O(N__47638),
            .I(bfn_10_8_0_));
    InMux I__7570 (
            .O(N__47635),
            .I(N__47632));
    LocalMux I__7569 (
            .O(N__47632),
            .I(\ppm_encoder_1.un1_elevator_cry_8_THRU_CO ));
    InMux I__7568 (
            .O(N__47629),
            .I(\ppm_encoder_1.un1_elevator_cry_8 ));
    InMux I__7567 (
            .O(N__47626),
            .I(N__47623));
    LocalMux I__7566 (
            .O(N__47623),
            .I(N__47620));
    Odrv4 I__7565 (
            .O(N__47620),
            .I(\ppm_encoder_1.un1_elevator_cry_9_THRU_CO ));
    InMux I__7564 (
            .O(N__47617),
            .I(\ppm_encoder_1.un1_elevator_cry_9 ));
    InMux I__7563 (
            .O(N__47614),
            .I(N__47611));
    LocalMux I__7562 (
            .O(N__47611),
            .I(N__47608));
    Odrv12 I__7561 (
            .O(N__47608),
            .I(\ppm_encoder_1.un1_elevator_cry_10_THRU_CO ));
    InMux I__7560 (
            .O(N__47605),
            .I(\ppm_encoder_1.un1_elevator_cry_10 ));
    InMux I__7559 (
            .O(N__47602),
            .I(N__47599));
    LocalMux I__7558 (
            .O(N__47599),
            .I(N__47596));
    Span4Mux_v I__7557 (
            .O(N__47596),
            .I(N__47593));
    Span4Mux_h I__7556 (
            .O(N__47593),
            .I(N__47590));
    Odrv4 I__7555 (
            .O(N__47590),
            .I(\ppm_encoder_1.un1_elevator_cry_11_THRU_CO ));
    InMux I__7554 (
            .O(N__47587),
            .I(\ppm_encoder_1.un1_elevator_cry_11 ));
    InMux I__7553 (
            .O(N__47584),
            .I(N__47581));
    LocalMux I__7552 (
            .O(N__47581),
            .I(N__47578));
    Span4Mux_v I__7551 (
            .O(N__47578),
            .I(N__47575));
    Odrv4 I__7550 (
            .O(N__47575),
            .I(\ppm_encoder_1.un1_elevator_cry_12_THRU_CO ));
    InMux I__7549 (
            .O(N__47572),
            .I(\ppm_encoder_1.un1_elevator_cry_12 ));
    InMux I__7548 (
            .O(N__47569),
            .I(\ppm_encoder_1.un1_elevator_cry_13 ));
    InMux I__7547 (
            .O(N__47566),
            .I(N__47563));
    LocalMux I__7546 (
            .O(N__47563),
            .I(N__47560));
    Span4Mux_h I__7545 (
            .O(N__47560),
            .I(N__47557));
    Odrv4 I__7544 (
            .O(N__47557),
            .I(\ppm_encoder_1.elevatorZ0Z_14 ));
    CascadeMux I__7543 (
            .O(N__47554),
            .I(N__47550));
    InMux I__7542 (
            .O(N__47553),
            .I(N__47546));
    InMux I__7541 (
            .O(N__47550),
            .I(N__47543));
    InMux I__7540 (
            .O(N__47549),
            .I(N__47540));
    LocalMux I__7539 (
            .O(N__47546),
            .I(N__47537));
    LocalMux I__7538 (
            .O(N__47543),
            .I(N__47534));
    LocalMux I__7537 (
            .O(N__47540),
            .I(N__47529));
    Span4Mux_v I__7536 (
            .O(N__47537),
            .I(N__47529));
    Span4Mux_h I__7535 (
            .O(N__47534),
            .I(N__47526));
    Odrv4 I__7534 (
            .O(N__47529),
            .I(\ppm_encoder_1.elevatorZ0Z_3 ));
    Odrv4 I__7533 (
            .O(N__47526),
            .I(\ppm_encoder_1.elevatorZ0Z_3 ));
    InMux I__7532 (
            .O(N__47521),
            .I(N__47517));
    InMux I__7531 (
            .O(N__47520),
            .I(N__47513));
    LocalMux I__7530 (
            .O(N__47517),
            .I(N__47509));
    InMux I__7529 (
            .O(N__47516),
            .I(N__47505));
    LocalMux I__7528 (
            .O(N__47513),
            .I(N__47502));
    InMux I__7527 (
            .O(N__47512),
            .I(N__47499));
    Span4Mux_v I__7526 (
            .O(N__47509),
            .I(N__47496));
    InMux I__7525 (
            .O(N__47508),
            .I(N__47493));
    LocalMux I__7524 (
            .O(N__47505),
            .I(N__47490));
    Span4Mux_v I__7523 (
            .O(N__47502),
            .I(N__47487));
    LocalMux I__7522 (
            .O(N__47499),
            .I(N__47484));
    Span4Mux_h I__7521 (
            .O(N__47496),
            .I(N__47475));
    LocalMux I__7520 (
            .O(N__47493),
            .I(N__47475));
    Span4Mux_v I__7519 (
            .O(N__47490),
            .I(N__47468));
    Span4Mux_h I__7518 (
            .O(N__47487),
            .I(N__47468));
    Span4Mux_s2_v I__7517 (
            .O(N__47484),
            .I(N__47468));
    InMux I__7516 (
            .O(N__47483),
            .I(N__47459));
    InMux I__7515 (
            .O(N__47482),
            .I(N__47459));
    InMux I__7514 (
            .O(N__47481),
            .I(N__47459));
    InMux I__7513 (
            .O(N__47480),
            .I(N__47459));
    Odrv4 I__7512 (
            .O(N__47475),
            .I(\ppm_encoder_1.N_513 ));
    Odrv4 I__7511 (
            .O(N__47468),
            .I(\ppm_encoder_1.N_513 ));
    LocalMux I__7510 (
            .O(N__47459),
            .I(\ppm_encoder_1.N_513 ));
    CascadeMux I__7509 (
            .O(N__47452),
            .I(N__47448));
    CascadeMux I__7508 (
            .O(N__47451),
            .I(N__47442));
    InMux I__7507 (
            .O(N__47448),
            .I(N__47439));
    InMux I__7506 (
            .O(N__47447),
            .I(N__47424));
    InMux I__7505 (
            .O(N__47446),
            .I(N__47424));
    InMux I__7504 (
            .O(N__47445),
            .I(N__47424));
    InMux I__7503 (
            .O(N__47442),
            .I(N__47421));
    LocalMux I__7502 (
            .O(N__47439),
            .I(N__47418));
    InMux I__7501 (
            .O(N__47438),
            .I(N__47415));
    InMux I__7500 (
            .O(N__47437),
            .I(N__47412));
    InMux I__7499 (
            .O(N__47436),
            .I(N__47404));
    InMux I__7498 (
            .O(N__47435),
            .I(N__47404));
    InMux I__7497 (
            .O(N__47434),
            .I(N__47399));
    InMux I__7496 (
            .O(N__47433),
            .I(N__47399));
    InMux I__7495 (
            .O(N__47432),
            .I(N__47394));
    InMux I__7494 (
            .O(N__47431),
            .I(N__47391));
    LocalMux I__7493 (
            .O(N__47424),
            .I(N__47388));
    LocalMux I__7492 (
            .O(N__47421),
            .I(N__47379));
    Span4Mux_s1_v I__7491 (
            .O(N__47418),
            .I(N__47379));
    LocalMux I__7490 (
            .O(N__47415),
            .I(N__47379));
    LocalMux I__7489 (
            .O(N__47412),
            .I(N__47379));
    InMux I__7488 (
            .O(N__47411),
            .I(N__47372));
    InMux I__7487 (
            .O(N__47410),
            .I(N__47372));
    InMux I__7486 (
            .O(N__47409),
            .I(N__47372));
    LocalMux I__7485 (
            .O(N__47404),
            .I(N__47369));
    LocalMux I__7484 (
            .O(N__47399),
            .I(N__47366));
    InMux I__7483 (
            .O(N__47398),
            .I(N__47361));
    InMux I__7482 (
            .O(N__47397),
            .I(N__47361));
    LocalMux I__7481 (
            .O(N__47394),
            .I(N__47358));
    LocalMux I__7480 (
            .O(N__47391),
            .I(N__47351));
    Span4Mux_h I__7479 (
            .O(N__47388),
            .I(N__47344));
    Span4Mux_v I__7478 (
            .O(N__47379),
            .I(N__47344));
    LocalMux I__7477 (
            .O(N__47372),
            .I(N__47344));
    Span12Mux_h I__7476 (
            .O(N__47369),
            .I(N__47339));
    Span4Mux_s3_v I__7475 (
            .O(N__47366),
            .I(N__47332));
    LocalMux I__7474 (
            .O(N__47361),
            .I(N__47332));
    Span4Mux_v I__7473 (
            .O(N__47358),
            .I(N__47332));
    InMux I__7472 (
            .O(N__47357),
            .I(N__47327));
    InMux I__7471 (
            .O(N__47356),
            .I(N__47327));
    InMux I__7470 (
            .O(N__47355),
            .I(N__47324));
    InMux I__7469 (
            .O(N__47354),
            .I(N__47321));
    Span4Mux_v I__7468 (
            .O(N__47351),
            .I(N__47316));
    Span4Mux_h I__7467 (
            .O(N__47344),
            .I(N__47316));
    InMux I__7466 (
            .O(N__47343),
            .I(N__47311));
    InMux I__7465 (
            .O(N__47342),
            .I(N__47311));
    Odrv12 I__7464 (
            .O(N__47339),
            .I(\ppm_encoder_1.N_300 ));
    Odrv4 I__7463 (
            .O(N__47332),
            .I(\ppm_encoder_1.N_300 ));
    LocalMux I__7462 (
            .O(N__47327),
            .I(\ppm_encoder_1.N_300 ));
    LocalMux I__7461 (
            .O(N__47324),
            .I(\ppm_encoder_1.N_300 ));
    LocalMux I__7460 (
            .O(N__47321),
            .I(\ppm_encoder_1.N_300 ));
    Odrv4 I__7459 (
            .O(N__47316),
            .I(\ppm_encoder_1.N_300 ));
    LocalMux I__7458 (
            .O(N__47311),
            .I(\ppm_encoder_1.N_300 ));
    InMux I__7457 (
            .O(N__47296),
            .I(N__47293));
    LocalMux I__7456 (
            .O(N__47293),
            .I(\ppm_encoder_1.pulses2count_9_0_0_0_3 ));
    InMux I__7455 (
            .O(N__47290),
            .I(N__47287));
    LocalMux I__7454 (
            .O(N__47287),
            .I(N__47284));
    Span4Mux_h I__7453 (
            .O(N__47284),
            .I(N__47281));
    Odrv4 I__7452 (
            .O(N__47281),
            .I(\ppm_encoder_1.un1_elevator_cry_0_THRU_CO ));
    InMux I__7451 (
            .O(N__47278),
            .I(\ppm_encoder_1.un1_elevator_cry_0 ));
    InMux I__7450 (
            .O(N__47275),
            .I(N__47272));
    LocalMux I__7449 (
            .O(N__47272),
            .I(N__47269));
    Span4Mux_h I__7448 (
            .O(N__47269),
            .I(N__47266));
    Odrv4 I__7447 (
            .O(N__47266),
            .I(\ppm_encoder_1.un1_elevator_cry_1_THRU_CO ));
    InMux I__7446 (
            .O(N__47263),
            .I(\ppm_encoder_1.un1_elevator_cry_1 ));
    InMux I__7445 (
            .O(N__47260),
            .I(N__47257));
    LocalMux I__7444 (
            .O(N__47257),
            .I(N__47254));
    Odrv12 I__7443 (
            .O(N__47254),
            .I(\ppm_encoder_1.un1_elevator_cry_2_THRU_CO ));
    InMux I__7442 (
            .O(N__47251),
            .I(\ppm_encoder_1.un1_elevator_cry_2 ));
    CascadeMux I__7441 (
            .O(N__47248),
            .I(N__47245));
    InMux I__7440 (
            .O(N__47245),
            .I(N__47242));
    LocalMux I__7439 (
            .O(N__47242),
            .I(N__47239));
    Odrv12 I__7438 (
            .O(N__47239),
            .I(\ppm_encoder_1.un1_elevator_cry_3_THRU_CO ));
    InMux I__7437 (
            .O(N__47236),
            .I(\ppm_encoder_1.un1_elevator_cry_3 ));
    InMux I__7436 (
            .O(N__47233),
            .I(\ppm_encoder_1.un1_elevator_cry_4 ));
    InMux I__7435 (
            .O(N__47230),
            .I(N__47225));
    InMux I__7434 (
            .O(N__47229),
            .I(N__47220));
    InMux I__7433 (
            .O(N__47228),
            .I(N__47220));
    LocalMux I__7432 (
            .O(N__47225),
            .I(N__47217));
    LocalMux I__7431 (
            .O(N__47220),
            .I(\ppm_encoder_1.elevatorZ0Z_0 ));
    Odrv4 I__7430 (
            .O(N__47217),
            .I(\ppm_encoder_1.elevatorZ0Z_0 ));
    CascadeMux I__7429 (
            .O(N__47212),
            .I(N__47209));
    InMux I__7428 (
            .O(N__47209),
            .I(N__47206));
    LocalMux I__7427 (
            .O(N__47206),
            .I(N__47203));
    Span4Mux_v I__7426 (
            .O(N__47203),
            .I(N__47200));
    Odrv4 I__7425 (
            .O(N__47200),
            .I(\ppm_encoder_1.N_393 ));
    CascadeMux I__7424 (
            .O(N__47197),
            .I(N__47194));
    InMux I__7423 (
            .O(N__47194),
            .I(N__47190));
    InMux I__7422 (
            .O(N__47193),
            .I(N__47187));
    LocalMux I__7421 (
            .O(N__47190),
            .I(N__47183));
    LocalMux I__7420 (
            .O(N__47187),
            .I(N__47180));
    CascadeMux I__7419 (
            .O(N__47186),
            .I(N__47177));
    Span4Mux_h I__7418 (
            .O(N__47183),
            .I(N__47174));
    Span4Mux_v I__7417 (
            .O(N__47180),
            .I(N__47171));
    InMux I__7416 (
            .O(N__47177),
            .I(N__47168));
    Span4Mux_h I__7415 (
            .O(N__47174),
            .I(N__47165));
    Span4Mux_h I__7414 (
            .O(N__47171),
            .I(N__47160));
    LocalMux I__7413 (
            .O(N__47168),
            .I(N__47160));
    Span4Mux_h I__7412 (
            .O(N__47165),
            .I(N__47157));
    Span4Mux_h I__7411 (
            .O(N__47160),
            .I(N__47154));
    Odrv4 I__7410 (
            .O(N__47157),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_ns_0 ));
    Odrv4 I__7409 (
            .O(N__47154),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_ns_0 ));
    CascadeMux I__7408 (
            .O(N__47149),
            .I(N__47146));
    InMux I__7407 (
            .O(N__47146),
            .I(N__47143));
    LocalMux I__7406 (
            .O(N__47143),
            .I(N__47139));
    InMux I__7405 (
            .O(N__47142),
            .I(N__47136));
    Span4Mux_v I__7404 (
            .O(N__47139),
            .I(N__47130));
    LocalMux I__7403 (
            .O(N__47136),
            .I(N__47130));
    InMux I__7402 (
            .O(N__47135),
            .I(N__47126));
    Span4Mux_v I__7401 (
            .O(N__47130),
            .I(N__47123));
    InMux I__7400 (
            .O(N__47129),
            .I(N__47120));
    LocalMux I__7399 (
            .O(N__47126),
            .I(N__47117));
    Span4Mux_h I__7398 (
            .O(N__47123),
            .I(N__47112));
    LocalMux I__7397 (
            .O(N__47120),
            .I(N__47112));
    Span4Mux_v I__7396 (
            .O(N__47117),
            .I(N__47109));
    Sp12to4 I__7395 (
            .O(N__47112),
            .I(N__47106));
    Odrv4 I__7394 (
            .O(N__47109),
            .I(\ppm_encoder_1.N_56 ));
    Odrv12 I__7393 (
            .O(N__47106),
            .I(\ppm_encoder_1.N_56 ));
    CascadeMux I__7392 (
            .O(N__47101),
            .I(N__47098));
    InMux I__7391 (
            .O(N__47098),
            .I(N__47095));
    LocalMux I__7390 (
            .O(N__47095),
            .I(N__47092));
    Odrv12 I__7389 (
            .O(N__47092),
            .I(\ppm_encoder_1.N_378 ));
    InMux I__7388 (
            .O(N__47089),
            .I(N__47086));
    LocalMux I__7387 (
            .O(N__47086),
            .I(N__47081));
    InMux I__7386 (
            .O(N__47085),
            .I(N__47078));
    InMux I__7385 (
            .O(N__47084),
            .I(N__47075));
    Span4Mux_v I__7384 (
            .O(N__47081),
            .I(N__47072));
    LocalMux I__7383 (
            .O(N__47078),
            .I(N__47069));
    LocalMux I__7382 (
            .O(N__47075),
            .I(\ppm_encoder_1.rudderZ0Z_10 ));
    Odrv4 I__7381 (
            .O(N__47072),
            .I(\ppm_encoder_1.rudderZ0Z_10 ));
    Odrv4 I__7380 (
            .O(N__47069),
            .I(\ppm_encoder_1.rudderZ0Z_10 ));
    CascadeMux I__7379 (
            .O(N__47062),
            .I(N__47059));
    InMux I__7378 (
            .O(N__47059),
            .I(N__47056));
    LocalMux I__7377 (
            .O(N__47056),
            .I(N__47053));
    Odrv12 I__7376 (
            .O(N__47053),
            .I(\ppm_encoder_1.N_406 ));
    InMux I__7375 (
            .O(N__47050),
            .I(N__47047));
    LocalMux I__7374 (
            .O(N__47047),
            .I(N__47043));
    CascadeMux I__7373 (
            .O(N__47046),
            .I(N__47040));
    Span4Mux_h I__7372 (
            .O(N__47043),
            .I(N__47037));
    InMux I__7371 (
            .O(N__47040),
            .I(N__47034));
    Odrv4 I__7370 (
            .O(N__47037),
            .I(scaler_4_data_4));
    LocalMux I__7369 (
            .O(N__47034),
            .I(scaler_4_data_4));
    CascadeMux I__7368 (
            .O(N__47029),
            .I(N__47026));
    InMux I__7367 (
            .O(N__47026),
            .I(N__47022));
    InMux I__7366 (
            .O(N__47025),
            .I(N__47019));
    LocalMux I__7365 (
            .O(N__47022),
            .I(N__47016));
    LocalMux I__7364 (
            .O(N__47019),
            .I(\ppm_encoder_1.rudderZ0Z_4 ));
    Odrv4 I__7363 (
            .O(N__47016),
            .I(\ppm_encoder_1.rudderZ0Z_4 ));
    CascadeMux I__7362 (
            .O(N__47011),
            .I(N__47008));
    InMux I__7361 (
            .O(N__47008),
            .I(N__47005));
    LocalMux I__7360 (
            .O(N__47005),
            .I(N__47002));
    Span4Mux_v I__7359 (
            .O(N__47002),
            .I(N__46999));
    Odrv4 I__7358 (
            .O(N__46999),
            .I(\ppm_encoder_1.N_420 ));
    InMux I__7357 (
            .O(N__46996),
            .I(N__46991));
    InMux I__7356 (
            .O(N__46995),
            .I(N__46988));
    CascadeMux I__7355 (
            .O(N__46994),
            .I(N__46985));
    LocalMux I__7354 (
            .O(N__46991),
            .I(N__46982));
    LocalMux I__7353 (
            .O(N__46988),
            .I(N__46979));
    InMux I__7352 (
            .O(N__46985),
            .I(N__46976));
    Span12Mux_h I__7351 (
            .O(N__46982),
            .I(N__46971));
    Span12Mux_s8_h I__7350 (
            .O(N__46979),
            .I(N__46971));
    LocalMux I__7349 (
            .O(N__46976),
            .I(\ppm_encoder_1.rudderZ0Z_8 ));
    Odrv12 I__7348 (
            .O(N__46971),
            .I(\ppm_encoder_1.rudderZ0Z_8 ));
    CascadeMux I__7347 (
            .O(N__46966),
            .I(N__46963));
    InMux I__7346 (
            .O(N__46963),
            .I(N__46959));
    InMux I__7345 (
            .O(N__46962),
            .I(N__46956));
    LocalMux I__7344 (
            .O(N__46959),
            .I(N__46952));
    LocalMux I__7343 (
            .O(N__46956),
            .I(N__46949));
    InMux I__7342 (
            .O(N__46955),
            .I(N__46946));
    Span4Mux_h I__7341 (
            .O(N__46952),
            .I(N__46943));
    Span4Mux_h I__7340 (
            .O(N__46949),
            .I(N__46940));
    LocalMux I__7339 (
            .O(N__46946),
            .I(\ppm_encoder_1.rudderZ0Z_9 ));
    Odrv4 I__7338 (
            .O(N__46943),
            .I(\ppm_encoder_1.rudderZ0Z_9 ));
    Odrv4 I__7337 (
            .O(N__46940),
            .I(\ppm_encoder_1.rudderZ0Z_9 ));
    InMux I__7336 (
            .O(N__46933),
            .I(N__46930));
    LocalMux I__7335 (
            .O(N__46930),
            .I(\ppm_encoder_1.N_425 ));
    InMux I__7334 (
            .O(N__46927),
            .I(N__46924));
    LocalMux I__7333 (
            .O(N__46924),
            .I(N__46921));
    Span4Mux_v I__7332 (
            .O(N__46921),
            .I(N__46918));
    Span4Mux_h I__7331 (
            .O(N__46918),
            .I(N__46915));
    Odrv4 I__7330 (
            .O(N__46915),
            .I(\ppm_encoder_1.pulses2count_9_i_2_9 ));
    CascadeMux I__7329 (
            .O(N__46912),
            .I(N__46909));
    InMux I__7328 (
            .O(N__46909),
            .I(N__46904));
    CascadeMux I__7327 (
            .O(N__46908),
            .I(N__46901));
    CascadeMux I__7326 (
            .O(N__46907),
            .I(N__46898));
    LocalMux I__7325 (
            .O(N__46904),
            .I(N__46895));
    InMux I__7324 (
            .O(N__46901),
            .I(N__46889));
    InMux I__7323 (
            .O(N__46898),
            .I(N__46889));
    Span4Mux_h I__7322 (
            .O(N__46895),
            .I(N__46886));
    InMux I__7321 (
            .O(N__46894),
            .I(N__46883));
    LocalMux I__7320 (
            .O(N__46889),
            .I(N__46880));
    Span4Mux_h I__7319 (
            .O(N__46886),
            .I(N__46877));
    LocalMux I__7318 (
            .O(N__46883),
            .I(N__46874));
    Span4Mux_h I__7317 (
            .O(N__46880),
            .I(N__46871));
    Odrv4 I__7316 (
            .O(N__46877),
            .I(\ppm_encoder_1.N_275 ));
    Odrv12 I__7315 (
            .O(N__46874),
            .I(\ppm_encoder_1.N_275 ));
    Odrv4 I__7314 (
            .O(N__46871),
            .I(\ppm_encoder_1.N_275 ));
    CascadeMux I__7313 (
            .O(N__46864),
            .I(N__46861));
    InMux I__7312 (
            .O(N__46861),
            .I(N__46858));
    LocalMux I__7311 (
            .O(N__46858),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_16 ));
    InMux I__7310 (
            .O(N__46855),
            .I(N__46852));
    LocalMux I__7309 (
            .O(N__46852),
            .I(N__46849));
    Span4Mux_h I__7308 (
            .O(N__46849),
            .I(N__46846));
    Odrv4 I__7307 (
            .O(N__46846),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_16 ));
    InMux I__7306 (
            .O(N__46843),
            .I(N__46840));
    LocalMux I__7305 (
            .O(N__46840),
            .I(N__46837));
    Span4Mux_h I__7304 (
            .O(N__46837),
            .I(N__46834));
    Odrv4 I__7303 (
            .O(N__46834),
            .I(\ppm_encoder_1.un1_init_pulses_11_8 ));
    InMux I__7302 (
            .O(N__46831),
            .I(N__46828));
    LocalMux I__7301 (
            .O(N__46828),
            .I(\ppm_encoder_1.un1_init_pulses_10_8 ));
    InMux I__7300 (
            .O(N__46825),
            .I(N__46822));
    LocalMux I__7299 (
            .O(N__46822),
            .I(N__46819));
    Span4Mux_v I__7298 (
            .O(N__46819),
            .I(N__46816));
    Odrv4 I__7297 (
            .O(N__46816),
            .I(\ppm_encoder_1.un1_init_pulses_11_11 ));
    InMux I__7296 (
            .O(N__46813),
            .I(N__46810));
    LocalMux I__7295 (
            .O(N__46810),
            .I(\ppm_encoder_1.un1_init_pulses_10_11 ));
    CascadeMux I__7294 (
            .O(N__46807),
            .I(N__46804));
    InMux I__7293 (
            .O(N__46804),
            .I(N__46800));
    CascadeMux I__7292 (
            .O(N__46803),
            .I(N__46797));
    LocalMux I__7291 (
            .O(N__46800),
            .I(N__46793));
    InMux I__7290 (
            .O(N__46797),
            .I(N__46789));
    InMux I__7289 (
            .O(N__46796),
            .I(N__46786));
    Span4Mux_h I__7288 (
            .O(N__46793),
            .I(N__46783));
    CascadeMux I__7287 (
            .O(N__46792),
            .I(N__46780));
    LocalMux I__7286 (
            .O(N__46789),
            .I(N__46777));
    LocalMux I__7285 (
            .O(N__46786),
            .I(N__46772));
    Span4Mux_s2_v I__7284 (
            .O(N__46783),
            .I(N__46772));
    InMux I__7283 (
            .O(N__46780),
            .I(N__46769));
    Span4Mux_h I__7282 (
            .O(N__46777),
            .I(N__46766));
    Odrv4 I__7281 (
            .O(N__46772),
            .I(\ppm_encoder_1.init_pulsesZ0Z_11 ));
    LocalMux I__7280 (
            .O(N__46769),
            .I(\ppm_encoder_1.init_pulsesZ0Z_11 ));
    Odrv4 I__7279 (
            .O(N__46766),
            .I(\ppm_encoder_1.init_pulsesZ0Z_11 ));
    InMux I__7278 (
            .O(N__46759),
            .I(N__46756));
    LocalMux I__7277 (
            .O(N__46756),
            .I(N__46753));
    Span4Mux_h I__7276 (
            .O(N__46753),
            .I(N__46750));
    Odrv4 I__7275 (
            .O(N__46750),
            .I(\ppm_encoder_1.un1_init_pulses_11_12 ));
    InMux I__7274 (
            .O(N__46747),
            .I(N__46744));
    LocalMux I__7273 (
            .O(N__46744),
            .I(\ppm_encoder_1.un1_init_pulses_10_12 ));
    InMux I__7272 (
            .O(N__46741),
            .I(N__46736));
    InMux I__7271 (
            .O(N__46740),
            .I(N__46733));
    CascadeMux I__7270 (
            .O(N__46739),
            .I(N__46730));
    LocalMux I__7269 (
            .O(N__46736),
            .I(N__46727));
    LocalMux I__7268 (
            .O(N__46733),
            .I(N__46724));
    InMux I__7267 (
            .O(N__46730),
            .I(N__46721));
    Span4Mux_h I__7266 (
            .O(N__46727),
            .I(N__46718));
    Span4Mux_v I__7265 (
            .O(N__46724),
            .I(N__46715));
    LocalMux I__7264 (
            .O(N__46721),
            .I(N__46710));
    Span4Mux_v I__7263 (
            .O(N__46718),
            .I(N__46710));
    Odrv4 I__7262 (
            .O(N__46715),
            .I(\ppm_encoder_1.aileronZ0Z_4 ));
    Odrv4 I__7261 (
            .O(N__46710),
            .I(\ppm_encoder_1.aileronZ0Z_4 ));
    InMux I__7260 (
            .O(N__46705),
            .I(N__46701));
    CascadeMux I__7259 (
            .O(N__46704),
            .I(N__46697));
    LocalMux I__7258 (
            .O(N__46701),
            .I(N__46694));
    InMux I__7257 (
            .O(N__46700),
            .I(N__46691));
    InMux I__7256 (
            .O(N__46697),
            .I(N__46688));
    Span4Mux_h I__7255 (
            .O(N__46694),
            .I(N__46685));
    LocalMux I__7254 (
            .O(N__46691),
            .I(\ppm_encoder_1.elevatorZ0Z_4 ));
    LocalMux I__7253 (
            .O(N__46688),
            .I(\ppm_encoder_1.elevatorZ0Z_4 ));
    Odrv4 I__7252 (
            .O(N__46685),
            .I(\ppm_encoder_1.elevatorZ0Z_4 ));
    InMux I__7251 (
            .O(N__46678),
            .I(\ppm_encoder_1.counter24_0_N_2 ));
    InMux I__7250 (
            .O(N__46675),
            .I(N__46672));
    LocalMux I__7249 (
            .O(N__46672),
            .I(\ppm_encoder_1.counter24_0_I_51_c_RNOZ0 ));
    InMux I__7248 (
            .O(N__46669),
            .I(N__46666));
    LocalMux I__7247 (
            .O(N__46666),
            .I(\ppm_encoder_1.counter24_0_I_39_c_RNOZ0 ));
    InMux I__7246 (
            .O(N__46663),
            .I(N__46660));
    LocalMux I__7245 (
            .O(N__46660),
            .I(N__46657));
    Span4Mux_v I__7244 (
            .O(N__46657),
            .I(N__46654));
    Odrv4 I__7243 (
            .O(N__46654),
            .I(\ppm_encoder_1.un1_init_pulses_11_2 ));
    InMux I__7242 (
            .O(N__46651),
            .I(N__46648));
    LocalMux I__7241 (
            .O(N__46648),
            .I(\ppm_encoder_1.un1_init_pulses_10_2 ));
    CascadeMux I__7240 (
            .O(N__46645),
            .I(N__46639));
    InMux I__7239 (
            .O(N__46644),
            .I(N__46634));
    InMux I__7238 (
            .O(N__46643),
            .I(N__46634));
    InMux I__7237 (
            .O(N__46642),
            .I(N__46629));
    InMux I__7236 (
            .O(N__46639),
            .I(N__46629));
    LocalMux I__7235 (
            .O(N__46634),
            .I(N__46626));
    LocalMux I__7234 (
            .O(N__46629),
            .I(N__46623));
    Span4Mux_v I__7233 (
            .O(N__46626),
            .I(N__46620));
    Span4Mux_s2_v I__7232 (
            .O(N__46623),
            .I(N__46617));
    Span4Mux_h I__7231 (
            .O(N__46620),
            .I(N__46612));
    Span4Mux_h I__7230 (
            .O(N__46617),
            .I(N__46612));
    Odrv4 I__7229 (
            .O(N__46612),
            .I(\ppm_encoder_1.init_pulsesZ0Z_2 ));
    CascadeMux I__7228 (
            .O(N__46609),
            .I(N__46606));
    InMux I__7227 (
            .O(N__46606),
            .I(N__46603));
    LocalMux I__7226 (
            .O(N__46603),
            .I(N__46600));
    Span4Mux_h I__7225 (
            .O(N__46600),
            .I(N__46597));
    Odrv4 I__7224 (
            .O(N__46597),
            .I(\ppm_encoder_1.un1_init_pulses_11_5 ));
    InMux I__7223 (
            .O(N__46594),
            .I(N__46591));
    LocalMux I__7222 (
            .O(N__46591),
            .I(\ppm_encoder_1.un1_init_pulses_10_5 ));
    InMux I__7221 (
            .O(N__46588),
            .I(N__46585));
    LocalMux I__7220 (
            .O(N__46585),
            .I(N__46582));
    Span4Mux_h I__7219 (
            .O(N__46582),
            .I(N__46579));
    Odrv4 I__7218 (
            .O(N__46579),
            .I(\ppm_encoder_1.un1_init_pulses_11_6 ));
    InMux I__7217 (
            .O(N__46576),
            .I(N__46573));
    LocalMux I__7216 (
            .O(N__46573),
            .I(\ppm_encoder_1.un1_init_pulses_10_6 ));
    CascadeMux I__7215 (
            .O(N__46570),
            .I(N__46567));
    InMux I__7214 (
            .O(N__46567),
            .I(N__46564));
    LocalMux I__7213 (
            .O(N__46564),
            .I(N__46561));
    Span4Mux_h I__7212 (
            .O(N__46561),
            .I(N__46558));
    Odrv4 I__7211 (
            .O(N__46558),
            .I(\ppm_encoder_1.un1_init_pulses_11_7 ));
    InMux I__7210 (
            .O(N__46555),
            .I(N__46552));
    LocalMux I__7209 (
            .O(N__46552),
            .I(\ppm_encoder_1.un1_init_pulses_10_7 ));
    InMux I__7208 (
            .O(N__46549),
            .I(N__46546));
    LocalMux I__7207 (
            .O(N__46546),
            .I(\ppm_encoder_1.un1_init_pulses_10_9 ));
    InMux I__7206 (
            .O(N__46543),
            .I(N__46540));
    LocalMux I__7205 (
            .O(N__46540),
            .I(N__46537));
    Span4Mux_h I__7204 (
            .O(N__46537),
            .I(N__46534));
    Odrv4 I__7203 (
            .O(N__46534),
            .I(\ppm_encoder_1.un1_init_pulses_11_9 ));
    InMux I__7202 (
            .O(N__46531),
            .I(N__46528));
    LocalMux I__7201 (
            .O(N__46528),
            .I(N__46524));
    InMux I__7200 (
            .O(N__46527),
            .I(N__46521));
    Span4Mux_v I__7199 (
            .O(N__46524),
            .I(N__46517));
    LocalMux I__7198 (
            .O(N__46521),
            .I(N__46514));
    CascadeMux I__7197 (
            .O(N__46520),
            .I(N__46510));
    Span4Mux_h I__7196 (
            .O(N__46517),
            .I(N__46507));
    Span4Mux_v I__7195 (
            .O(N__46514),
            .I(N__46504));
    InMux I__7194 (
            .O(N__46513),
            .I(N__46499));
    InMux I__7193 (
            .O(N__46510),
            .I(N__46499));
    Sp12to4 I__7192 (
            .O(N__46507),
            .I(N__46496));
    Span4Mux_h I__7191 (
            .O(N__46504),
            .I(N__46493));
    LocalMux I__7190 (
            .O(N__46499),
            .I(N__46490));
    Odrv12 I__7189 (
            .O(N__46496),
            .I(\ppm_encoder_1.init_pulsesZ0Z_9 ));
    Odrv4 I__7188 (
            .O(N__46493),
            .I(\ppm_encoder_1.init_pulsesZ0Z_9 ));
    Odrv4 I__7187 (
            .O(N__46490),
            .I(\ppm_encoder_1.init_pulsesZ0Z_9 ));
    InMux I__7186 (
            .O(N__46483),
            .I(N__46480));
    LocalMux I__7185 (
            .O(N__46480),
            .I(N__46476));
    CascadeMux I__7184 (
            .O(N__46479),
            .I(N__46473));
    Span4Mux_s3_v I__7183 (
            .O(N__46476),
            .I(N__46469));
    InMux I__7182 (
            .O(N__46473),
            .I(N__46466));
    InMux I__7181 (
            .O(N__46472),
            .I(N__46463));
    Span4Mux_h I__7180 (
            .O(N__46469),
            .I(N__46458));
    LocalMux I__7179 (
            .O(N__46466),
            .I(N__46458));
    LocalMux I__7178 (
            .O(N__46463),
            .I(N__46453));
    Span4Mux_v I__7177 (
            .O(N__46458),
            .I(N__46453));
    Odrv4 I__7176 (
            .O(N__46453),
            .I(\ppm_encoder_1.throttleZ0Z_10 ));
    InMux I__7175 (
            .O(N__46450),
            .I(N__46447));
    LocalMux I__7174 (
            .O(N__46447),
            .I(\dron_frame_decoder_1.state_ns_0_i_a2_0_3_3 ));
    InMux I__7173 (
            .O(N__46444),
            .I(N__46432));
    InMux I__7172 (
            .O(N__46443),
            .I(N__46432));
    InMux I__7171 (
            .O(N__46442),
            .I(N__46432));
    InMux I__7170 (
            .O(N__46441),
            .I(N__46427));
    InMux I__7169 (
            .O(N__46440),
            .I(N__46427));
    InMux I__7168 (
            .O(N__46439),
            .I(N__46424));
    LocalMux I__7167 (
            .O(N__46432),
            .I(\dron_frame_decoder_1.stateZ0Z_6 ));
    LocalMux I__7166 (
            .O(N__46427),
            .I(\dron_frame_decoder_1.stateZ0Z_6 ));
    LocalMux I__7165 (
            .O(N__46424),
            .I(\dron_frame_decoder_1.stateZ0Z_6 ));
    InMux I__7164 (
            .O(N__46417),
            .I(N__46414));
    LocalMux I__7163 (
            .O(N__46414),
            .I(N__46411));
    Span4Mux_v I__7162 (
            .O(N__46411),
            .I(N__46408));
    Span4Mux_v I__7161 (
            .O(N__46408),
            .I(N__46405));
    Odrv4 I__7160 (
            .O(N__46405),
            .I(\pid_alt.state_RNIFCSD1Z0Z_0 ));
    InMux I__7159 (
            .O(N__46402),
            .I(N__46399));
    LocalMux I__7158 (
            .O(N__46399),
            .I(N__46396));
    Span4Mux_h I__7157 (
            .O(N__46396),
            .I(N__46393));
    Odrv4 I__7156 (
            .O(N__46393),
            .I(\Commands_frame_decoder.state_ns_0_a3_0_1 ));
    InMux I__7155 (
            .O(N__46390),
            .I(N__46387));
    LocalMux I__7154 (
            .O(N__46387),
            .I(N__46384));
    Sp12to4 I__7153 (
            .O(N__46384),
            .I(N__46381));
    Span12Mux_v I__7152 (
            .O(N__46381),
            .I(N__46378));
    Odrv12 I__7151 (
            .O(N__46378),
            .I(\pid_front.O_0_6 ));
    InMux I__7150 (
            .O(N__46375),
            .I(N__46372));
    LocalMux I__7149 (
            .O(N__46372),
            .I(N__46369));
    Odrv12 I__7148 (
            .O(N__46369),
            .I(drone_altitude_i_9));
    InMux I__7147 (
            .O(N__46366),
            .I(N__46362));
    InMux I__7146 (
            .O(N__46365),
            .I(N__46359));
    LocalMux I__7145 (
            .O(N__46362),
            .I(N__46356));
    LocalMux I__7144 (
            .O(N__46359),
            .I(N__46353));
    Odrv4 I__7143 (
            .O(N__46356),
            .I(\dron_frame_decoder_1.state_RNI4N6KZ0Z_2 ));
    Odrv4 I__7142 (
            .O(N__46353),
            .I(\dron_frame_decoder_1.state_RNI4N6KZ0Z_2 ));
    InMux I__7141 (
            .O(N__46348),
            .I(N__46345));
    LocalMux I__7140 (
            .O(N__46345),
            .I(\dron_frame_decoder_1.un1_sink_data_valid_5_i_0 ));
    CascadeMux I__7139 (
            .O(N__46342),
            .I(\dron_frame_decoder_1.un1_sink_data_valid_5_i_0_cascade_ ));
    InMux I__7138 (
            .O(N__46339),
            .I(N__46335));
    CascadeMux I__7137 (
            .O(N__46338),
            .I(N__46331));
    LocalMux I__7136 (
            .O(N__46335),
            .I(N__46326));
    InMux I__7135 (
            .O(N__46334),
            .I(N__46321));
    InMux I__7134 (
            .O(N__46331),
            .I(N__46321));
    InMux I__7133 (
            .O(N__46330),
            .I(N__46316));
    InMux I__7132 (
            .O(N__46329),
            .I(N__46316));
    Span4Mux_h I__7131 (
            .O(N__46326),
            .I(N__46313));
    LocalMux I__7130 (
            .O(N__46321),
            .I(\dron_frame_decoder_1.stateZ0Z_4 ));
    LocalMux I__7129 (
            .O(N__46316),
            .I(\dron_frame_decoder_1.stateZ0Z_4 ));
    Odrv4 I__7128 (
            .O(N__46313),
            .I(\dron_frame_decoder_1.stateZ0Z_4 ));
    InMux I__7127 (
            .O(N__46306),
            .I(N__46294));
    InMux I__7126 (
            .O(N__46305),
            .I(N__46294));
    InMux I__7125 (
            .O(N__46304),
            .I(N__46294));
    InMux I__7124 (
            .O(N__46303),
            .I(N__46294));
    LocalMux I__7123 (
            .O(N__46294),
            .I(\dron_frame_decoder_1.stateZ0Z_5 ));
    CascadeMux I__7122 (
            .O(N__46291),
            .I(\dron_frame_decoder_1.state_ns_0_i_a2_0_2_3_cascade_ ));
    CascadeMux I__7121 (
            .O(N__46288),
            .I(N__46283));
    InMux I__7120 (
            .O(N__46287),
            .I(N__46280));
    InMux I__7119 (
            .O(N__46286),
            .I(N__46275));
    InMux I__7118 (
            .O(N__46283),
            .I(N__46275));
    LocalMux I__7117 (
            .O(N__46280),
            .I(\dron_frame_decoder_1.stateZ0Z_3 ));
    LocalMux I__7116 (
            .O(N__46275),
            .I(\dron_frame_decoder_1.stateZ0Z_3 ));
    InMux I__7115 (
            .O(N__46270),
            .I(N__46256));
    InMux I__7114 (
            .O(N__46269),
            .I(N__46256));
    InMux I__7113 (
            .O(N__46268),
            .I(N__46256));
    InMux I__7112 (
            .O(N__46267),
            .I(N__46256));
    InMux I__7111 (
            .O(N__46266),
            .I(N__46251));
    InMux I__7110 (
            .O(N__46265),
            .I(N__46251));
    LocalMux I__7109 (
            .O(N__46256),
            .I(\uart_pc.timer_Count_RNIMQ8T1Z0Z_2 ));
    LocalMux I__7108 (
            .O(N__46251),
            .I(\uart_pc.timer_Count_RNIMQ8T1Z0Z_2 ));
    CascadeMux I__7107 (
            .O(N__46246),
            .I(N__46243));
    InMux I__7106 (
            .O(N__46243),
            .I(N__46239));
    InMux I__7105 (
            .O(N__46242),
            .I(N__46236));
    LocalMux I__7104 (
            .O(N__46239),
            .I(\uart_pc.data_AuxZ1Z_1 ));
    LocalMux I__7103 (
            .O(N__46236),
            .I(\uart_pc.data_AuxZ1Z_1 ));
    InMux I__7102 (
            .O(N__46231),
            .I(N__46228));
    LocalMux I__7101 (
            .O(N__46228),
            .I(N__46225));
    Span4Mux_h I__7100 (
            .O(N__46225),
            .I(N__46221));
    InMux I__7099 (
            .O(N__46224),
            .I(N__46218));
    Span4Mux_h I__7098 (
            .O(N__46221),
            .I(N__46215));
    LocalMux I__7097 (
            .O(N__46218),
            .I(\pid_alt.drone_altitude_i_0 ));
    Odrv4 I__7096 (
            .O(N__46215),
            .I(\pid_alt.drone_altitude_i_0 ));
    InMux I__7095 (
            .O(N__46210),
            .I(N__46207));
    LocalMux I__7094 (
            .O(N__46207),
            .I(N__46203));
    InMux I__7093 (
            .O(N__46206),
            .I(N__46200));
    Odrv12 I__7092 (
            .O(N__46203),
            .I(frame_decoder_OFF4data_7));
    LocalMux I__7091 (
            .O(N__46200),
            .I(frame_decoder_OFF4data_7));
    InMux I__7090 (
            .O(N__46195),
            .I(N__46192));
    LocalMux I__7089 (
            .O(N__46192),
            .I(N__46188));
    InMux I__7088 (
            .O(N__46191),
            .I(N__46185));
    Span12Mux_v I__7087 (
            .O(N__46188),
            .I(N__46182));
    LocalMux I__7086 (
            .O(N__46185),
            .I(N__46179));
    Odrv12 I__7085 (
            .O(N__46182),
            .I(frame_decoder_CH4data_7));
    Odrv4 I__7084 (
            .O(N__46179),
            .I(frame_decoder_CH4data_7));
    InMux I__7083 (
            .O(N__46174),
            .I(N__46171));
    LocalMux I__7082 (
            .O(N__46171),
            .I(N__46168));
    Span4Mux_v I__7081 (
            .O(N__46168),
            .I(N__46165));
    Odrv4 I__7080 (
            .O(N__46165),
            .I(\scaler_4.N_2928_i_l_ofxZ0 ));
    InMux I__7079 (
            .O(N__46162),
            .I(N__46159));
    LocalMux I__7078 (
            .O(N__46159),
            .I(N__46156));
    Odrv12 I__7077 (
            .O(N__46156),
            .I(drone_altitude_i_4));
    InMux I__7076 (
            .O(N__46153),
            .I(N__46150));
    LocalMux I__7075 (
            .O(N__46150),
            .I(N__46147));
    Odrv12 I__7074 (
            .O(N__46147),
            .I(drone_altitude_i_5));
    CascadeMux I__7073 (
            .O(N__46144),
            .I(N__46141));
    InMux I__7072 (
            .O(N__46141),
            .I(N__46138));
    LocalMux I__7071 (
            .O(N__46138),
            .I(N__46135));
    Span4Mux_h I__7070 (
            .O(N__46135),
            .I(N__46132));
    Odrv4 I__7069 (
            .O(N__46132),
            .I(drone_altitude_i_6));
    CascadeMux I__7068 (
            .O(N__46129),
            .I(N__46126));
    InMux I__7067 (
            .O(N__46126),
            .I(N__46123));
    LocalMux I__7066 (
            .O(N__46123),
            .I(N__46120));
    Odrv12 I__7065 (
            .O(N__46120),
            .I(drone_altitude_i_7));
    InMux I__7064 (
            .O(N__46117),
            .I(N__46114));
    LocalMux I__7063 (
            .O(N__46114),
            .I(N__46110));
    InMux I__7062 (
            .O(N__46113),
            .I(N__46107));
    Span4Mux_v I__7061 (
            .O(N__46110),
            .I(N__46104));
    LocalMux I__7060 (
            .O(N__46107),
            .I(N__46101));
    Span4Mux_v I__7059 (
            .O(N__46104),
            .I(N__46096));
    Span4Mux_v I__7058 (
            .O(N__46101),
            .I(N__46096));
    Span4Mux_h I__7057 (
            .O(N__46096),
            .I(N__46093));
    Span4Mux_h I__7056 (
            .O(N__46093),
            .I(N__46090));
    Span4Mux_h I__7055 (
            .O(N__46090),
            .I(N__46087));
    Odrv4 I__7054 (
            .O(N__46087),
            .I(xy_kd_1));
    InMux I__7053 (
            .O(N__46084),
            .I(N__46081));
    LocalMux I__7052 (
            .O(N__46081),
            .I(\uart_pc.data_Auxce_0_5 ));
    CascadeMux I__7051 (
            .O(N__46078),
            .I(N__46070));
    InMux I__7050 (
            .O(N__46077),
            .I(N__46066));
    InMux I__7049 (
            .O(N__46076),
            .I(N__46057));
    InMux I__7048 (
            .O(N__46075),
            .I(N__46057));
    InMux I__7047 (
            .O(N__46074),
            .I(N__46057));
    InMux I__7046 (
            .O(N__46073),
            .I(N__46057));
    InMux I__7045 (
            .O(N__46070),
            .I(N__46052));
    InMux I__7044 (
            .O(N__46069),
            .I(N__46052));
    LocalMux I__7043 (
            .O(N__46066),
            .I(\uart_pc.un1_state_2_0 ));
    LocalMux I__7042 (
            .O(N__46057),
            .I(\uart_pc.un1_state_2_0 ));
    LocalMux I__7041 (
            .O(N__46052),
            .I(\uart_pc.un1_state_2_0 ));
    InMux I__7040 (
            .O(N__46045),
            .I(N__46042));
    LocalMux I__7039 (
            .O(N__46042),
            .I(N__46039));
    Span4Mux_h I__7038 (
            .O(N__46039),
            .I(N__46036));
    Odrv4 I__7037 (
            .O(N__46036),
            .I(\uart_pc.data_Auxce_0_6 ));
    InMux I__7036 (
            .O(N__46033),
            .I(N__46029));
    InMux I__7035 (
            .O(N__46032),
            .I(N__46026));
    LocalMux I__7034 (
            .O(N__46029),
            .I(\uart_pc.data_AuxZ0Z_6 ));
    LocalMux I__7033 (
            .O(N__46026),
            .I(\uart_pc.data_AuxZ0Z_6 ));
    SRMux I__7032 (
            .O(N__46021),
            .I(N__46018));
    LocalMux I__7031 (
            .O(N__46018),
            .I(N__46014));
    SRMux I__7030 (
            .O(N__46017),
            .I(N__46011));
    Span4Mux_h I__7029 (
            .O(N__46014),
            .I(N__46008));
    LocalMux I__7028 (
            .O(N__46011),
            .I(N__46003));
    Span4Mux_h I__7027 (
            .O(N__46008),
            .I(N__46003));
    Odrv4 I__7026 (
            .O(N__46003),
            .I(\uart_pc.state_RNIEAGSZ0Z_4 ));
    InMux I__7025 (
            .O(N__46000),
            .I(N__45996));
    InMux I__7024 (
            .O(N__45999),
            .I(N__45993));
    LocalMux I__7023 (
            .O(N__45996),
            .I(\uart_pc.data_AuxZ1Z_2 ));
    LocalMux I__7022 (
            .O(N__45993),
            .I(\uart_pc.data_AuxZ1Z_2 ));
    CascadeMux I__7021 (
            .O(N__45988),
            .I(\Commands_frame_decoder.state_ns_0_a3_0_1Z0Z_2_cascade_ ));
    InMux I__7020 (
            .O(N__45985),
            .I(N__45981));
    InMux I__7019 (
            .O(N__45984),
            .I(N__45976));
    LocalMux I__7018 (
            .O(N__45981),
            .I(N__45973));
    InMux I__7017 (
            .O(N__45980),
            .I(N__45968));
    InMux I__7016 (
            .O(N__45979),
            .I(N__45968));
    LocalMux I__7015 (
            .O(N__45976),
            .I(\Commands_frame_decoder.stateZ0Z_1 ));
    Odrv4 I__7014 (
            .O(N__45973),
            .I(\Commands_frame_decoder.stateZ0Z_1 ));
    LocalMux I__7013 (
            .O(N__45968),
            .I(\Commands_frame_decoder.stateZ0Z_1 ));
    InMux I__7012 (
            .O(N__45961),
            .I(N__45957));
    InMux I__7011 (
            .O(N__45960),
            .I(N__45954));
    LocalMux I__7010 (
            .O(N__45957),
            .I(N__45949));
    LocalMux I__7009 (
            .O(N__45954),
            .I(N__45949));
    Odrv12 I__7008 (
            .O(N__45949),
            .I(\Commands_frame_decoder.N_406 ));
    InMux I__7007 (
            .O(N__45946),
            .I(N__45942));
    InMux I__7006 (
            .O(N__45945),
            .I(N__45939));
    LocalMux I__7005 (
            .O(N__45942),
            .I(\uart_pc.data_AuxZ1Z_0 ));
    LocalMux I__7004 (
            .O(N__45939),
            .I(\uart_pc.data_AuxZ1Z_0 ));
    CascadeMux I__7003 (
            .O(N__45934),
            .I(N__45930));
    InMux I__7002 (
            .O(N__45933),
            .I(N__45927));
    InMux I__7001 (
            .O(N__45930),
            .I(N__45924));
    LocalMux I__7000 (
            .O(N__45927),
            .I(\uart_pc.data_AuxZ0Z_5 ));
    LocalMux I__6999 (
            .O(N__45924),
            .I(\uart_pc.data_AuxZ0Z_5 ));
    CascadeMux I__6998 (
            .O(N__45919),
            .I(N__45915));
    CascadeMux I__6997 (
            .O(N__45918),
            .I(N__45909));
    InMux I__6996 (
            .O(N__45915),
            .I(N__45898));
    InMux I__6995 (
            .O(N__45914),
            .I(N__45898));
    InMux I__6994 (
            .O(N__45913),
            .I(N__45898));
    InMux I__6993 (
            .O(N__45912),
            .I(N__45898));
    InMux I__6992 (
            .O(N__45909),
            .I(N__45891));
    InMux I__6991 (
            .O(N__45908),
            .I(N__45891));
    InMux I__6990 (
            .O(N__45907),
            .I(N__45891));
    LocalMux I__6989 (
            .O(N__45898),
            .I(\uart_pc.timer_Count_RNILR1B2Z0Z_2 ));
    LocalMux I__6988 (
            .O(N__45891),
            .I(\uart_pc.timer_Count_RNILR1B2Z0Z_2 ));
    CEMux I__6987 (
            .O(N__45886),
            .I(N__45883));
    LocalMux I__6986 (
            .O(N__45883),
            .I(N__45880));
    Span4Mux_v I__6985 (
            .O(N__45880),
            .I(N__45877));
    Odrv4 I__6984 (
            .O(N__45877),
            .I(\Commands_frame_decoder.source_CH4data_1_sqmuxa_0 ));
    InMux I__6983 (
            .O(N__45874),
            .I(N__45871));
    LocalMux I__6982 (
            .O(N__45871),
            .I(N__45867));
    InMux I__6981 (
            .O(N__45870),
            .I(N__45864));
    Span4Mux_h I__6980 (
            .O(N__45867),
            .I(N__45861));
    LocalMux I__6979 (
            .O(N__45864),
            .I(\uart_pc.N_126_li ));
    Odrv4 I__6978 (
            .O(N__45861),
            .I(\uart_pc.N_126_li ));
    InMux I__6977 (
            .O(N__45856),
            .I(N__45852));
    InMux I__6976 (
            .O(N__45855),
            .I(N__45849));
    LocalMux I__6975 (
            .O(N__45852),
            .I(N__45844));
    LocalMux I__6974 (
            .O(N__45849),
            .I(N__45844));
    Span4Mux_h I__6973 (
            .O(N__45844),
            .I(N__45837));
    InMux I__6972 (
            .O(N__45843),
            .I(N__45834));
    InMux I__6971 (
            .O(N__45842),
            .I(N__45831));
    InMux I__6970 (
            .O(N__45841),
            .I(N__45826));
    InMux I__6969 (
            .O(N__45840),
            .I(N__45826));
    Sp12to4 I__6968 (
            .O(N__45837),
            .I(N__45821));
    LocalMux I__6967 (
            .O(N__45834),
            .I(N__45821));
    LocalMux I__6966 (
            .O(N__45831),
            .I(N__45816));
    LocalMux I__6965 (
            .O(N__45826),
            .I(N__45816));
    Odrv12 I__6964 (
            .O(N__45821),
            .I(\uart_pc.stateZ0Z_4 ));
    Odrv4 I__6963 (
            .O(N__45816),
            .I(\uart_pc.stateZ0Z_4 ));
    CascadeMux I__6962 (
            .O(N__45811),
            .I(N__45808));
    InMux I__6961 (
            .O(N__45808),
            .I(N__45805));
    LocalMux I__6960 (
            .O(N__45805),
            .I(N__45802));
    Span4Mux_h I__6959 (
            .O(N__45802),
            .I(N__45799));
    Odrv4 I__6958 (
            .O(N__45799),
            .I(\uart_pc.un1_state_2_0_a3_0 ));
    InMux I__6957 (
            .O(N__45796),
            .I(N__45791));
    InMux I__6956 (
            .O(N__45795),
            .I(N__45786));
    CascadeMux I__6955 (
            .O(N__45794),
            .I(N__45782));
    LocalMux I__6954 (
            .O(N__45791),
            .I(N__45777));
    InMux I__6953 (
            .O(N__45790),
            .I(N__45772));
    InMux I__6952 (
            .O(N__45789),
            .I(N__45772));
    LocalMux I__6951 (
            .O(N__45786),
            .I(N__45769));
    InMux I__6950 (
            .O(N__45785),
            .I(N__45766));
    InMux I__6949 (
            .O(N__45782),
            .I(N__45759));
    InMux I__6948 (
            .O(N__45781),
            .I(N__45759));
    InMux I__6947 (
            .O(N__45780),
            .I(N__45759));
    Odrv12 I__6946 (
            .O(N__45777),
            .I(\uart_pc.stateZ0Z_3 ));
    LocalMux I__6945 (
            .O(N__45772),
            .I(\uart_pc.stateZ0Z_3 ));
    Odrv4 I__6944 (
            .O(N__45769),
            .I(\uart_pc.stateZ0Z_3 ));
    LocalMux I__6943 (
            .O(N__45766),
            .I(\uart_pc.stateZ0Z_3 ));
    LocalMux I__6942 (
            .O(N__45759),
            .I(\uart_pc.stateZ0Z_3 ));
    CascadeMux I__6941 (
            .O(N__45748),
            .I(\uart_pc.un1_state_2_0_cascade_ ));
    InMux I__6940 (
            .O(N__45745),
            .I(N__45742));
    LocalMux I__6939 (
            .O(N__45742),
            .I(\uart_pc.data_Auxce_0_0_0 ));
    InMux I__6938 (
            .O(N__45739),
            .I(N__45736));
    LocalMux I__6937 (
            .O(N__45736),
            .I(\uart_pc.data_Auxce_0_1 ));
    InMux I__6936 (
            .O(N__45733),
            .I(N__45730));
    LocalMux I__6935 (
            .O(N__45730),
            .I(\uart_pc.data_Auxce_0_0_2 ));
    InMux I__6934 (
            .O(N__45727),
            .I(N__45724));
    LocalMux I__6933 (
            .O(N__45724),
            .I(\uart_pc.data_Auxce_0_3 ));
    CascadeMux I__6932 (
            .O(N__45721),
            .I(N__45718));
    InMux I__6931 (
            .O(N__45718),
            .I(N__45715));
    LocalMux I__6930 (
            .O(N__45715),
            .I(N__45711));
    InMux I__6929 (
            .O(N__45714),
            .I(N__45708));
    Odrv4 I__6928 (
            .O(N__45711),
            .I(\uart_pc.data_AuxZ0Z_3 ));
    LocalMux I__6927 (
            .O(N__45708),
            .I(\uart_pc.data_AuxZ0Z_3 ));
    InMux I__6926 (
            .O(N__45703),
            .I(N__45700));
    LocalMux I__6925 (
            .O(N__45700),
            .I(\uart_pc.data_Auxce_0_0_4 ));
    InMux I__6924 (
            .O(N__45697),
            .I(N__45693));
    InMux I__6923 (
            .O(N__45696),
            .I(N__45690));
    LocalMux I__6922 (
            .O(N__45693),
            .I(\uart_pc.data_AuxZ0Z_4 ));
    LocalMux I__6921 (
            .O(N__45690),
            .I(\uart_pc.data_AuxZ0Z_4 ));
    InMux I__6920 (
            .O(N__45685),
            .I(N__45682));
    LocalMux I__6919 (
            .O(N__45682),
            .I(N__45678));
    InMux I__6918 (
            .O(N__45681),
            .I(N__45675));
    Span4Mux_s3_h I__6917 (
            .O(N__45678),
            .I(N__45672));
    LocalMux I__6916 (
            .O(N__45675),
            .I(N__45669));
    Span4Mux_h I__6915 (
            .O(N__45672),
            .I(N__45666));
    Span4Mux_v I__6914 (
            .O(N__45669),
            .I(N__45663));
    Span4Mux_h I__6913 (
            .O(N__45666),
            .I(N__45660));
    Span4Mux_h I__6912 (
            .O(N__45663),
            .I(N__45657));
    Span4Mux_h I__6911 (
            .O(N__45660),
            .I(N__45654));
    Span4Mux_h I__6910 (
            .O(N__45657),
            .I(N__45651));
    Odrv4 I__6909 (
            .O(N__45654),
            .I(xy_kp_3));
    Odrv4 I__6908 (
            .O(N__45651),
            .I(xy_kp_3));
    InMux I__6907 (
            .O(N__45646),
            .I(N__45642));
    InMux I__6906 (
            .O(N__45645),
            .I(N__45639));
    LocalMux I__6905 (
            .O(N__45642),
            .I(N__45636));
    LocalMux I__6904 (
            .O(N__45639),
            .I(N__45633));
    Span4Mux_s2_h I__6903 (
            .O(N__45636),
            .I(N__45630));
    Span12Mux_v I__6902 (
            .O(N__45633),
            .I(N__45627));
    Span4Mux_h I__6901 (
            .O(N__45630),
            .I(N__45624));
    Span12Mux_h I__6900 (
            .O(N__45627),
            .I(N__45621));
    Span4Mux_h I__6899 (
            .O(N__45624),
            .I(N__45618));
    Odrv12 I__6898 (
            .O(N__45621),
            .I(xy_kp_5));
    Odrv4 I__6897 (
            .O(N__45618),
            .I(xy_kp_5));
    InMux I__6896 (
            .O(N__45613),
            .I(N__45610));
    LocalMux I__6895 (
            .O(N__45610),
            .I(N__45607));
    Span4Mux_s2_h I__6894 (
            .O(N__45607),
            .I(N__45603));
    InMux I__6893 (
            .O(N__45606),
            .I(N__45600));
    Span4Mux_v I__6892 (
            .O(N__45603),
            .I(N__45597));
    LocalMux I__6891 (
            .O(N__45600),
            .I(N__45594));
    Sp12to4 I__6890 (
            .O(N__45597),
            .I(N__45591));
    Span4Mux_v I__6889 (
            .O(N__45594),
            .I(N__45588));
    Span12Mux_h I__6888 (
            .O(N__45591),
            .I(N__45585));
    Sp12to4 I__6887 (
            .O(N__45588),
            .I(N__45582));
    Odrv12 I__6886 (
            .O(N__45585),
            .I(xy_kp_6));
    Odrv12 I__6885 (
            .O(N__45582),
            .I(xy_kp_6));
    InMux I__6884 (
            .O(N__45577),
            .I(N__45574));
    LocalMux I__6883 (
            .O(N__45574),
            .I(N__45571));
    Span4Mux_s3_h I__6882 (
            .O(N__45571),
            .I(N__45567));
    InMux I__6881 (
            .O(N__45570),
            .I(N__45564));
    Span4Mux_h I__6880 (
            .O(N__45567),
            .I(N__45561));
    LocalMux I__6879 (
            .O(N__45564),
            .I(N__45558));
    Span4Mux_h I__6878 (
            .O(N__45561),
            .I(N__45555));
    Span4Mux_v I__6877 (
            .O(N__45558),
            .I(N__45552));
    Span4Mux_h I__6876 (
            .O(N__45555),
            .I(N__45549));
    Sp12to4 I__6875 (
            .O(N__45552),
            .I(N__45546));
    Odrv4 I__6874 (
            .O(N__45549),
            .I(xy_kp_7));
    Odrv12 I__6873 (
            .O(N__45546),
            .I(xy_kp_7));
    CascadeMux I__6872 (
            .O(N__45541),
            .I(N__45538));
    InMux I__6871 (
            .O(N__45538),
            .I(N__45533));
    InMux I__6870 (
            .O(N__45537),
            .I(N__45530));
    InMux I__6869 (
            .O(N__45536),
            .I(N__45527));
    LocalMux I__6868 (
            .O(N__45533),
            .I(\uart_pc.N_152 ));
    LocalMux I__6867 (
            .O(N__45530),
            .I(\uart_pc.N_152 ));
    LocalMux I__6866 (
            .O(N__45527),
            .I(\uart_pc.N_152 ));
    InMux I__6865 (
            .O(N__45520),
            .I(N__45517));
    LocalMux I__6864 (
            .O(N__45517),
            .I(N__45513));
    CascadeMux I__6863 (
            .O(N__45516),
            .I(N__45510));
    Span4Mux_v I__6862 (
            .O(N__45513),
            .I(N__45507));
    InMux I__6861 (
            .O(N__45510),
            .I(N__45504));
    Odrv4 I__6860 (
            .O(N__45507),
            .I(\uart_pc.data_AuxZ0Z_7 ));
    LocalMux I__6859 (
            .O(N__45504),
            .I(\uart_pc.data_AuxZ0Z_7 ));
    CEMux I__6858 (
            .O(N__45499),
            .I(N__45496));
    LocalMux I__6857 (
            .O(N__45496),
            .I(N__45492));
    CEMux I__6856 (
            .O(N__45495),
            .I(N__45489));
    Span4Mux_v I__6855 (
            .O(N__45492),
            .I(N__45484));
    LocalMux I__6854 (
            .O(N__45489),
            .I(N__45484));
    Span4Mux_v I__6853 (
            .O(N__45484),
            .I(N__45481));
    Span4Mux_h I__6852 (
            .O(N__45481),
            .I(N__45478));
    Odrv4 I__6851 (
            .O(N__45478),
            .I(\Commands_frame_decoder.un1_sink_data_valid_2_0_0 ));
    InMux I__6850 (
            .O(N__45475),
            .I(N__45472));
    LocalMux I__6849 (
            .O(N__45472),
            .I(N__45469));
    Sp12to4 I__6848 (
            .O(N__45469),
            .I(N__45466));
    Odrv12 I__6847 (
            .O(N__45466),
            .I(\Commands_frame_decoder.source_offset4data_1_sqmuxa ));
    CascadeMux I__6846 (
            .O(N__45463),
            .I(\Commands_frame_decoder.source_offset4data_1_sqmuxa_cascade_ ));
    CEMux I__6845 (
            .O(N__45460),
            .I(N__45457));
    LocalMux I__6844 (
            .O(N__45457),
            .I(N__45454));
    Odrv12 I__6843 (
            .O(N__45454),
            .I(\Commands_frame_decoder.source_offset4data_1_sqmuxa_0 ));
    CascadeMux I__6842 (
            .O(N__45451),
            .I(N__45448));
    InMux I__6841 (
            .O(N__45448),
            .I(N__45445));
    LocalMux I__6840 (
            .O(N__45445),
            .I(N__45442));
    Odrv4 I__6839 (
            .O(N__45442),
            .I(frame_decoder_OFF4data_1));
    CascadeMux I__6838 (
            .O(N__45439),
            .I(N__45436));
    InMux I__6837 (
            .O(N__45436),
            .I(N__45433));
    LocalMux I__6836 (
            .O(N__45433),
            .I(N__45430));
    Odrv4 I__6835 (
            .O(N__45430),
            .I(frame_decoder_OFF4data_2));
    CascadeMux I__6834 (
            .O(N__45427),
            .I(N__45424));
    InMux I__6833 (
            .O(N__45424),
            .I(N__45421));
    LocalMux I__6832 (
            .O(N__45421),
            .I(N__45418));
    Odrv4 I__6831 (
            .O(N__45418),
            .I(frame_decoder_OFF4data_3));
    CascadeMux I__6830 (
            .O(N__45415),
            .I(N__45412));
    InMux I__6829 (
            .O(N__45412),
            .I(N__45409));
    LocalMux I__6828 (
            .O(N__45409),
            .I(N__45406));
    Odrv4 I__6827 (
            .O(N__45406),
            .I(frame_decoder_OFF4data_4));
    CascadeMux I__6826 (
            .O(N__45403),
            .I(N__45400));
    InMux I__6825 (
            .O(N__45400),
            .I(N__45397));
    LocalMux I__6824 (
            .O(N__45397),
            .I(N__45394));
    Odrv4 I__6823 (
            .O(N__45394),
            .I(frame_decoder_OFF4data_5));
    CascadeMux I__6822 (
            .O(N__45391),
            .I(N__45388));
    InMux I__6821 (
            .O(N__45388),
            .I(N__45385));
    LocalMux I__6820 (
            .O(N__45385),
            .I(N__45382));
    Odrv4 I__6819 (
            .O(N__45382),
            .I(frame_decoder_OFF4data_6));
    InMux I__6818 (
            .O(N__45379),
            .I(N__45376));
    LocalMux I__6817 (
            .O(N__45376),
            .I(N__45372));
    InMux I__6816 (
            .O(N__45375),
            .I(N__45369));
    Span4Mux_s3_h I__6815 (
            .O(N__45372),
            .I(N__45366));
    LocalMux I__6814 (
            .O(N__45369),
            .I(N__45363));
    Span4Mux_h I__6813 (
            .O(N__45366),
            .I(N__45360));
    Span4Mux_s2_h I__6812 (
            .O(N__45363),
            .I(N__45357));
    Span4Mux_h I__6811 (
            .O(N__45360),
            .I(N__45354));
    Span4Mux_h I__6810 (
            .O(N__45357),
            .I(N__45351));
    Span4Mux_h I__6809 (
            .O(N__45354),
            .I(N__45348));
    Span4Mux_h I__6808 (
            .O(N__45351),
            .I(N__45345));
    Odrv4 I__6807 (
            .O(N__45348),
            .I(xy_kp_0));
    Odrv4 I__6806 (
            .O(N__45345),
            .I(xy_kp_0));
    InMux I__6805 (
            .O(N__45340),
            .I(N__45336));
    InMux I__6804 (
            .O(N__45339),
            .I(N__45333));
    LocalMux I__6803 (
            .O(N__45336),
            .I(N__45330));
    LocalMux I__6802 (
            .O(N__45333),
            .I(N__45327));
    Span4Mux_s1_h I__6801 (
            .O(N__45330),
            .I(N__45324));
    Span12Mux_s4_h I__6800 (
            .O(N__45327),
            .I(N__45321));
    Span4Mux_h I__6799 (
            .O(N__45324),
            .I(N__45318));
    Span12Mux_h I__6798 (
            .O(N__45321),
            .I(N__45315));
    Span4Mux_h I__6797 (
            .O(N__45318),
            .I(N__45312));
    Odrv12 I__6796 (
            .O(N__45315),
            .I(xy_kp_1));
    Odrv4 I__6795 (
            .O(N__45312),
            .I(xy_kp_1));
    InMux I__6794 (
            .O(N__45307),
            .I(N__45304));
    LocalMux I__6793 (
            .O(N__45304),
            .I(N__45301));
    Span4Mux_s3_h I__6792 (
            .O(N__45301),
            .I(N__45298));
    Span4Mux_h I__6791 (
            .O(N__45298),
            .I(N__45294));
    InMux I__6790 (
            .O(N__45297),
            .I(N__45291));
    Span4Mux_h I__6789 (
            .O(N__45294),
            .I(N__45288));
    LocalMux I__6788 (
            .O(N__45291),
            .I(N__45285));
    Span4Mux_h I__6787 (
            .O(N__45288),
            .I(N__45282));
    Span12Mux_s9_h I__6786 (
            .O(N__45285),
            .I(N__45279));
    Odrv4 I__6785 (
            .O(N__45282),
            .I(xy_kp_2));
    Odrv12 I__6784 (
            .O(N__45279),
            .I(xy_kp_2));
    CascadeMux I__6783 (
            .O(N__45274),
            .I(\uart_drone.N_126_li_cascade_ ));
    CascadeMux I__6782 (
            .O(N__45271),
            .I(\uart_drone.N_143_cascade_ ));
    InMux I__6781 (
            .O(N__45268),
            .I(N__45263));
    CascadeMux I__6780 (
            .O(N__45267),
            .I(N__45260));
    InMux I__6779 (
            .O(N__45266),
            .I(N__45256));
    LocalMux I__6778 (
            .O(N__45263),
            .I(N__45253));
    InMux I__6777 (
            .O(N__45260),
            .I(N__45248));
    InMux I__6776 (
            .O(N__45259),
            .I(N__45248));
    LocalMux I__6775 (
            .O(N__45256),
            .I(\scaler_4.un2_source_data_0 ));
    Odrv12 I__6774 (
            .O(N__45253),
            .I(\scaler_4.un2_source_data_0 ));
    LocalMux I__6773 (
            .O(N__45248),
            .I(\scaler_4.un2_source_data_0 ));
    InMux I__6772 (
            .O(N__45241),
            .I(N__45238));
    LocalMux I__6771 (
            .O(N__45238),
            .I(N__45232));
    InMux I__6770 (
            .O(N__45237),
            .I(N__45229));
    InMux I__6769 (
            .O(N__45236),
            .I(N__45226));
    InMux I__6768 (
            .O(N__45235),
            .I(N__45223));
    Odrv12 I__6767 (
            .O(N__45232),
            .I(frame_decoder_CH4data_0));
    LocalMux I__6766 (
            .O(N__45229),
            .I(frame_decoder_CH4data_0));
    LocalMux I__6765 (
            .O(N__45226),
            .I(frame_decoder_CH4data_0));
    LocalMux I__6764 (
            .O(N__45223),
            .I(frame_decoder_CH4data_0));
    CascadeMux I__6763 (
            .O(N__45214),
            .I(N__45211));
    InMux I__6762 (
            .O(N__45211),
            .I(N__45208));
    LocalMux I__6761 (
            .O(N__45208),
            .I(N__45205));
    Odrv4 I__6760 (
            .O(N__45205),
            .I(\scaler_4.un2_source_data_0_cry_1_c_RNOZ0 ));
    IoInMux I__6759 (
            .O(N__45202),
            .I(N__45199));
    LocalMux I__6758 (
            .O(N__45199),
            .I(N__45196));
    Span4Mux_s2_v I__6757 (
            .O(N__45196),
            .I(N__45193));
    Sp12to4 I__6756 (
            .O(N__45193),
            .I(N__45190));
    Span12Mux_h I__6755 (
            .O(N__45190),
            .I(N__45187));
    Odrv12 I__6754 (
            .O(N__45187),
            .I(\pid_alt.N_933_0 ));
    CascadeMux I__6753 (
            .O(N__45184),
            .I(N__45178));
    InMux I__6752 (
            .O(N__45183),
            .I(N__45175));
    InMux I__6751 (
            .O(N__45182),
            .I(N__45172));
    InMux I__6750 (
            .O(N__45181),
            .I(N__45169));
    InMux I__6749 (
            .O(N__45178),
            .I(N__45166));
    LocalMux I__6748 (
            .O(N__45175),
            .I(N__45163));
    LocalMux I__6747 (
            .O(N__45172),
            .I(N__45156));
    LocalMux I__6746 (
            .O(N__45169),
            .I(N__45156));
    LocalMux I__6745 (
            .O(N__45166),
            .I(N__45156));
    Odrv4 I__6744 (
            .O(N__45163),
            .I(frame_decoder_OFF4data_0));
    Odrv4 I__6743 (
            .O(N__45156),
            .I(frame_decoder_OFF4data_0));
    InMux I__6742 (
            .O(N__45151),
            .I(N__45148));
    LocalMux I__6741 (
            .O(N__45148),
            .I(N__45145));
    Span4Mux_h I__6740 (
            .O(N__45145),
            .I(N__45142));
    Span4Mux_h I__6739 (
            .O(N__45142),
            .I(N__45139));
    Odrv4 I__6738 (
            .O(N__45139),
            .I(\ppm_encoder_1.un1_throttle_cry_6_THRU_CO ));
    InMux I__6737 (
            .O(N__45136),
            .I(N__45133));
    LocalMux I__6736 (
            .O(N__45133),
            .I(N__45129));
    CascadeMux I__6735 (
            .O(N__45132),
            .I(N__45125));
    Span4Mux_v I__6734 (
            .O(N__45129),
            .I(N__45122));
    InMux I__6733 (
            .O(N__45128),
            .I(N__45119));
    InMux I__6732 (
            .O(N__45125),
            .I(N__45116));
    Span4Mux_h I__6731 (
            .O(N__45122),
            .I(N__45111));
    LocalMux I__6730 (
            .O(N__45119),
            .I(N__45111));
    LocalMux I__6729 (
            .O(N__45116),
            .I(throttle_order_7));
    Odrv4 I__6728 (
            .O(N__45111),
            .I(throttle_order_7));
    InMux I__6727 (
            .O(N__45106),
            .I(N__45103));
    LocalMux I__6726 (
            .O(N__45103),
            .I(N__45099));
    CascadeMux I__6725 (
            .O(N__45102),
            .I(N__45096));
    Span4Mux_h I__6724 (
            .O(N__45099),
            .I(N__45093));
    InMux I__6723 (
            .O(N__45096),
            .I(N__45089));
    Span4Mux_h I__6722 (
            .O(N__45093),
            .I(N__45086));
    InMux I__6721 (
            .O(N__45092),
            .I(N__45083));
    LocalMux I__6720 (
            .O(N__45089),
            .I(throttle_order_8));
    Odrv4 I__6719 (
            .O(N__45086),
            .I(throttle_order_8));
    LocalMux I__6718 (
            .O(N__45083),
            .I(throttle_order_8));
    InMux I__6717 (
            .O(N__45076),
            .I(N__45073));
    LocalMux I__6716 (
            .O(N__45073),
            .I(N__45070));
    Span4Mux_v I__6715 (
            .O(N__45070),
            .I(N__45067));
    Span4Mux_h I__6714 (
            .O(N__45067),
            .I(N__45064));
    Odrv4 I__6713 (
            .O(N__45064),
            .I(\ppm_encoder_1.un1_throttle_cry_7_THRU_CO ));
    InMux I__6712 (
            .O(N__45061),
            .I(N__45056));
    InMux I__6711 (
            .O(N__45060),
            .I(N__45053));
    CascadeMux I__6710 (
            .O(N__45059),
            .I(N__45050));
    LocalMux I__6709 (
            .O(N__45056),
            .I(N__45047));
    LocalMux I__6708 (
            .O(N__45053),
            .I(N__45044));
    InMux I__6707 (
            .O(N__45050),
            .I(N__45041));
    Span4Mux_h I__6706 (
            .O(N__45047),
            .I(N__45038));
    Span4Mux_h I__6705 (
            .O(N__45044),
            .I(N__45035));
    LocalMux I__6704 (
            .O(N__45041),
            .I(\ppm_encoder_1.throttleZ0Z_8 ));
    Odrv4 I__6703 (
            .O(N__45038),
            .I(\ppm_encoder_1.throttleZ0Z_8 ));
    Odrv4 I__6702 (
            .O(N__45035),
            .I(\ppm_encoder_1.throttleZ0Z_8 ));
    InMux I__6701 (
            .O(N__45028),
            .I(N__45025));
    LocalMux I__6700 (
            .O(N__45025),
            .I(N__45022));
    Span4Mux_h I__6699 (
            .O(N__45022),
            .I(N__45018));
    InMux I__6698 (
            .O(N__45021),
            .I(N__45014));
    Span4Mux_h I__6697 (
            .O(N__45018),
            .I(N__45011));
    InMux I__6696 (
            .O(N__45017),
            .I(N__45008));
    LocalMux I__6695 (
            .O(N__45014),
            .I(throttle_order_9));
    Odrv4 I__6694 (
            .O(N__45011),
            .I(throttle_order_9));
    LocalMux I__6693 (
            .O(N__45008),
            .I(throttle_order_9));
    InMux I__6692 (
            .O(N__45001),
            .I(N__44998));
    LocalMux I__6691 (
            .O(N__44998),
            .I(N__44995));
    Span4Mux_v I__6690 (
            .O(N__44995),
            .I(N__44992));
    Span4Mux_h I__6689 (
            .O(N__44992),
            .I(N__44989));
    Odrv4 I__6688 (
            .O(N__44989),
            .I(\ppm_encoder_1.un1_throttle_cry_8_THRU_CO ));
    CascadeMux I__6687 (
            .O(N__44986),
            .I(N__44983));
    InMux I__6686 (
            .O(N__44983),
            .I(N__44979));
    InMux I__6685 (
            .O(N__44982),
            .I(N__44975));
    LocalMux I__6684 (
            .O(N__44979),
            .I(N__44972));
    InMux I__6683 (
            .O(N__44978),
            .I(N__44969));
    LocalMux I__6682 (
            .O(N__44975),
            .I(N__44966));
    Span4Mux_h I__6681 (
            .O(N__44972),
            .I(N__44963));
    LocalMux I__6680 (
            .O(N__44969),
            .I(\ppm_encoder_1.throttleZ0Z_9 ));
    Odrv4 I__6679 (
            .O(N__44966),
            .I(\ppm_encoder_1.throttleZ0Z_9 ));
    Odrv4 I__6678 (
            .O(N__44963),
            .I(\ppm_encoder_1.throttleZ0Z_9 ));
    InMux I__6677 (
            .O(N__44956),
            .I(N__44952));
    InMux I__6676 (
            .O(N__44955),
            .I(N__44949));
    LocalMux I__6675 (
            .O(N__44952),
            .I(N__44946));
    LocalMux I__6674 (
            .O(N__44949),
            .I(\ppm_encoder_1.aileronZ0Z_6 ));
    Odrv4 I__6673 (
            .O(N__44946),
            .I(\ppm_encoder_1.aileronZ0Z_6 ));
    CascadeMux I__6672 (
            .O(N__44941),
            .I(N__44938));
    InMux I__6671 (
            .O(N__44938),
            .I(N__44934));
    InMux I__6670 (
            .O(N__44937),
            .I(N__44931));
    LocalMux I__6669 (
            .O(N__44934),
            .I(N__44928));
    LocalMux I__6668 (
            .O(N__44931),
            .I(\ppm_encoder_1.throttleZ0Z_6 ));
    Odrv12 I__6667 (
            .O(N__44928),
            .I(\ppm_encoder_1.throttleZ0Z_6 ));
    InMux I__6666 (
            .O(N__44923),
            .I(N__44916));
    InMux I__6665 (
            .O(N__44922),
            .I(N__44916));
    InMux I__6664 (
            .O(N__44921),
            .I(N__44913));
    LocalMux I__6663 (
            .O(N__44916),
            .I(N__44908));
    LocalMux I__6662 (
            .O(N__44913),
            .I(N__44908));
    Span4Mux_v I__6661 (
            .O(N__44908),
            .I(N__44902));
    InMux I__6660 (
            .O(N__44907),
            .I(N__44899));
    InMux I__6659 (
            .O(N__44906),
            .I(N__44892));
    InMux I__6658 (
            .O(N__44905),
            .I(N__44892));
    Span4Mux_h I__6657 (
            .O(N__44902),
            .I(N__44886));
    LocalMux I__6656 (
            .O(N__44899),
            .I(N__44886));
    InMux I__6655 (
            .O(N__44898),
            .I(N__44881));
    InMux I__6654 (
            .O(N__44897),
            .I(N__44881));
    LocalMux I__6653 (
            .O(N__44892),
            .I(N__44878));
    InMux I__6652 (
            .O(N__44891),
            .I(N__44875));
    Odrv4 I__6651 (
            .O(N__44886),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ));
    LocalMux I__6650 (
            .O(N__44881),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ));
    Odrv4 I__6649 (
            .O(N__44878),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ));
    LocalMux I__6648 (
            .O(N__44875),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ));
    InMux I__6647 (
            .O(N__44866),
            .I(N__44862));
    CascadeMux I__6646 (
            .O(N__44865),
            .I(N__44859));
    LocalMux I__6645 (
            .O(N__44862),
            .I(N__44856));
    InMux I__6644 (
            .O(N__44859),
            .I(N__44853));
    Span4Mux_h I__6643 (
            .O(N__44856),
            .I(N__44848));
    LocalMux I__6642 (
            .O(N__44853),
            .I(N__44845));
    InMux I__6641 (
            .O(N__44852),
            .I(N__44842));
    CascadeMux I__6640 (
            .O(N__44851),
            .I(N__44839));
    Span4Mux_v I__6639 (
            .O(N__44848),
            .I(N__44836));
    Span4Mux_s1_v I__6638 (
            .O(N__44845),
            .I(N__44833));
    LocalMux I__6637 (
            .O(N__44842),
            .I(N__44830));
    InMux I__6636 (
            .O(N__44839),
            .I(N__44827));
    Odrv4 I__6635 (
            .O(N__44836),
            .I(\ppm_encoder_1.init_pulsesZ0Z_3 ));
    Odrv4 I__6634 (
            .O(N__44833),
            .I(\ppm_encoder_1.init_pulsesZ0Z_3 ));
    Odrv12 I__6633 (
            .O(N__44830),
            .I(\ppm_encoder_1.init_pulsesZ0Z_3 ));
    LocalMux I__6632 (
            .O(N__44827),
            .I(\ppm_encoder_1.init_pulsesZ0Z_3 ));
    InMux I__6631 (
            .O(N__44818),
            .I(N__44815));
    LocalMux I__6630 (
            .O(N__44815),
            .I(N__44811));
    CascadeMux I__6629 (
            .O(N__44814),
            .I(N__44808));
    Span4Mux_h I__6628 (
            .O(N__44811),
            .I(N__44805));
    InMux I__6627 (
            .O(N__44808),
            .I(N__44801));
    Span4Mux_h I__6626 (
            .O(N__44805),
            .I(N__44798));
    InMux I__6625 (
            .O(N__44804),
            .I(N__44795));
    LocalMux I__6624 (
            .O(N__44801),
            .I(\ppm_encoder_1.aileronZ0Z_8 ));
    Odrv4 I__6623 (
            .O(N__44798),
            .I(\ppm_encoder_1.aileronZ0Z_8 ));
    LocalMux I__6622 (
            .O(N__44795),
            .I(\ppm_encoder_1.aileronZ0Z_8 ));
    CascadeMux I__6621 (
            .O(N__44788),
            .I(N__44785));
    InMux I__6620 (
            .O(N__44785),
            .I(N__44782));
    LocalMux I__6619 (
            .O(N__44782),
            .I(N__44779));
    Span4Mux_v I__6618 (
            .O(N__44779),
            .I(N__44775));
    InMux I__6617 (
            .O(N__44778),
            .I(N__44771));
    Span4Mux_h I__6616 (
            .O(N__44775),
            .I(N__44768));
    InMux I__6615 (
            .O(N__44774),
            .I(N__44765));
    LocalMux I__6614 (
            .O(N__44771),
            .I(\ppm_encoder_1.elevatorZ0Z_8 ));
    Odrv4 I__6613 (
            .O(N__44768),
            .I(\ppm_encoder_1.elevatorZ0Z_8 ));
    LocalMux I__6612 (
            .O(N__44765),
            .I(\ppm_encoder_1.elevatorZ0Z_8 ));
    InMux I__6611 (
            .O(N__44758),
            .I(N__44755));
    LocalMux I__6610 (
            .O(N__44755),
            .I(N__44750));
    InMux I__6609 (
            .O(N__44754),
            .I(N__44747));
    InMux I__6608 (
            .O(N__44753),
            .I(N__44744));
    Span4Mux_v I__6607 (
            .O(N__44750),
            .I(N__44741));
    LocalMux I__6606 (
            .O(N__44747),
            .I(\ppm_encoder_1.aileronZ0Z_9 ));
    LocalMux I__6605 (
            .O(N__44744),
            .I(\ppm_encoder_1.aileronZ0Z_9 ));
    Odrv4 I__6604 (
            .O(N__44741),
            .I(\ppm_encoder_1.aileronZ0Z_9 ));
    CascadeMux I__6603 (
            .O(N__44734),
            .I(N__44731));
    InMux I__6602 (
            .O(N__44731),
            .I(N__44728));
    LocalMux I__6601 (
            .O(N__44728),
            .I(N__44725));
    Span4Mux_h I__6600 (
            .O(N__44725),
            .I(N__44722));
    Span4Mux_v I__6599 (
            .O(N__44722),
            .I(N__44719));
    Odrv4 I__6598 (
            .O(N__44719),
            .I(\ppm_encoder_1.pulses2count_9_i_1_9 ));
    CascadeMux I__6597 (
            .O(N__44716),
            .I(N__44713));
    InMux I__6596 (
            .O(N__44713),
            .I(N__44710));
    LocalMux I__6595 (
            .O(N__44710),
            .I(N__44705));
    InMux I__6594 (
            .O(N__44709),
            .I(N__44700));
    InMux I__6593 (
            .O(N__44708),
            .I(N__44700));
    Span4Mux_v I__6592 (
            .O(N__44705),
            .I(N__44697));
    LocalMux I__6591 (
            .O(N__44700),
            .I(\ppm_encoder_1.elevatorZ0Z_9 ));
    Odrv4 I__6590 (
            .O(N__44697),
            .I(\ppm_encoder_1.elevatorZ0Z_9 ));
    InMux I__6589 (
            .O(N__44692),
            .I(N__44689));
    LocalMux I__6588 (
            .O(N__44689),
            .I(\ppm_encoder_1.N_293 ));
    InMux I__6587 (
            .O(N__44686),
            .I(N__44683));
    LocalMux I__6586 (
            .O(N__44683),
            .I(N__44675));
    InMux I__6585 (
            .O(N__44682),
            .I(N__44672));
    InMux I__6584 (
            .O(N__44681),
            .I(N__44669));
    InMux I__6583 (
            .O(N__44680),
            .I(N__44665));
    InMux I__6582 (
            .O(N__44679),
            .I(N__44662));
    InMux I__6581 (
            .O(N__44678),
            .I(N__44659));
    Span4Mux_h I__6580 (
            .O(N__44675),
            .I(N__44656));
    LocalMux I__6579 (
            .O(N__44672),
            .I(N__44651));
    LocalMux I__6578 (
            .O(N__44669),
            .I(N__44651));
    CascadeMux I__6577 (
            .O(N__44668),
            .I(N__44645));
    LocalMux I__6576 (
            .O(N__44665),
            .I(N__44638));
    LocalMux I__6575 (
            .O(N__44662),
            .I(N__44638));
    LocalMux I__6574 (
            .O(N__44659),
            .I(N__44638));
    Span4Mux_h I__6573 (
            .O(N__44656),
            .I(N__44635));
    Span4Mux_h I__6572 (
            .O(N__44651),
            .I(N__44632));
    InMux I__6571 (
            .O(N__44650),
            .I(N__44627));
    InMux I__6570 (
            .O(N__44649),
            .I(N__44627));
    InMux I__6569 (
            .O(N__44648),
            .I(N__44622));
    InMux I__6568 (
            .O(N__44645),
            .I(N__44622));
    Span4Mux_h I__6567 (
            .O(N__44638),
            .I(N__44619));
    Odrv4 I__6566 (
            .O(N__44635),
            .I(\ppm_encoder_1.N_507 ));
    Odrv4 I__6565 (
            .O(N__44632),
            .I(\ppm_encoder_1.N_507 ));
    LocalMux I__6564 (
            .O(N__44627),
            .I(\ppm_encoder_1.N_507 ));
    LocalMux I__6563 (
            .O(N__44622),
            .I(\ppm_encoder_1.N_507 ));
    Odrv4 I__6562 (
            .O(N__44619),
            .I(\ppm_encoder_1.N_507 ));
    InMux I__6561 (
            .O(N__44608),
            .I(N__44604));
    InMux I__6560 (
            .O(N__44607),
            .I(N__44601));
    LocalMux I__6559 (
            .O(N__44604),
            .I(N__44598));
    LocalMux I__6558 (
            .O(N__44601),
            .I(N__44590));
    Span4Mux_v I__6557 (
            .O(N__44598),
            .I(N__44587));
    InMux I__6556 (
            .O(N__44597),
            .I(N__44584));
    InMux I__6555 (
            .O(N__44596),
            .I(N__44581));
    InMux I__6554 (
            .O(N__44595),
            .I(N__44578));
    InMux I__6553 (
            .O(N__44594),
            .I(N__44575));
    InMux I__6552 (
            .O(N__44593),
            .I(N__44567));
    Span4Mux_h I__6551 (
            .O(N__44590),
            .I(N__44564));
    Span4Mux_h I__6550 (
            .O(N__44587),
            .I(N__44559));
    LocalMux I__6549 (
            .O(N__44584),
            .I(N__44559));
    LocalMux I__6548 (
            .O(N__44581),
            .I(N__44552));
    LocalMux I__6547 (
            .O(N__44578),
            .I(N__44552));
    LocalMux I__6546 (
            .O(N__44575),
            .I(N__44552));
    InMux I__6545 (
            .O(N__44574),
            .I(N__44547));
    InMux I__6544 (
            .O(N__44573),
            .I(N__44547));
    InMux I__6543 (
            .O(N__44572),
            .I(N__44544));
    InMux I__6542 (
            .O(N__44571),
            .I(N__44539));
    InMux I__6541 (
            .O(N__44570),
            .I(N__44539));
    LocalMux I__6540 (
            .O(N__44567),
            .I(N__44536));
    Odrv4 I__6539 (
            .O(N__44564),
            .I(\ppm_encoder_1.N_509 ));
    Odrv4 I__6538 (
            .O(N__44559),
            .I(\ppm_encoder_1.N_509 ));
    Odrv12 I__6537 (
            .O(N__44552),
            .I(\ppm_encoder_1.N_509 ));
    LocalMux I__6536 (
            .O(N__44547),
            .I(\ppm_encoder_1.N_509 ));
    LocalMux I__6535 (
            .O(N__44544),
            .I(\ppm_encoder_1.N_509 ));
    LocalMux I__6534 (
            .O(N__44539),
            .I(\ppm_encoder_1.N_509 ));
    Odrv4 I__6533 (
            .O(N__44536),
            .I(\ppm_encoder_1.N_509 ));
    CascadeMux I__6532 (
            .O(N__44521),
            .I(\ppm_encoder_1.un2_throttle_iv_i_i_0_14_cascade_ ));
    CascadeMux I__6531 (
            .O(N__44518),
            .I(N__44515));
    InMux I__6530 (
            .O(N__44515),
            .I(N__44506));
    InMux I__6529 (
            .O(N__44514),
            .I(N__44503));
    InMux I__6528 (
            .O(N__44513),
            .I(N__44499));
    InMux I__6527 (
            .O(N__44512),
            .I(N__44496));
    InMux I__6526 (
            .O(N__44511),
            .I(N__44493));
    InMux I__6525 (
            .O(N__44510),
            .I(N__44490));
    InMux I__6524 (
            .O(N__44509),
            .I(N__44487));
    LocalMux I__6523 (
            .O(N__44506),
            .I(N__44482));
    LocalMux I__6522 (
            .O(N__44503),
            .I(N__44482));
    InMux I__6521 (
            .O(N__44502),
            .I(N__44479));
    LocalMux I__6520 (
            .O(N__44499),
            .I(N__44475));
    LocalMux I__6519 (
            .O(N__44496),
            .I(N__44468));
    LocalMux I__6518 (
            .O(N__44493),
            .I(N__44468));
    LocalMux I__6517 (
            .O(N__44490),
            .I(N__44468));
    LocalMux I__6516 (
            .O(N__44487),
            .I(N__44459));
    Span4Mux_v I__6515 (
            .O(N__44482),
            .I(N__44459));
    LocalMux I__6514 (
            .O(N__44479),
            .I(N__44459));
    InMux I__6513 (
            .O(N__44478),
            .I(N__44453));
    Span4Mux_s2_v I__6512 (
            .O(N__44475),
            .I(N__44448));
    Span4Mux_v I__6511 (
            .O(N__44468),
            .I(N__44448));
    InMux I__6510 (
            .O(N__44467),
            .I(N__44445));
    InMux I__6509 (
            .O(N__44466),
            .I(N__44442));
    Span4Mux_h I__6508 (
            .O(N__44459),
            .I(N__44439));
    InMux I__6507 (
            .O(N__44458),
            .I(N__44434));
    InMux I__6506 (
            .O(N__44457),
            .I(N__44434));
    InMux I__6505 (
            .O(N__44456),
            .I(N__44431));
    LocalMux I__6504 (
            .O(N__44453),
            .I(N__44422));
    Span4Mux_h I__6503 (
            .O(N__44448),
            .I(N__44422));
    LocalMux I__6502 (
            .O(N__44445),
            .I(N__44422));
    LocalMux I__6501 (
            .O(N__44442),
            .I(N__44422));
    Odrv4 I__6500 (
            .O(N__44439),
            .I(\ppm_encoder_1.N_303 ));
    LocalMux I__6499 (
            .O(N__44434),
            .I(\ppm_encoder_1.N_303 ));
    LocalMux I__6498 (
            .O(N__44431),
            .I(\ppm_encoder_1.N_303 ));
    Odrv4 I__6497 (
            .O(N__44422),
            .I(\ppm_encoder_1.N_303 ));
    CascadeMux I__6496 (
            .O(N__44413),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_14_cascade_ ));
    InMux I__6495 (
            .O(N__44410),
            .I(N__44407));
    LocalMux I__6494 (
            .O(N__44407),
            .I(N__44404));
    Odrv4 I__6493 (
            .O(N__44404),
            .I(\ppm_encoder_1.init_pulses_RNIP98N6Z0Z_14 ));
    InMux I__6492 (
            .O(N__44401),
            .I(N__44398));
    LocalMux I__6491 (
            .O(N__44398),
            .I(N__44395));
    Span4Mux_h I__6490 (
            .O(N__44395),
            .I(N__44392));
    Odrv4 I__6489 (
            .O(N__44392),
            .I(\ppm_encoder_1.rudderZ0Z_14 ));
    CascadeMux I__6488 (
            .O(N__44389),
            .I(N__44386));
    InMux I__6487 (
            .O(N__44386),
            .I(N__44383));
    LocalMux I__6486 (
            .O(N__44383),
            .I(N__44379));
    InMux I__6485 (
            .O(N__44382),
            .I(N__44376));
    Odrv12 I__6484 (
            .O(N__44379),
            .I(\ppm_encoder_1.N_269_i_i ));
    LocalMux I__6483 (
            .O(N__44376),
            .I(\ppm_encoder_1.N_269_i_i ));
    InMux I__6482 (
            .O(N__44371),
            .I(N__44368));
    LocalMux I__6481 (
            .O(N__44368),
            .I(N__44365));
    Odrv4 I__6480 (
            .O(N__44365),
            .I(\ppm_encoder_1.pulses2count_9_0_0_11 ));
    CascadeMux I__6479 (
            .O(N__44362),
            .I(N__44359));
    InMux I__6478 (
            .O(N__44359),
            .I(N__44356));
    LocalMux I__6477 (
            .O(N__44356),
            .I(N__44353));
    Odrv4 I__6476 (
            .O(N__44353),
            .I(\ppm_encoder_1.N_431 ));
    InMux I__6475 (
            .O(N__44350),
            .I(N__44347));
    LocalMux I__6474 (
            .O(N__44347),
            .I(\ppm_encoder_1.N_269_i ));
    InMux I__6473 (
            .O(N__44344),
            .I(N__44340));
    InMux I__6472 (
            .O(N__44343),
            .I(N__44337));
    LocalMux I__6471 (
            .O(N__44340),
            .I(N__44334));
    LocalMux I__6470 (
            .O(N__44337),
            .I(N__44331));
    Span4Mux_h I__6469 (
            .O(N__44334),
            .I(N__44325));
    Span4Mux_s2_v I__6468 (
            .O(N__44331),
            .I(N__44322));
    InMux I__6467 (
            .O(N__44330),
            .I(N__44319));
    InMux I__6466 (
            .O(N__44329),
            .I(N__44314));
    InMux I__6465 (
            .O(N__44328),
            .I(N__44314));
    Odrv4 I__6464 (
            .O(N__44325),
            .I(\ppm_encoder_1.init_pulses_4_sqmuxa_i_0_0_0 ));
    Odrv4 I__6463 (
            .O(N__44322),
            .I(\ppm_encoder_1.init_pulses_4_sqmuxa_i_0_0_0 ));
    LocalMux I__6462 (
            .O(N__44319),
            .I(\ppm_encoder_1.init_pulses_4_sqmuxa_i_0_0_0 ));
    LocalMux I__6461 (
            .O(N__44314),
            .I(\ppm_encoder_1.init_pulses_4_sqmuxa_i_0_0_0 ));
    InMux I__6460 (
            .O(N__44305),
            .I(N__44301));
    InMux I__6459 (
            .O(N__44304),
            .I(N__44298));
    LocalMux I__6458 (
            .O(N__44301),
            .I(\ppm_encoder_1.un2_throttle_iv_0_1_0 ));
    LocalMux I__6457 (
            .O(N__44298),
            .I(\ppm_encoder_1.un2_throttle_iv_0_1_0 ));
    InMux I__6456 (
            .O(N__44293),
            .I(N__44289));
    InMux I__6455 (
            .O(N__44292),
            .I(N__44286));
    LocalMux I__6454 (
            .O(N__44289),
            .I(\ppm_encoder_1.un2_throttle_iv_0_0_0 ));
    LocalMux I__6453 (
            .O(N__44286),
            .I(\ppm_encoder_1.un2_throttle_iv_0_0_0 ));
    CascadeMux I__6452 (
            .O(N__44281),
            .I(N__44275));
    InMux I__6451 (
            .O(N__44280),
            .I(N__44272));
    CascadeMux I__6450 (
            .O(N__44279),
            .I(N__44269));
    InMux I__6449 (
            .O(N__44278),
            .I(N__44266));
    InMux I__6448 (
            .O(N__44275),
            .I(N__44263));
    LocalMux I__6447 (
            .O(N__44272),
            .I(N__44260));
    InMux I__6446 (
            .O(N__44269),
            .I(N__44257));
    LocalMux I__6445 (
            .O(N__44266),
            .I(N__44251));
    LocalMux I__6444 (
            .O(N__44263),
            .I(N__44251));
    Span4Mux_h I__6443 (
            .O(N__44260),
            .I(N__44246));
    LocalMux I__6442 (
            .O(N__44257),
            .I(N__44246));
    InMux I__6441 (
            .O(N__44256),
            .I(N__44243));
    Span4Mux_s1_v I__6440 (
            .O(N__44251),
            .I(N__44240));
    Odrv4 I__6439 (
            .O(N__44246),
            .I(\ppm_encoder_1.N_257_i_i ));
    LocalMux I__6438 (
            .O(N__44243),
            .I(\ppm_encoder_1.N_257_i_i ));
    Odrv4 I__6437 (
            .O(N__44240),
            .I(\ppm_encoder_1.N_257_i_i ));
    InMux I__6436 (
            .O(N__44233),
            .I(N__44230));
    LocalMux I__6435 (
            .O(N__44230),
            .I(N__44227));
    Odrv4 I__6434 (
            .O(N__44227),
            .I(\ppm_encoder_1.throttle_RNI0EA05Z0Z_0 ));
    CascadeMux I__6433 (
            .O(N__44224),
            .I(N__44221));
    InMux I__6432 (
            .O(N__44221),
            .I(N__44217));
    InMux I__6431 (
            .O(N__44220),
            .I(N__44214));
    LocalMux I__6430 (
            .O(N__44217),
            .I(\ppm_encoder_1.N_266_i_i ));
    LocalMux I__6429 (
            .O(N__44214),
            .I(\ppm_encoder_1.N_266_i_i ));
    InMux I__6428 (
            .O(N__44209),
            .I(N__44206));
    LocalMux I__6427 (
            .O(N__44206),
            .I(N__44203));
    Span4Mux_h I__6426 (
            .O(N__44203),
            .I(N__44200));
    Odrv4 I__6425 (
            .O(N__44200),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_11 ));
    InMux I__6424 (
            .O(N__44197),
            .I(N__44194));
    LocalMux I__6423 (
            .O(N__44194),
            .I(\ppm_encoder_1.init_pulses_RNIU1F76Z0Z_11 ));
    CascadeMux I__6422 (
            .O(N__44191),
            .I(\ppm_encoder_1.N_263_i_cascade_ ));
    CascadeMux I__6421 (
            .O(N__44188),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_7_cascade_ ));
    InMux I__6420 (
            .O(N__44185),
            .I(N__44182));
    LocalMux I__6419 (
            .O(N__44182),
            .I(N__44179));
    Odrv4 I__6418 (
            .O(N__44179),
            .I(\ppm_encoder_1.init_pulses_RNISD9M6Z0Z_7 ));
    InMux I__6417 (
            .O(N__44176),
            .I(N__44173));
    LocalMux I__6416 (
            .O(N__44173),
            .I(\ppm_encoder_1.un2_throttle_iv_0_0_0_7 ));
    CascadeMux I__6415 (
            .O(N__44170),
            .I(N__44167));
    InMux I__6414 (
            .O(N__44167),
            .I(N__44164));
    LocalMux I__6413 (
            .O(N__44164),
            .I(N__44160));
    InMux I__6412 (
            .O(N__44163),
            .I(N__44157));
    Span4Mux_v I__6411 (
            .O(N__44160),
            .I(N__44154));
    LocalMux I__6410 (
            .O(N__44157),
            .I(\ppm_encoder_1.rudderZ0Z_7 ));
    Odrv4 I__6409 (
            .O(N__44154),
            .I(\ppm_encoder_1.rudderZ0Z_7 ));
    CascadeMux I__6408 (
            .O(N__44149),
            .I(N__44146));
    InMux I__6407 (
            .O(N__44146),
            .I(N__44143));
    LocalMux I__6406 (
            .O(N__44143),
            .I(N__44139));
    InMux I__6405 (
            .O(N__44142),
            .I(N__44136));
    Odrv4 I__6404 (
            .O(N__44139),
            .I(\ppm_encoder_1.N_263_i_i ));
    LocalMux I__6403 (
            .O(N__44136),
            .I(\ppm_encoder_1.N_263_i_i ));
    InMux I__6402 (
            .O(N__44131),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_11 ));
    InMux I__6401 (
            .O(N__44128),
            .I(N__44125));
    LocalMux I__6400 (
            .O(N__44125),
            .I(\ppm_encoder_1.init_pulses_RNI8L3H5Z0Z_13 ));
    CascadeMux I__6399 (
            .O(N__44122),
            .I(N__44119));
    InMux I__6398 (
            .O(N__44119),
            .I(N__44115));
    InMux I__6397 (
            .O(N__44118),
            .I(N__44110));
    LocalMux I__6396 (
            .O(N__44115),
            .I(N__44107));
    InMux I__6395 (
            .O(N__44114),
            .I(N__44104));
    InMux I__6394 (
            .O(N__44113),
            .I(N__44101));
    LocalMux I__6393 (
            .O(N__44110),
            .I(\ppm_encoder_1.N_268_i_i ));
    Odrv12 I__6392 (
            .O(N__44107),
            .I(\ppm_encoder_1.N_268_i_i ));
    LocalMux I__6391 (
            .O(N__44104),
            .I(\ppm_encoder_1.N_268_i_i ));
    LocalMux I__6390 (
            .O(N__44101),
            .I(\ppm_encoder_1.N_268_i_i ));
    InMux I__6389 (
            .O(N__44092),
            .I(N__44089));
    LocalMux I__6388 (
            .O(N__44089),
            .I(\ppm_encoder_1.un1_init_pulses_10_13 ));
    InMux I__6387 (
            .O(N__44086),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_12 ));
    InMux I__6386 (
            .O(N__44083),
            .I(N__44080));
    LocalMux I__6385 (
            .O(N__44080),
            .I(\ppm_encoder_1.un1_init_pulses_10_14 ));
    InMux I__6384 (
            .O(N__44077),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_13 ));
    InMux I__6383 (
            .O(N__44074),
            .I(N__44071));
    LocalMux I__6382 (
            .O(N__44071),
            .I(\ppm_encoder_1.init_pulses_RNILFR51Z0Z_15 ));
    CascadeMux I__6381 (
            .O(N__44068),
            .I(N__44065));
    InMux I__6380 (
            .O(N__44065),
            .I(N__44062));
    LocalMux I__6379 (
            .O(N__44062),
            .I(\ppm_encoder_1.N_254_i_i ));
    InMux I__6378 (
            .O(N__44059),
            .I(N__44056));
    LocalMux I__6377 (
            .O(N__44056),
            .I(\ppm_encoder_1.un1_init_pulses_10_15 ));
    InMux I__6376 (
            .O(N__44053),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_14 ));
    InMux I__6375 (
            .O(N__44050),
            .I(N__44047));
    LocalMux I__6374 (
            .O(N__44047),
            .I(\ppm_encoder_1.un1_init_pulses_10_16 ));
    InMux I__6373 (
            .O(N__44044),
            .I(bfn_9_4_0_));
    InMux I__6372 (
            .O(N__44041),
            .I(N__44038));
    LocalMux I__6371 (
            .O(N__44038),
            .I(N__44035));
    Span4Mux_h I__6370 (
            .O(N__44035),
            .I(N__44032));
    Odrv4 I__6369 (
            .O(N__44032),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_17 ));
    InMux I__6368 (
            .O(N__44029),
            .I(N__44026));
    LocalMux I__6367 (
            .O(N__44026),
            .I(\ppm_encoder_1.un1_init_pulses_10_17 ));
    InMux I__6366 (
            .O(N__44023),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_16 ));
    InMux I__6365 (
            .O(N__44020),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_17 ));
    InMux I__6364 (
            .O(N__44017),
            .I(N__44014));
    LocalMux I__6363 (
            .O(N__44014),
            .I(\ppm_encoder_1.un1_init_pulses_10_18 ));
    InMux I__6362 (
            .O(N__44011),
            .I(N__44008));
    LocalMux I__6361 (
            .O(N__44008),
            .I(N__44005));
    Span4Mux_s2_v I__6360 (
            .O(N__44005),
            .I(N__44002));
    Span4Mux_h I__6359 (
            .O(N__44002),
            .I(N__43999));
    Odrv4 I__6358 (
            .O(N__43999),
            .I(\ppm_encoder_1.init_pulses_RNIFTCL6Z0Z_4 ));
    CascadeMux I__6357 (
            .O(N__43996),
            .I(N__43993));
    InMux I__6356 (
            .O(N__43993),
            .I(N__43990));
    LocalMux I__6355 (
            .O(N__43990),
            .I(N__43987));
    Span4Mux_h I__6354 (
            .O(N__43987),
            .I(N__43983));
    InMux I__6353 (
            .O(N__43986),
            .I(N__43980));
    Odrv4 I__6352 (
            .O(N__43983),
            .I(\ppm_encoder_1.N_260_i_i ));
    LocalMux I__6351 (
            .O(N__43980),
            .I(\ppm_encoder_1.N_260_i_i ));
    InMux I__6350 (
            .O(N__43975),
            .I(N__43972));
    LocalMux I__6349 (
            .O(N__43972),
            .I(N__43969));
    Odrv12 I__6348 (
            .O(N__43969),
            .I(\ppm_encoder_1.un1_init_pulses_10_4 ));
    InMux I__6347 (
            .O(N__43966),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_3 ));
    InMux I__6346 (
            .O(N__43963),
            .I(N__43960));
    LocalMux I__6345 (
            .O(N__43960),
            .I(N__43957));
    Odrv12 I__6344 (
            .O(N__43957),
            .I(\ppm_encoder_1.init_pulses_RNI3K6R5Z0Z_5 ));
    CascadeMux I__6343 (
            .O(N__43954),
            .I(N__43951));
    InMux I__6342 (
            .O(N__43951),
            .I(N__43948));
    LocalMux I__6341 (
            .O(N__43948),
            .I(N__43945));
    Span4Mux_h I__6340 (
            .O(N__43945),
            .I(N__43941));
    InMux I__6339 (
            .O(N__43944),
            .I(N__43938));
    Odrv4 I__6338 (
            .O(N__43941),
            .I(\ppm_encoder_1.N_261_i_i ));
    LocalMux I__6337 (
            .O(N__43938),
            .I(\ppm_encoder_1.N_261_i_i ));
    InMux I__6336 (
            .O(N__43933),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_4 ));
    InMux I__6335 (
            .O(N__43930),
            .I(N__43927));
    LocalMux I__6334 (
            .O(N__43927),
            .I(\ppm_encoder_1.init_pulses_RNI20JF6Z0Z_6 ));
    InMux I__6333 (
            .O(N__43924),
            .I(N__43920));
    CascadeMux I__6332 (
            .O(N__43923),
            .I(N__43917));
    LocalMux I__6331 (
            .O(N__43920),
            .I(N__43913));
    InMux I__6330 (
            .O(N__43917),
            .I(N__43910));
    InMux I__6329 (
            .O(N__43916),
            .I(N__43907));
    Odrv4 I__6328 (
            .O(N__43913),
            .I(\ppm_encoder_1.N_262_i_i ));
    LocalMux I__6327 (
            .O(N__43910),
            .I(\ppm_encoder_1.N_262_i_i ));
    LocalMux I__6326 (
            .O(N__43907),
            .I(\ppm_encoder_1.N_262_i_i ));
    InMux I__6325 (
            .O(N__43900),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_5 ));
    InMux I__6324 (
            .O(N__43897),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_6 ));
    InMux I__6323 (
            .O(N__43894),
            .I(N__43891));
    LocalMux I__6322 (
            .O(N__43891),
            .I(N__43888));
    Span12Mux_s5_v I__6321 (
            .O(N__43888),
            .I(N__43885));
    Odrv12 I__6320 (
            .O(N__43885),
            .I(\ppm_encoder_1.init_pulses_RNIL76H6Z0Z_8 ));
    CascadeMux I__6319 (
            .O(N__43882),
            .I(N__43879));
    InMux I__6318 (
            .O(N__43879),
            .I(N__43876));
    LocalMux I__6317 (
            .O(N__43876),
            .I(N__43873));
    Span4Mux_h I__6316 (
            .O(N__43873),
            .I(N__43870));
    Span4Mux_h I__6315 (
            .O(N__43870),
            .I(N__43867));
    Odrv4 I__6314 (
            .O(N__43867),
            .I(\ppm_encoder_1.N_264_i_i ));
    InMux I__6313 (
            .O(N__43864),
            .I(bfn_9_3_0_));
    InMux I__6312 (
            .O(N__43861),
            .I(N__43858));
    LocalMux I__6311 (
            .O(N__43858),
            .I(N__43855));
    Span4Mux_h I__6310 (
            .O(N__43855),
            .I(N__43852));
    Odrv4 I__6309 (
            .O(N__43852),
            .I(\ppm_encoder_1.init_pulses_RNIOCUG6Z0Z_9 ));
    CascadeMux I__6308 (
            .O(N__43849),
            .I(N__43846));
    InMux I__6307 (
            .O(N__43846),
            .I(N__43842));
    InMux I__6306 (
            .O(N__43845),
            .I(N__43839));
    LocalMux I__6305 (
            .O(N__43842),
            .I(N__43836));
    LocalMux I__6304 (
            .O(N__43839),
            .I(N__43833));
    Span4Mux_s2_v I__6303 (
            .O(N__43836),
            .I(N__43828));
    Span4Mux_v I__6302 (
            .O(N__43833),
            .I(N__43828));
    Odrv4 I__6301 (
            .O(N__43828),
            .I(\ppm_encoder_1.N_265_i_i ));
    InMux I__6300 (
            .O(N__43825),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_8 ));
    InMux I__6299 (
            .O(N__43822),
            .I(N__43819));
    LocalMux I__6298 (
            .O(N__43819),
            .I(N__43816));
    Span4Mux_h I__6297 (
            .O(N__43816),
            .I(N__43813));
    Odrv4 I__6296 (
            .O(N__43813),
            .I(\ppm_encoder_1.init_pulses_RNI8E326Z0Z_10 ));
    CascadeMux I__6295 (
            .O(N__43810),
            .I(N__43807));
    InMux I__6294 (
            .O(N__43807),
            .I(N__43804));
    LocalMux I__6293 (
            .O(N__43804),
            .I(N__43800));
    InMux I__6292 (
            .O(N__43803),
            .I(N__43797));
    Odrv4 I__6291 (
            .O(N__43800),
            .I(\ppm_encoder_1.N_255_i_i ));
    LocalMux I__6290 (
            .O(N__43797),
            .I(\ppm_encoder_1.N_255_i_i ));
    InMux I__6289 (
            .O(N__43792),
            .I(N__43789));
    LocalMux I__6288 (
            .O(N__43789),
            .I(\ppm_encoder_1.un1_init_pulses_10_10 ));
    InMux I__6287 (
            .O(N__43786),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_9 ));
    InMux I__6286 (
            .O(N__43783),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_10 ));
    InMux I__6285 (
            .O(N__43780),
            .I(N__43774));
    InMux I__6284 (
            .O(N__43779),
            .I(N__43774));
    LocalMux I__6283 (
            .O(N__43774),
            .I(\ppm_encoder_1.elevatorZ0Z_6 ));
    InMux I__6282 (
            .O(N__43771),
            .I(N__43768));
    LocalMux I__6281 (
            .O(N__43768),
            .I(N__43765));
    Span4Mux_h I__6280 (
            .O(N__43765),
            .I(N__43761));
    InMux I__6279 (
            .O(N__43764),
            .I(N__43758));
    Sp12to4 I__6278 (
            .O(N__43761),
            .I(N__43755));
    LocalMux I__6277 (
            .O(N__43758),
            .I(N__43752));
    Odrv12 I__6276 (
            .O(N__43755),
            .I(scaler_4_data_6));
    Odrv4 I__6275 (
            .O(N__43752),
            .I(scaler_4_data_6));
    InMux I__6274 (
            .O(N__43747),
            .I(N__43741));
    InMux I__6273 (
            .O(N__43746),
            .I(N__43741));
    LocalMux I__6272 (
            .O(N__43741),
            .I(\ppm_encoder_1.rudderZ0Z_6 ));
    InMux I__6271 (
            .O(N__43738),
            .I(N__43731));
    InMux I__6270 (
            .O(N__43737),
            .I(N__43731));
    CascadeMux I__6269 (
            .O(N__43736),
            .I(N__43728));
    LocalMux I__6268 (
            .O(N__43731),
            .I(N__43723));
    InMux I__6267 (
            .O(N__43728),
            .I(N__43718));
    InMux I__6266 (
            .O(N__43727),
            .I(N__43718));
    CascadeMux I__6265 (
            .O(N__43726),
            .I(N__43714));
    Span4Mux_s2_v I__6264 (
            .O(N__43723),
            .I(N__43708));
    LocalMux I__6263 (
            .O(N__43718),
            .I(N__43705));
    CascadeMux I__6262 (
            .O(N__43717),
            .I(N__43702));
    InMux I__6261 (
            .O(N__43714),
            .I(N__43698));
    InMux I__6260 (
            .O(N__43713),
            .I(N__43691));
    InMux I__6259 (
            .O(N__43712),
            .I(N__43691));
    InMux I__6258 (
            .O(N__43711),
            .I(N__43691));
    Span4Mux_h I__6257 (
            .O(N__43708),
            .I(N__43686));
    Span4Mux_s2_v I__6256 (
            .O(N__43705),
            .I(N__43686));
    InMux I__6255 (
            .O(N__43702),
            .I(N__43681));
    InMux I__6254 (
            .O(N__43701),
            .I(N__43681));
    LocalMux I__6253 (
            .O(N__43698),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z1 ));
    LocalMux I__6252 (
            .O(N__43691),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z1 ));
    Odrv4 I__6251 (
            .O(N__43686),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z1 ));
    LocalMux I__6250 (
            .O(N__43681),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z1 ));
    CascadeMux I__6249 (
            .O(N__43672),
            .I(\ppm_encoder_1.N_262_i_i_cascade_ ));
    InMux I__6248 (
            .O(N__43669),
            .I(N__43666));
    LocalMux I__6247 (
            .O(N__43666),
            .I(N__43663));
    Span4Mux_s2_v I__6246 (
            .O(N__43663),
            .I(N__43660));
    Span4Mux_h I__6245 (
            .O(N__43660),
            .I(N__43657));
    Odrv4 I__6244 (
            .O(N__43657),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_6 ));
    CascadeMux I__6243 (
            .O(N__43654),
            .I(N__43651));
    InMux I__6242 (
            .O(N__43651),
            .I(N__43648));
    LocalMux I__6241 (
            .O(N__43648),
            .I(\ppm_encoder_1.init_pulses_RNIQOIP3Z0Z_6 ));
    InMux I__6240 (
            .O(N__43645),
            .I(N__43642));
    LocalMux I__6239 (
            .O(N__43642),
            .I(N__43639));
    Span4Mux_h I__6238 (
            .O(N__43639),
            .I(N__43636));
    Odrv4 I__6237 (
            .O(N__43636),
            .I(\ppm_encoder_1.init_pulses_RNI29LM5Z0Z_1 ));
    CascadeMux I__6236 (
            .O(N__43633),
            .I(N__43630));
    InMux I__6235 (
            .O(N__43630),
            .I(N__43627));
    LocalMux I__6234 (
            .O(N__43627),
            .I(N__43623));
    InMux I__6233 (
            .O(N__43626),
            .I(N__43620));
    Span4Mux_h I__6232 (
            .O(N__43623),
            .I(N__43617));
    LocalMux I__6231 (
            .O(N__43620),
            .I(N__43614));
    Odrv4 I__6230 (
            .O(N__43617),
            .I(\ppm_encoder_1.N_258_i_i ));
    Odrv4 I__6229 (
            .O(N__43614),
            .I(\ppm_encoder_1.N_258_i_i ));
    InMux I__6228 (
            .O(N__43609),
            .I(N__43606));
    LocalMux I__6227 (
            .O(N__43606),
            .I(N__43603));
    Odrv12 I__6226 (
            .O(N__43603),
            .I(\ppm_encoder_1.un1_init_pulses_10_1 ));
    InMux I__6225 (
            .O(N__43600),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_0 ));
    InMux I__6224 (
            .O(N__43597),
            .I(N__43594));
    LocalMux I__6223 (
            .O(N__43594),
            .I(N__43591));
    Span12Mux_s4_v I__6222 (
            .O(N__43591),
            .I(N__43588));
    Odrv12 I__6221 (
            .O(N__43588),
            .I(\ppm_encoder_1.init_pulses_RNIIIS46Z0Z_2 ));
    CascadeMux I__6220 (
            .O(N__43585),
            .I(N__43581));
    InMux I__6219 (
            .O(N__43584),
            .I(N__43578));
    InMux I__6218 (
            .O(N__43581),
            .I(N__43575));
    LocalMux I__6217 (
            .O(N__43578),
            .I(N__43570));
    LocalMux I__6216 (
            .O(N__43575),
            .I(N__43570));
    Span4Mux_s3_v I__6215 (
            .O(N__43570),
            .I(N__43566));
    InMux I__6214 (
            .O(N__43569),
            .I(N__43563));
    Span4Mux_h I__6213 (
            .O(N__43566),
            .I(N__43559));
    LocalMux I__6212 (
            .O(N__43563),
            .I(N__43556));
    InMux I__6211 (
            .O(N__43562),
            .I(N__43553));
    Odrv4 I__6210 (
            .O(N__43559),
            .I(\ppm_encoder_1.N_259_i_i ));
    Odrv4 I__6209 (
            .O(N__43556),
            .I(\ppm_encoder_1.N_259_i_i ));
    LocalMux I__6208 (
            .O(N__43553),
            .I(\ppm_encoder_1.N_259_i_i ));
    InMux I__6207 (
            .O(N__43546),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_1 ));
    InMux I__6206 (
            .O(N__43543),
            .I(N__43540));
    LocalMux I__6205 (
            .O(N__43540),
            .I(N__43537));
    Span4Mux_h I__6204 (
            .O(N__43537),
            .I(N__43534));
    Odrv4 I__6203 (
            .O(N__43534),
            .I(\ppm_encoder_1.init_pulses_RNINNS46Z0Z_3 ));
    CascadeMux I__6202 (
            .O(N__43531),
            .I(N__43528));
    InMux I__6201 (
            .O(N__43528),
            .I(N__43525));
    LocalMux I__6200 (
            .O(N__43525),
            .I(N__43521));
    InMux I__6199 (
            .O(N__43524),
            .I(N__43518));
    Span4Mux_s1_v I__6198 (
            .O(N__43521),
            .I(N__43515));
    LocalMux I__6197 (
            .O(N__43518),
            .I(N__43512));
    Odrv4 I__6196 (
            .O(N__43515),
            .I(\ppm_encoder_1.N_256_i_i ));
    Odrv12 I__6195 (
            .O(N__43512),
            .I(\ppm_encoder_1.N_256_i_i ));
    InMux I__6194 (
            .O(N__43507),
            .I(N__43504));
    LocalMux I__6193 (
            .O(N__43504),
            .I(N__43501));
    Odrv12 I__6192 (
            .O(N__43501),
            .I(\ppm_encoder_1.un1_init_pulses_10_3 ));
    InMux I__6191 (
            .O(N__43498),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_2 ));
    InMux I__6190 (
            .O(N__43495),
            .I(N__43490));
    InMux I__6189 (
            .O(N__43494),
            .I(N__43485));
    InMux I__6188 (
            .O(N__43493),
            .I(N__43485));
    LocalMux I__6187 (
            .O(N__43490),
            .I(\dron_frame_decoder_1.WDTZ0Z_12 ));
    LocalMux I__6186 (
            .O(N__43485),
            .I(\dron_frame_decoder_1.WDTZ0Z_12 ));
    CascadeMux I__6185 (
            .O(N__43480),
            .I(N__43476));
    InMux I__6184 (
            .O(N__43479),
            .I(N__43471));
    InMux I__6183 (
            .O(N__43476),
            .I(N__43468));
    InMux I__6182 (
            .O(N__43475),
            .I(N__43463));
    InMux I__6181 (
            .O(N__43474),
            .I(N__43463));
    LocalMux I__6180 (
            .O(N__43471),
            .I(\dron_frame_decoder_1.WDTZ0Z_13 ));
    LocalMux I__6179 (
            .O(N__43468),
            .I(\dron_frame_decoder_1.WDTZ0Z_13 ));
    LocalMux I__6178 (
            .O(N__43463),
            .I(\dron_frame_decoder_1.WDTZ0Z_13 ));
    InMux I__6177 (
            .O(N__43456),
            .I(N__43453));
    LocalMux I__6176 (
            .O(N__43453),
            .I(\dron_frame_decoder_1.WDT10lt12_0 ));
    CascadeMux I__6175 (
            .O(N__43450),
            .I(N__43445));
    InMux I__6174 (
            .O(N__43449),
            .I(N__43442));
    InMux I__6173 (
            .O(N__43448),
            .I(N__43437));
    InMux I__6172 (
            .O(N__43445),
            .I(N__43437));
    LocalMux I__6171 (
            .O(N__43442),
            .I(\dron_frame_decoder_1.WDTZ0Z_14 ));
    LocalMux I__6170 (
            .O(N__43437),
            .I(\dron_frame_decoder_1.WDTZ0Z_14 ));
    CascadeMux I__6169 (
            .O(N__43432),
            .I(\dron_frame_decoder_1.WDT10lt14_0_cascade_ ));
    InMux I__6168 (
            .O(N__43429),
            .I(N__43424));
    InMux I__6167 (
            .O(N__43428),
            .I(N__43419));
    InMux I__6166 (
            .O(N__43427),
            .I(N__43419));
    LocalMux I__6165 (
            .O(N__43424),
            .I(\dron_frame_decoder_1.WDTZ0Z_15 ));
    LocalMux I__6164 (
            .O(N__43419),
            .I(\dron_frame_decoder_1.WDTZ0Z_15 ));
    CascadeMux I__6163 (
            .O(N__43414),
            .I(\dron_frame_decoder_1.N_218_cascade_ ));
    InMux I__6162 (
            .O(N__43411),
            .I(N__43406));
    InMux I__6161 (
            .O(N__43410),
            .I(N__43403));
    InMux I__6160 (
            .O(N__43409),
            .I(N__43400));
    LocalMux I__6159 (
            .O(N__43406),
            .I(\dron_frame_decoder_1.stateZ0Z_2 ));
    LocalMux I__6158 (
            .O(N__43403),
            .I(\dron_frame_decoder_1.stateZ0Z_2 ));
    LocalMux I__6157 (
            .O(N__43400),
            .I(\dron_frame_decoder_1.stateZ0Z_2 ));
    CascadeMux I__6156 (
            .O(N__43393),
            .I(\ppm_encoder_1.N_262_i_cascade_ ));
    CascadeMux I__6155 (
            .O(N__43390),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_6_cascade_ ));
    InMux I__6154 (
            .O(N__43387),
            .I(\dron_frame_decoder_1.un1_WDT_cry_11 ));
    InMux I__6153 (
            .O(N__43384),
            .I(\dron_frame_decoder_1.un1_WDT_cry_12 ));
    InMux I__6152 (
            .O(N__43381),
            .I(\dron_frame_decoder_1.un1_WDT_cry_13 ));
    InMux I__6151 (
            .O(N__43378),
            .I(\dron_frame_decoder_1.un1_WDT_cry_14 ));
    SRMux I__6150 (
            .O(N__43375),
            .I(N__43372));
    LocalMux I__6149 (
            .O(N__43372),
            .I(N__43368));
    SRMux I__6148 (
            .O(N__43371),
            .I(N__43365));
    Span4Mux_h I__6147 (
            .O(N__43368),
            .I(N__43362));
    LocalMux I__6146 (
            .O(N__43365),
            .I(N__43359));
    Span4Mux_h I__6145 (
            .O(N__43362),
            .I(N__43356));
    Span4Mux_h I__6144 (
            .O(N__43359),
            .I(N__43353));
    Odrv4 I__6143 (
            .O(N__43356),
            .I(\dron_frame_decoder_1.source_data_valid_2_sqmuxa_iZ0 ));
    Odrv4 I__6142 (
            .O(N__43353),
            .I(\dron_frame_decoder_1.source_data_valid_2_sqmuxa_iZ0 ));
    InMux I__6141 (
            .O(N__43348),
            .I(N__43344));
    InMux I__6140 (
            .O(N__43347),
            .I(N__43341));
    LocalMux I__6139 (
            .O(N__43344),
            .I(N__43338));
    LocalMux I__6138 (
            .O(N__43341),
            .I(\dron_frame_decoder_1.WDTZ0Z_6 ));
    Odrv4 I__6137 (
            .O(N__43338),
            .I(\dron_frame_decoder_1.WDTZ0Z_6 ));
    InMux I__6136 (
            .O(N__43333),
            .I(N__43329));
    InMux I__6135 (
            .O(N__43332),
            .I(N__43326));
    LocalMux I__6134 (
            .O(N__43329),
            .I(N__43323));
    LocalMux I__6133 (
            .O(N__43326),
            .I(\dron_frame_decoder_1.WDTZ0Z_7 ));
    Odrv4 I__6132 (
            .O(N__43323),
            .I(\dron_frame_decoder_1.WDTZ0Z_7 ));
    CascadeMux I__6131 (
            .O(N__43318),
            .I(N__43314));
    InMux I__6130 (
            .O(N__43317),
            .I(N__43311));
    InMux I__6129 (
            .O(N__43314),
            .I(N__43308));
    LocalMux I__6128 (
            .O(N__43311),
            .I(\dron_frame_decoder_1.WDTZ0Z_10 ));
    LocalMux I__6127 (
            .O(N__43308),
            .I(\dron_frame_decoder_1.WDTZ0Z_10 ));
    CascadeMux I__6126 (
            .O(N__43303),
            .I(\dron_frame_decoder_1.WDT10lt12_0_cascade_ ));
    CascadeMux I__6125 (
            .O(N__43300),
            .I(N__43296));
    InMux I__6124 (
            .O(N__43299),
            .I(N__43293));
    InMux I__6123 (
            .O(N__43296),
            .I(N__43290));
    LocalMux I__6122 (
            .O(N__43293),
            .I(N__43285));
    LocalMux I__6121 (
            .O(N__43290),
            .I(N__43285));
    Odrv4 I__6120 (
            .O(N__43285),
            .I(\dron_frame_decoder_1.WDT10_0_i ));
    InMux I__6119 (
            .O(N__43282),
            .I(N__43279));
    LocalMux I__6118 (
            .O(N__43279),
            .I(\dron_frame_decoder_1.WDT10_0_i_1 ));
    InMux I__6117 (
            .O(N__43276),
            .I(N__43272));
    InMux I__6116 (
            .O(N__43275),
            .I(N__43269));
    LocalMux I__6115 (
            .O(N__43272),
            .I(\dron_frame_decoder_1.WDTZ0Z_8 ));
    LocalMux I__6114 (
            .O(N__43269),
            .I(\dron_frame_decoder_1.WDTZ0Z_8 ));
    InMux I__6113 (
            .O(N__43264),
            .I(N__43260));
    InMux I__6112 (
            .O(N__43263),
            .I(N__43257));
    LocalMux I__6111 (
            .O(N__43260),
            .I(N__43254));
    LocalMux I__6110 (
            .O(N__43257),
            .I(\dron_frame_decoder_1.WDTZ0Z_5 ));
    Odrv4 I__6109 (
            .O(N__43254),
            .I(\dron_frame_decoder_1.WDTZ0Z_5 ));
    CascadeMux I__6108 (
            .O(N__43249),
            .I(N__43245));
    InMux I__6107 (
            .O(N__43248),
            .I(N__43242));
    InMux I__6106 (
            .O(N__43245),
            .I(N__43239));
    LocalMux I__6105 (
            .O(N__43242),
            .I(\dron_frame_decoder_1.WDTZ0Z_9 ));
    LocalMux I__6104 (
            .O(N__43239),
            .I(\dron_frame_decoder_1.WDTZ0Z_9 ));
    InMux I__6103 (
            .O(N__43234),
            .I(N__43230));
    InMux I__6102 (
            .O(N__43233),
            .I(N__43227));
    LocalMux I__6101 (
            .O(N__43230),
            .I(N__43224));
    LocalMux I__6100 (
            .O(N__43227),
            .I(\dron_frame_decoder_1.WDTZ0Z_4 ));
    Odrv4 I__6099 (
            .O(N__43224),
            .I(\dron_frame_decoder_1.WDTZ0Z_4 ));
    InMux I__6098 (
            .O(N__43219),
            .I(N__43216));
    LocalMux I__6097 (
            .O(N__43216),
            .I(\dron_frame_decoder_1.WDT10lto9_3 ));
    InMux I__6096 (
            .O(N__43213),
            .I(N__43208));
    InMux I__6095 (
            .O(N__43212),
            .I(N__43203));
    InMux I__6094 (
            .O(N__43211),
            .I(N__43203));
    LocalMux I__6093 (
            .O(N__43208),
            .I(\dron_frame_decoder_1.WDTZ0Z_11 ));
    LocalMux I__6092 (
            .O(N__43203),
            .I(\dron_frame_decoder_1.WDTZ0Z_11 ));
    InMux I__6091 (
            .O(N__43198),
            .I(N__43195));
    LocalMux I__6090 (
            .O(N__43195),
            .I(\dron_frame_decoder_1.WDTZ0Z_3 ));
    InMux I__6089 (
            .O(N__43192),
            .I(\dron_frame_decoder_1.un1_WDT_cry_2 ));
    InMux I__6088 (
            .O(N__43189),
            .I(\dron_frame_decoder_1.un1_WDT_cry_3 ));
    InMux I__6087 (
            .O(N__43186),
            .I(\dron_frame_decoder_1.un1_WDT_cry_4 ));
    InMux I__6086 (
            .O(N__43183),
            .I(\dron_frame_decoder_1.un1_WDT_cry_5 ));
    InMux I__6085 (
            .O(N__43180),
            .I(\dron_frame_decoder_1.un1_WDT_cry_6 ));
    InMux I__6084 (
            .O(N__43177),
            .I(bfn_8_19_0_));
    InMux I__6083 (
            .O(N__43174),
            .I(\dron_frame_decoder_1.un1_WDT_cry_8 ));
    InMux I__6082 (
            .O(N__43171),
            .I(\dron_frame_decoder_1.un1_WDT_cry_9 ));
    InMux I__6081 (
            .O(N__43168),
            .I(\dron_frame_decoder_1.un1_WDT_cry_10 ));
    CascadeMux I__6080 (
            .O(N__43165),
            .I(\uart_pc.timer_Count_RNILR1B2Z0Z_2_cascade_ ));
    CascadeMux I__6079 (
            .O(N__43162),
            .I(\Commands_frame_decoder.state_ns_i_a2_2_1Z0Z_0_cascade_ ));
    InMux I__6078 (
            .O(N__43159),
            .I(N__43154));
    InMux I__6077 (
            .O(N__43158),
            .I(N__43149));
    InMux I__6076 (
            .O(N__43157),
            .I(N__43149));
    LocalMux I__6075 (
            .O(N__43154),
            .I(N__43146));
    LocalMux I__6074 (
            .O(N__43149),
            .I(\Commands_frame_decoder.N_410 ));
    Odrv4 I__6073 (
            .O(N__43146),
            .I(\Commands_frame_decoder.N_410 ));
    CascadeMux I__6072 (
            .O(N__43141),
            .I(\uart_pc.timer_Count_RNIMQ8T1Z0Z_2_cascade_ ));
    InMux I__6071 (
            .O(N__43138),
            .I(N__43135));
    LocalMux I__6070 (
            .O(N__43135),
            .I(\dron_frame_decoder_1.WDTZ0Z_0 ));
    InMux I__6069 (
            .O(N__43132),
            .I(N__43129));
    LocalMux I__6068 (
            .O(N__43129),
            .I(\dron_frame_decoder_1.WDTZ0Z_1 ));
    InMux I__6067 (
            .O(N__43126),
            .I(\dron_frame_decoder_1.un1_WDT_cry_0 ));
    InMux I__6066 (
            .O(N__43123),
            .I(N__43120));
    LocalMux I__6065 (
            .O(N__43120),
            .I(\dron_frame_decoder_1.WDTZ0Z_2 ));
    InMux I__6064 (
            .O(N__43117),
            .I(\dron_frame_decoder_1.un1_WDT_cry_1 ));
    CascadeMux I__6063 (
            .O(N__43114),
            .I(\uart_pc.CO0_cascade_ ));
    InMux I__6062 (
            .O(N__43111),
            .I(N__43105));
    InMux I__6061 (
            .O(N__43110),
            .I(N__43105));
    LocalMux I__6060 (
            .O(N__43105),
            .I(\uart_pc.un1_state_7_0 ));
    InMux I__6059 (
            .O(N__43102),
            .I(N__43092));
    InMux I__6058 (
            .O(N__43101),
            .I(N__43092));
    InMux I__6057 (
            .O(N__43100),
            .I(N__43092));
    InMux I__6056 (
            .O(N__43099),
            .I(N__43089));
    LocalMux I__6055 (
            .O(N__43092),
            .I(\uart_pc.un1_state_4_0 ));
    LocalMux I__6054 (
            .O(N__43089),
            .I(\uart_pc.un1_state_4_0 ));
    InMux I__6053 (
            .O(N__43084),
            .I(N__43063));
    InMux I__6052 (
            .O(N__43083),
            .I(N__43063));
    InMux I__6051 (
            .O(N__43082),
            .I(N__43063));
    InMux I__6050 (
            .O(N__43081),
            .I(N__43063));
    InMux I__6049 (
            .O(N__43080),
            .I(N__43063));
    InMux I__6048 (
            .O(N__43079),
            .I(N__43050));
    InMux I__6047 (
            .O(N__43078),
            .I(N__43050));
    InMux I__6046 (
            .O(N__43077),
            .I(N__43050));
    InMux I__6045 (
            .O(N__43076),
            .I(N__43050));
    InMux I__6044 (
            .O(N__43075),
            .I(N__43050));
    InMux I__6043 (
            .O(N__43074),
            .I(N__43050));
    LocalMux I__6042 (
            .O(N__43063),
            .I(\uart_pc.bit_CountZ0Z_0 ));
    LocalMux I__6041 (
            .O(N__43050),
            .I(\uart_pc.bit_CountZ0Z_0 ));
    CascadeMux I__6040 (
            .O(N__43045),
            .I(N__43038));
    CascadeMux I__6039 (
            .O(N__43044),
            .I(N__43035));
    CascadeMux I__6038 (
            .O(N__43043),
            .I(N__43030));
    CascadeMux I__6037 (
            .O(N__43042),
            .I(N__43026));
    InMux I__6036 (
            .O(N__43041),
            .I(N__43015));
    InMux I__6035 (
            .O(N__43038),
            .I(N__43015));
    InMux I__6034 (
            .O(N__43035),
            .I(N__43015));
    InMux I__6033 (
            .O(N__43034),
            .I(N__43015));
    InMux I__6032 (
            .O(N__43033),
            .I(N__43002));
    InMux I__6031 (
            .O(N__43030),
            .I(N__43002));
    InMux I__6030 (
            .O(N__43029),
            .I(N__43002));
    InMux I__6029 (
            .O(N__43026),
            .I(N__43002));
    InMux I__6028 (
            .O(N__43025),
            .I(N__43002));
    InMux I__6027 (
            .O(N__43024),
            .I(N__43002));
    LocalMux I__6026 (
            .O(N__43015),
            .I(\uart_pc.bit_CountZ0Z_1 ));
    LocalMux I__6025 (
            .O(N__43002),
            .I(\uart_pc.bit_CountZ0Z_1 ));
    InMux I__6024 (
            .O(N__42997),
            .I(N__42986));
    InMux I__6023 (
            .O(N__42996),
            .I(N__42981));
    InMux I__6022 (
            .O(N__42995),
            .I(N__42981));
    InMux I__6021 (
            .O(N__42994),
            .I(N__42968));
    InMux I__6020 (
            .O(N__42993),
            .I(N__42968));
    InMux I__6019 (
            .O(N__42992),
            .I(N__42968));
    InMux I__6018 (
            .O(N__42991),
            .I(N__42968));
    InMux I__6017 (
            .O(N__42990),
            .I(N__42968));
    InMux I__6016 (
            .O(N__42989),
            .I(N__42968));
    LocalMux I__6015 (
            .O(N__42986),
            .I(\uart_pc.bit_CountZ0Z_2 ));
    LocalMux I__6014 (
            .O(N__42981),
            .I(\uart_pc.bit_CountZ0Z_2 ));
    LocalMux I__6013 (
            .O(N__42968),
            .I(\uart_pc.bit_CountZ0Z_2 ));
    InMux I__6012 (
            .O(N__42961),
            .I(\Commands_frame_decoder.un1_WDT_cry_13 ));
    InMux I__6011 (
            .O(N__42958),
            .I(\Commands_frame_decoder.un1_WDT_cry_14 ));
    InMux I__6010 (
            .O(N__42955),
            .I(N__42952));
    LocalMux I__6009 (
            .O(N__42952),
            .I(N__42949));
    Span4Mux_h I__6008 (
            .O(N__42949),
            .I(N__42946));
    Span4Mux_v I__6007 (
            .O(N__42946),
            .I(N__42943));
    Span4Mux_h I__6006 (
            .O(N__42943),
            .I(N__42940));
    Odrv4 I__6005 (
            .O(N__42940),
            .I(scaler_4_data_5));
    CascadeMux I__6004 (
            .O(N__42937),
            .I(\uart_pc.N_152_cascade_ ));
    InMux I__6003 (
            .O(N__42934),
            .I(\Commands_frame_decoder.un1_WDT_cry_4 ));
    InMux I__6002 (
            .O(N__42931),
            .I(N__42926));
    InMux I__6001 (
            .O(N__42930),
            .I(N__42923));
    InMux I__6000 (
            .O(N__42929),
            .I(N__42920));
    LocalMux I__5999 (
            .O(N__42926),
            .I(\Commands_frame_decoder.WDTZ0Z_6 ));
    LocalMux I__5998 (
            .O(N__42923),
            .I(\Commands_frame_decoder.WDTZ0Z_6 ));
    LocalMux I__5997 (
            .O(N__42920),
            .I(\Commands_frame_decoder.WDTZ0Z_6 ));
    InMux I__5996 (
            .O(N__42913),
            .I(\Commands_frame_decoder.un1_WDT_cry_5 ));
    CascadeMux I__5995 (
            .O(N__42910),
            .I(N__42905));
    CascadeMux I__5994 (
            .O(N__42909),
            .I(N__42902));
    InMux I__5993 (
            .O(N__42908),
            .I(N__42899));
    InMux I__5992 (
            .O(N__42905),
            .I(N__42896));
    InMux I__5991 (
            .O(N__42902),
            .I(N__42893));
    LocalMux I__5990 (
            .O(N__42899),
            .I(\Commands_frame_decoder.WDTZ0Z_7 ));
    LocalMux I__5989 (
            .O(N__42896),
            .I(\Commands_frame_decoder.WDTZ0Z_7 ));
    LocalMux I__5988 (
            .O(N__42893),
            .I(\Commands_frame_decoder.WDTZ0Z_7 ));
    InMux I__5987 (
            .O(N__42886),
            .I(\Commands_frame_decoder.un1_WDT_cry_6 ));
    InMux I__5986 (
            .O(N__42883),
            .I(N__42878));
    InMux I__5985 (
            .O(N__42882),
            .I(N__42873));
    InMux I__5984 (
            .O(N__42881),
            .I(N__42873));
    LocalMux I__5983 (
            .O(N__42878),
            .I(\Commands_frame_decoder.WDTZ0Z_8 ));
    LocalMux I__5982 (
            .O(N__42873),
            .I(\Commands_frame_decoder.WDTZ0Z_8 ));
    InMux I__5981 (
            .O(N__42868),
            .I(bfn_8_14_0_));
    CascadeMux I__5980 (
            .O(N__42865),
            .I(N__42861));
    InMux I__5979 (
            .O(N__42864),
            .I(N__42857));
    InMux I__5978 (
            .O(N__42861),
            .I(N__42852));
    InMux I__5977 (
            .O(N__42860),
            .I(N__42852));
    LocalMux I__5976 (
            .O(N__42857),
            .I(\Commands_frame_decoder.WDTZ0Z_9 ));
    LocalMux I__5975 (
            .O(N__42852),
            .I(\Commands_frame_decoder.WDTZ0Z_9 ));
    InMux I__5974 (
            .O(N__42847),
            .I(\Commands_frame_decoder.un1_WDT_cry_8 ));
    InMux I__5973 (
            .O(N__42844),
            .I(N__42839));
    InMux I__5972 (
            .O(N__42843),
            .I(N__42836));
    InMux I__5971 (
            .O(N__42842),
            .I(N__42833));
    LocalMux I__5970 (
            .O(N__42839),
            .I(\Commands_frame_decoder.WDTZ0Z_10 ));
    LocalMux I__5969 (
            .O(N__42836),
            .I(\Commands_frame_decoder.WDTZ0Z_10 ));
    LocalMux I__5968 (
            .O(N__42833),
            .I(\Commands_frame_decoder.WDTZ0Z_10 ));
    InMux I__5967 (
            .O(N__42826),
            .I(\Commands_frame_decoder.un1_WDT_cry_9 ));
    InMux I__5966 (
            .O(N__42823),
            .I(N__42817));
    InMux I__5965 (
            .O(N__42822),
            .I(N__42812));
    InMux I__5964 (
            .O(N__42821),
            .I(N__42812));
    InMux I__5963 (
            .O(N__42820),
            .I(N__42809));
    LocalMux I__5962 (
            .O(N__42817),
            .I(\Commands_frame_decoder.WDTZ0Z_11 ));
    LocalMux I__5961 (
            .O(N__42812),
            .I(\Commands_frame_decoder.WDTZ0Z_11 ));
    LocalMux I__5960 (
            .O(N__42809),
            .I(\Commands_frame_decoder.WDTZ0Z_11 ));
    InMux I__5959 (
            .O(N__42802),
            .I(\Commands_frame_decoder.un1_WDT_cry_10 ));
    CascadeMux I__5958 (
            .O(N__42799),
            .I(N__42795));
    InMux I__5957 (
            .O(N__42798),
            .I(N__42790));
    InMux I__5956 (
            .O(N__42795),
            .I(N__42785));
    InMux I__5955 (
            .O(N__42794),
            .I(N__42785));
    InMux I__5954 (
            .O(N__42793),
            .I(N__42782));
    LocalMux I__5953 (
            .O(N__42790),
            .I(\Commands_frame_decoder.WDTZ0Z_12 ));
    LocalMux I__5952 (
            .O(N__42785),
            .I(\Commands_frame_decoder.WDTZ0Z_12 ));
    LocalMux I__5951 (
            .O(N__42782),
            .I(\Commands_frame_decoder.WDTZ0Z_12 ));
    InMux I__5950 (
            .O(N__42775),
            .I(\Commands_frame_decoder.un1_WDT_cry_11 ));
    InMux I__5949 (
            .O(N__42772),
            .I(N__42767));
    InMux I__5948 (
            .O(N__42771),
            .I(N__42764));
    InMux I__5947 (
            .O(N__42770),
            .I(N__42761));
    LocalMux I__5946 (
            .O(N__42767),
            .I(\Commands_frame_decoder.WDTZ0Z_13 ));
    LocalMux I__5945 (
            .O(N__42764),
            .I(\Commands_frame_decoder.WDTZ0Z_13 ));
    LocalMux I__5944 (
            .O(N__42761),
            .I(\Commands_frame_decoder.WDTZ0Z_13 ));
    InMux I__5943 (
            .O(N__42754),
            .I(\Commands_frame_decoder.un1_WDT_cry_12 ));
    InMux I__5942 (
            .O(N__42751),
            .I(\scaler_4.un3_source_data_0_cry_8 ));
    CascadeMux I__5941 (
            .O(N__42748),
            .I(N__42745));
    InMux I__5940 (
            .O(N__42745),
            .I(N__42742));
    LocalMux I__5939 (
            .O(N__42742),
            .I(\scaler_4.un3_source_data_0_cry_8_c_RNIS918 ));
    CEMux I__5938 (
            .O(N__42739),
            .I(N__42736));
    LocalMux I__5937 (
            .O(N__42736),
            .I(N__42732));
    CEMux I__5936 (
            .O(N__42735),
            .I(N__42729));
    Span4Mux_v I__5935 (
            .O(N__42732),
            .I(N__42726));
    LocalMux I__5934 (
            .O(N__42729),
            .I(N__42723));
    Sp12to4 I__5933 (
            .O(N__42726),
            .I(N__42718));
    Span12Mux_s11_v I__5932 (
            .O(N__42723),
            .I(N__42718));
    Odrv12 I__5931 (
            .O(N__42718),
            .I(\Commands_frame_decoder.state_RNIQRI31Z0Z_10 ));
    InMux I__5930 (
            .O(N__42715),
            .I(N__42712));
    LocalMux I__5929 (
            .O(N__42712),
            .I(\scaler_4.un3_source_data_0_axb_7 ));
    InMux I__5928 (
            .O(N__42709),
            .I(N__42705));
    CascadeMux I__5927 (
            .O(N__42708),
            .I(N__42702));
    LocalMux I__5926 (
            .O(N__42705),
            .I(N__42699));
    InMux I__5925 (
            .O(N__42702),
            .I(N__42696));
    Odrv4 I__5924 (
            .O(N__42699),
            .I(\Commands_frame_decoder.state_0_sqmuxa ));
    LocalMux I__5923 (
            .O(N__42696),
            .I(\Commands_frame_decoder.state_0_sqmuxa ));
    InMux I__5922 (
            .O(N__42691),
            .I(N__42688));
    LocalMux I__5921 (
            .O(N__42688),
            .I(\Commands_frame_decoder.WDTZ0Z_0 ));
    InMux I__5920 (
            .O(N__42685),
            .I(N__42682));
    LocalMux I__5919 (
            .O(N__42682),
            .I(\Commands_frame_decoder.WDTZ0Z_1 ));
    InMux I__5918 (
            .O(N__42679),
            .I(\Commands_frame_decoder.un1_WDT_cry_0 ));
    InMux I__5917 (
            .O(N__42676),
            .I(N__42673));
    LocalMux I__5916 (
            .O(N__42673),
            .I(\Commands_frame_decoder.WDTZ0Z_2 ));
    InMux I__5915 (
            .O(N__42670),
            .I(\Commands_frame_decoder.un1_WDT_cry_1 ));
    InMux I__5914 (
            .O(N__42667),
            .I(N__42664));
    LocalMux I__5913 (
            .O(N__42664),
            .I(\Commands_frame_decoder.WDTZ0Z_3 ));
    InMux I__5912 (
            .O(N__42661),
            .I(\Commands_frame_decoder.un1_WDT_cry_2 ));
    InMux I__5911 (
            .O(N__42658),
            .I(N__42653));
    InMux I__5910 (
            .O(N__42657),
            .I(N__42650));
    InMux I__5909 (
            .O(N__42656),
            .I(N__42647));
    LocalMux I__5908 (
            .O(N__42653),
            .I(\Commands_frame_decoder.WDTZ0Z_4 ));
    LocalMux I__5907 (
            .O(N__42650),
            .I(\Commands_frame_decoder.WDTZ0Z_4 ));
    LocalMux I__5906 (
            .O(N__42647),
            .I(\Commands_frame_decoder.WDTZ0Z_4 ));
    InMux I__5905 (
            .O(N__42640),
            .I(\Commands_frame_decoder.un1_WDT_cry_3 ));
    InMux I__5904 (
            .O(N__42637),
            .I(N__42632));
    InMux I__5903 (
            .O(N__42636),
            .I(N__42629));
    InMux I__5902 (
            .O(N__42635),
            .I(N__42626));
    LocalMux I__5901 (
            .O(N__42632),
            .I(\Commands_frame_decoder.WDTZ0Z_5 ));
    LocalMux I__5900 (
            .O(N__42629),
            .I(\Commands_frame_decoder.WDTZ0Z_5 ));
    LocalMux I__5899 (
            .O(N__42626),
            .I(\Commands_frame_decoder.WDTZ0Z_5 ));
    InMux I__5898 (
            .O(N__42619),
            .I(N__42616));
    LocalMux I__5897 (
            .O(N__42616),
            .I(frame_decoder_CH4data_1));
    InMux I__5896 (
            .O(N__42613),
            .I(\scaler_4.un3_source_data_0_cry_0 ));
    InMux I__5895 (
            .O(N__42610),
            .I(N__42607));
    LocalMux I__5894 (
            .O(N__42607),
            .I(frame_decoder_CH4data_2));
    CascadeMux I__5893 (
            .O(N__42604),
            .I(N__42601));
    InMux I__5892 (
            .O(N__42601),
            .I(N__42595));
    InMux I__5891 (
            .O(N__42600),
            .I(N__42595));
    LocalMux I__5890 (
            .O(N__42595),
            .I(\scaler_4.un3_source_data_0_cry_1_c_RNI74CL ));
    InMux I__5889 (
            .O(N__42592),
            .I(\scaler_4.un3_source_data_0_cry_1 ));
    InMux I__5888 (
            .O(N__42589),
            .I(N__42586));
    LocalMux I__5887 (
            .O(N__42586),
            .I(frame_decoder_CH4data_3));
    CascadeMux I__5886 (
            .O(N__42583),
            .I(N__42580));
    InMux I__5885 (
            .O(N__42580),
            .I(N__42574));
    InMux I__5884 (
            .O(N__42579),
            .I(N__42574));
    LocalMux I__5883 (
            .O(N__42574),
            .I(\scaler_4.un3_source_data_0_cry_2_c_RNIA8DL ));
    InMux I__5882 (
            .O(N__42571),
            .I(\scaler_4.un3_source_data_0_cry_2 ));
    InMux I__5881 (
            .O(N__42568),
            .I(N__42565));
    LocalMux I__5880 (
            .O(N__42565),
            .I(frame_decoder_CH4data_4));
    CascadeMux I__5879 (
            .O(N__42562),
            .I(N__42559));
    InMux I__5878 (
            .O(N__42559),
            .I(N__42553));
    InMux I__5877 (
            .O(N__42558),
            .I(N__42553));
    LocalMux I__5876 (
            .O(N__42553),
            .I(\scaler_4.un3_source_data_0_cry_3_c_RNIDCEL ));
    InMux I__5875 (
            .O(N__42550),
            .I(\scaler_4.un3_source_data_0_cry_3 ));
    InMux I__5874 (
            .O(N__42547),
            .I(N__42544));
    LocalMux I__5873 (
            .O(N__42544),
            .I(frame_decoder_CH4data_5));
    CascadeMux I__5872 (
            .O(N__42541),
            .I(N__42538));
    InMux I__5871 (
            .O(N__42538),
            .I(N__42532));
    InMux I__5870 (
            .O(N__42537),
            .I(N__42532));
    LocalMux I__5869 (
            .O(N__42532),
            .I(\scaler_4.un3_source_data_0_cry_4_c_RNIGGFL ));
    InMux I__5868 (
            .O(N__42529),
            .I(\scaler_4.un3_source_data_0_cry_4 ));
    InMux I__5867 (
            .O(N__42526),
            .I(N__42523));
    LocalMux I__5866 (
            .O(N__42523),
            .I(frame_decoder_CH4data_6));
    CascadeMux I__5865 (
            .O(N__42520),
            .I(N__42517));
    InMux I__5864 (
            .O(N__42517),
            .I(N__42511));
    InMux I__5863 (
            .O(N__42516),
            .I(N__42511));
    LocalMux I__5862 (
            .O(N__42511),
            .I(\scaler_4.un3_source_data_0_cry_5_c_RNIJKGL ));
    InMux I__5861 (
            .O(N__42508),
            .I(\scaler_4.un3_source_data_0_cry_5 ));
    CascadeMux I__5860 (
            .O(N__42505),
            .I(N__42502));
    InMux I__5859 (
            .O(N__42502),
            .I(N__42496));
    InMux I__5858 (
            .O(N__42501),
            .I(N__42496));
    LocalMux I__5857 (
            .O(N__42496),
            .I(\scaler_4.un3_source_data_0_cry_6_c_RNIOUNN ));
    InMux I__5856 (
            .O(N__42493),
            .I(\scaler_4.un3_source_data_0_cry_6 ));
    InMux I__5855 (
            .O(N__42490),
            .I(N__42486));
    InMux I__5854 (
            .O(N__42489),
            .I(N__42483));
    LocalMux I__5853 (
            .O(N__42486),
            .I(\scaler_4.un3_source_data_0_cry_7_c_RNIP0PN ));
    LocalMux I__5852 (
            .O(N__42483),
            .I(\scaler_4.un3_source_data_0_cry_7_c_RNIP0PN ));
    InMux I__5851 (
            .O(N__42478),
            .I(bfn_8_12_0_));
    InMux I__5850 (
            .O(N__42475),
            .I(N__42471));
    InMux I__5849 (
            .O(N__42474),
            .I(N__42468));
    LocalMux I__5848 (
            .O(N__42471),
            .I(N__42463));
    LocalMux I__5847 (
            .O(N__42468),
            .I(N__42463));
    Odrv4 I__5846 (
            .O(N__42463),
            .I(scaler_4_data_12));
    InMux I__5845 (
            .O(N__42460),
            .I(N__42457));
    LocalMux I__5844 (
            .O(N__42457),
            .I(\ppm_encoder_1.un1_rudder_cry_11_THRU_CO ));
    CascadeMux I__5843 (
            .O(N__42454),
            .I(N__42449));
    InMux I__5842 (
            .O(N__42453),
            .I(N__42444));
    InMux I__5841 (
            .O(N__42452),
            .I(N__42444));
    InMux I__5840 (
            .O(N__42449),
            .I(N__42441));
    LocalMux I__5839 (
            .O(N__42444),
            .I(N__42438));
    LocalMux I__5838 (
            .O(N__42441),
            .I(N__42433));
    Span12Mux_s8_v I__5837 (
            .O(N__42438),
            .I(N__42433));
    Odrv12 I__5836 (
            .O(N__42433),
            .I(\ppm_encoder_1.rudderZ0Z_12 ));
    InMux I__5835 (
            .O(N__42430),
            .I(N__42426));
    CascadeMux I__5834 (
            .O(N__42429),
            .I(N__42423));
    LocalMux I__5833 (
            .O(N__42426),
            .I(N__42420));
    InMux I__5832 (
            .O(N__42423),
            .I(N__42416));
    Span4Mux_h I__5831 (
            .O(N__42420),
            .I(N__42413));
    InMux I__5830 (
            .O(N__42419),
            .I(N__42410));
    LocalMux I__5829 (
            .O(N__42416),
            .I(\ppm_encoder_1.elevatorZ0Z_10 ));
    Odrv4 I__5828 (
            .O(N__42413),
            .I(\ppm_encoder_1.elevatorZ0Z_10 ));
    LocalMux I__5827 (
            .O(N__42410),
            .I(\ppm_encoder_1.elevatorZ0Z_10 ));
    InMux I__5826 (
            .O(N__42403),
            .I(N__42400));
    LocalMux I__5825 (
            .O(N__42400),
            .I(\ppm_encoder_1.un1_rudder_cry_7_THRU_CO ));
    InMux I__5824 (
            .O(N__42397),
            .I(N__42393));
    InMux I__5823 (
            .O(N__42396),
            .I(N__42390));
    LocalMux I__5822 (
            .O(N__42393),
            .I(N__42387));
    LocalMux I__5821 (
            .O(N__42390),
            .I(N__42384));
    Odrv4 I__5820 (
            .O(N__42387),
            .I(scaler_4_data_8));
    Odrv4 I__5819 (
            .O(N__42384),
            .I(scaler_4_data_8));
    CascadeMux I__5818 (
            .O(N__42379),
            .I(N__42375));
    InMux I__5817 (
            .O(N__42378),
            .I(N__42371));
    InMux I__5816 (
            .O(N__42375),
            .I(N__42368));
    CascadeMux I__5815 (
            .O(N__42374),
            .I(N__42365));
    LocalMux I__5814 (
            .O(N__42371),
            .I(N__42362));
    LocalMux I__5813 (
            .O(N__42368),
            .I(N__42359));
    InMux I__5812 (
            .O(N__42365),
            .I(N__42356));
    Span4Mux_v I__5811 (
            .O(N__42362),
            .I(N__42351));
    Span4Mux_v I__5810 (
            .O(N__42359),
            .I(N__42351));
    LocalMux I__5809 (
            .O(N__42356),
            .I(\ppm_encoder_1.elevatorZ0Z_13 ));
    Odrv4 I__5808 (
            .O(N__42351),
            .I(\ppm_encoder_1.elevatorZ0Z_13 ));
    InMux I__5807 (
            .O(N__42346),
            .I(N__42343));
    LocalMux I__5806 (
            .O(N__42343),
            .I(\ppm_encoder_1.un1_rudder_cry_9_THRU_CO ));
    InMux I__5805 (
            .O(N__42340),
            .I(N__42336));
    InMux I__5804 (
            .O(N__42339),
            .I(N__42333));
    LocalMux I__5803 (
            .O(N__42336),
            .I(N__42328));
    LocalMux I__5802 (
            .O(N__42333),
            .I(N__42328));
    Odrv4 I__5801 (
            .O(N__42328),
            .I(scaler_4_data_10));
    InMux I__5800 (
            .O(N__42325),
            .I(N__42322));
    LocalMux I__5799 (
            .O(N__42322),
            .I(\ppm_encoder_1.un1_rudder_cry_12_THRU_CO ));
    InMux I__5798 (
            .O(N__42319),
            .I(N__42316));
    LocalMux I__5797 (
            .O(N__42316),
            .I(N__42312));
    InMux I__5796 (
            .O(N__42315),
            .I(N__42309));
    Span4Mux_h I__5795 (
            .O(N__42312),
            .I(N__42306));
    LocalMux I__5794 (
            .O(N__42309),
            .I(N__42303));
    Odrv4 I__5793 (
            .O(N__42306),
            .I(scaler_4_data_13));
    Odrv4 I__5792 (
            .O(N__42303),
            .I(scaler_4_data_13));
    InMux I__5791 (
            .O(N__42298),
            .I(N__42294));
    CascadeMux I__5790 (
            .O(N__42297),
            .I(N__42291));
    LocalMux I__5789 (
            .O(N__42294),
            .I(N__42288));
    InMux I__5788 (
            .O(N__42291),
            .I(N__42285));
    Span4Mux_v I__5787 (
            .O(N__42288),
            .I(N__42282));
    LocalMux I__5786 (
            .O(N__42285),
            .I(\ppm_encoder_1.rudderZ0Z_13 ));
    Odrv4 I__5785 (
            .O(N__42282),
            .I(\ppm_encoder_1.rudderZ0Z_13 ));
    InMux I__5784 (
            .O(N__42277),
            .I(N__42274));
    LocalMux I__5783 (
            .O(N__42274),
            .I(\ppm_encoder_1.N_266_i ));
    InMux I__5782 (
            .O(N__42271),
            .I(N__42266));
    InMux I__5781 (
            .O(N__42270),
            .I(N__42261));
    InMux I__5780 (
            .O(N__42269),
            .I(N__42261));
    LocalMux I__5779 (
            .O(N__42266),
            .I(\ppm_encoder_1.aileronZ0Z_0 ));
    LocalMux I__5778 (
            .O(N__42261),
            .I(\ppm_encoder_1.aileronZ0Z_0 ));
    CascadeMux I__5777 (
            .O(N__42256),
            .I(N__42252));
    CascadeMux I__5776 (
            .O(N__42255),
            .I(N__42248));
    InMux I__5775 (
            .O(N__42252),
            .I(N__42245));
    InMux I__5774 (
            .O(N__42251),
            .I(N__42240));
    InMux I__5773 (
            .O(N__42248),
            .I(N__42240));
    LocalMux I__5772 (
            .O(N__42245),
            .I(\ppm_encoder_1.throttleZ0Z_0 ));
    LocalMux I__5771 (
            .O(N__42240),
            .I(\ppm_encoder_1.throttleZ0Z_0 ));
    CascadeMux I__5770 (
            .O(N__42235),
            .I(N__42231));
    CascadeMux I__5769 (
            .O(N__42234),
            .I(N__42228));
    InMux I__5768 (
            .O(N__42231),
            .I(N__42225));
    InMux I__5767 (
            .O(N__42228),
            .I(N__42221));
    LocalMux I__5766 (
            .O(N__42225),
            .I(N__42218));
    InMux I__5765 (
            .O(N__42224),
            .I(N__42215));
    LocalMux I__5764 (
            .O(N__42221),
            .I(\ppm_encoder_1.aileronZ0Z_10 ));
    Odrv4 I__5763 (
            .O(N__42218),
            .I(\ppm_encoder_1.aileronZ0Z_10 ));
    LocalMux I__5762 (
            .O(N__42215),
            .I(\ppm_encoder_1.aileronZ0Z_10 ));
    InMux I__5761 (
            .O(N__42208),
            .I(N__42199));
    InMux I__5760 (
            .O(N__42207),
            .I(N__42199));
    CascadeMux I__5759 (
            .O(N__42206),
            .I(N__42194));
    InMux I__5758 (
            .O(N__42205),
            .I(N__42189));
    InMux I__5757 (
            .O(N__42204),
            .I(N__42186));
    LocalMux I__5756 (
            .O(N__42199),
            .I(N__42183));
    InMux I__5755 (
            .O(N__42198),
            .I(N__42180));
    InMux I__5754 (
            .O(N__42197),
            .I(N__42176));
    InMux I__5753 (
            .O(N__42194),
            .I(N__42173));
    CascadeMux I__5752 (
            .O(N__42193),
            .I(N__42167));
    CascadeMux I__5751 (
            .O(N__42192),
            .I(N__42163));
    LocalMux I__5750 (
            .O(N__42189),
            .I(N__42157));
    LocalMux I__5749 (
            .O(N__42186),
            .I(N__42157));
    Span4Mux_v I__5748 (
            .O(N__42183),
            .I(N__42150));
    LocalMux I__5747 (
            .O(N__42180),
            .I(N__42150));
    InMux I__5746 (
            .O(N__42179),
            .I(N__42147));
    LocalMux I__5745 (
            .O(N__42176),
            .I(N__42144));
    LocalMux I__5744 (
            .O(N__42173),
            .I(N__42141));
    InMux I__5743 (
            .O(N__42172),
            .I(N__42138));
    InMux I__5742 (
            .O(N__42171),
            .I(N__42135));
    InMux I__5741 (
            .O(N__42170),
            .I(N__42132));
    InMux I__5740 (
            .O(N__42167),
            .I(N__42123));
    InMux I__5739 (
            .O(N__42166),
            .I(N__42123));
    InMux I__5738 (
            .O(N__42163),
            .I(N__42123));
    InMux I__5737 (
            .O(N__42162),
            .I(N__42123));
    Span4Mux_h I__5736 (
            .O(N__42157),
            .I(N__42120));
    InMux I__5735 (
            .O(N__42156),
            .I(N__42115));
    InMux I__5734 (
            .O(N__42155),
            .I(N__42115));
    Span4Mux_h I__5733 (
            .O(N__42150),
            .I(N__42106));
    LocalMux I__5732 (
            .O(N__42147),
            .I(N__42106));
    Span4Mux_s2_v I__5731 (
            .O(N__42144),
            .I(N__42106));
    Span4Mux_s2_v I__5730 (
            .O(N__42141),
            .I(N__42106));
    LocalMux I__5729 (
            .O(N__42138),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1 ));
    LocalMux I__5728 (
            .O(N__42135),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1 ));
    LocalMux I__5727 (
            .O(N__42132),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1 ));
    LocalMux I__5726 (
            .O(N__42123),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1 ));
    Odrv4 I__5725 (
            .O(N__42120),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1 ));
    LocalMux I__5724 (
            .O(N__42115),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1 ));
    Odrv4 I__5723 (
            .O(N__42106),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1 ));
    InMux I__5722 (
            .O(N__42091),
            .I(N__42084));
    InMux I__5721 (
            .O(N__42090),
            .I(N__42084));
    InMux I__5720 (
            .O(N__42089),
            .I(N__42081));
    LocalMux I__5719 (
            .O(N__42084),
            .I(N__42075));
    LocalMux I__5718 (
            .O(N__42081),
            .I(N__42072));
    CascadeMux I__5717 (
            .O(N__42080),
            .I(N__42068));
    InMux I__5716 (
            .O(N__42079),
            .I(N__42064));
    InMux I__5715 (
            .O(N__42078),
            .I(N__42061));
    Span4Mux_h I__5714 (
            .O(N__42075),
            .I(N__42056));
    Span4Mux_v I__5713 (
            .O(N__42072),
            .I(N__42056));
    InMux I__5712 (
            .O(N__42071),
            .I(N__42049));
    InMux I__5711 (
            .O(N__42068),
            .I(N__42049));
    InMux I__5710 (
            .O(N__42067),
            .I(N__42049));
    LocalMux I__5709 (
            .O(N__42064),
            .I(N__42044));
    LocalMux I__5708 (
            .O(N__42061),
            .I(N__42044));
    Odrv4 I__5707 (
            .O(N__42056),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ));
    LocalMux I__5706 (
            .O(N__42049),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ));
    Odrv4 I__5705 (
            .O(N__42044),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ));
    CascadeMux I__5704 (
            .O(N__42037),
            .I(\ppm_encoder_1.N_508_cascade_ ));
    InMux I__5703 (
            .O(N__42034),
            .I(N__42031));
    LocalMux I__5702 (
            .O(N__42031),
            .I(N__42028));
    Span4Mux_h I__5701 (
            .O(N__42028),
            .I(N__42024));
    InMux I__5700 (
            .O(N__42027),
            .I(N__42021));
    Odrv4 I__5699 (
            .O(N__42024),
            .I(throttle_order_12));
    LocalMux I__5698 (
            .O(N__42021),
            .I(throttle_order_12));
    InMux I__5697 (
            .O(N__42016),
            .I(N__42013));
    LocalMux I__5696 (
            .O(N__42013),
            .I(N__42010));
    Span4Mux_v I__5695 (
            .O(N__42010),
            .I(N__42007));
    Odrv4 I__5694 (
            .O(N__42007),
            .I(\ppm_encoder_1.un1_throttle_cry_11_THRU_CO ));
    InMux I__5693 (
            .O(N__42004),
            .I(N__42001));
    LocalMux I__5692 (
            .O(N__42001),
            .I(N__41998));
    Odrv4 I__5691 (
            .O(N__41998),
            .I(\ppm_encoder_1.un1_init_pulses_11_15 ));
    InMux I__5690 (
            .O(N__41995),
            .I(N__41992));
    LocalMux I__5689 (
            .O(N__41992),
            .I(N__41989));
    Span4Mux_v I__5688 (
            .O(N__41989),
            .I(N__41985));
    CascadeMux I__5687 (
            .O(N__41988),
            .I(N__41979));
    Span4Mux_h I__5686 (
            .O(N__41985),
            .I(N__41976));
    InMux I__5685 (
            .O(N__41984),
            .I(N__41971));
    InMux I__5684 (
            .O(N__41983),
            .I(N__41971));
    InMux I__5683 (
            .O(N__41982),
            .I(N__41966));
    InMux I__5682 (
            .O(N__41979),
            .I(N__41966));
    Odrv4 I__5681 (
            .O(N__41976),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3 ));
    LocalMux I__5680 (
            .O(N__41971),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3 ));
    LocalMux I__5679 (
            .O(N__41966),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3 ));
    CascadeMux I__5678 (
            .O(N__41959),
            .I(\ppm_encoder_1.N_257_i_i_cascade_ ));
    InMux I__5677 (
            .O(N__41956),
            .I(N__41953));
    LocalMux I__5676 (
            .O(N__41953),
            .I(N__41950));
    Span4Mux_h I__5675 (
            .O(N__41950),
            .I(N__41946));
    InMux I__5674 (
            .O(N__41949),
            .I(N__41943));
    Span4Mux_v I__5673 (
            .O(N__41946),
            .I(N__41940));
    LocalMux I__5672 (
            .O(N__41943),
            .I(N__41937));
    Odrv4 I__5671 (
            .O(N__41940),
            .I(throttle_order_0));
    Odrv4 I__5670 (
            .O(N__41937),
            .I(throttle_order_0));
    CascadeMux I__5669 (
            .O(N__41932),
            .I(\ppm_encoder_1.N_254_i_i_cascade_ ));
    InMux I__5668 (
            .O(N__41929),
            .I(N__41926));
    LocalMux I__5667 (
            .O(N__41926),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_17 ));
    CascadeMux I__5666 (
            .O(N__41923),
            .I(N__41920));
    InMux I__5665 (
            .O(N__41920),
            .I(N__41917));
    LocalMux I__5664 (
            .O(N__41917),
            .I(\ppm_encoder_1.un1_init_pulses_11_16 ));
    InMux I__5663 (
            .O(N__41914),
            .I(N__41911));
    LocalMux I__5662 (
            .O(N__41911),
            .I(N__41908));
    Odrv4 I__5661 (
            .O(N__41908),
            .I(\ppm_encoder_1.un1_init_pulses_11_10 ));
    CascadeMux I__5660 (
            .O(N__41905),
            .I(\ppm_encoder_1.N_298_cascade_ ));
    InMux I__5659 (
            .O(N__41902),
            .I(N__41899));
    LocalMux I__5658 (
            .O(N__41899),
            .I(\ppm_encoder_1.un1_init_pulses_11_17 ));
    InMux I__5657 (
            .O(N__41896),
            .I(N__41893));
    LocalMux I__5656 (
            .O(N__41893),
            .I(\ppm_encoder_1.un1_init_pulses_11_18 ));
    InMux I__5655 (
            .O(N__41890),
            .I(N__41887));
    LocalMux I__5654 (
            .O(N__41887),
            .I(N__41884));
    Odrv4 I__5653 (
            .O(N__41884),
            .I(\ppm_encoder_1.un1_init_pulses_11_13 ));
    InMux I__5652 (
            .O(N__41881),
            .I(N__41877));
    CascadeMux I__5651 (
            .O(N__41880),
            .I(N__41874));
    LocalMux I__5650 (
            .O(N__41877),
            .I(N__41870));
    InMux I__5649 (
            .O(N__41874),
            .I(N__41867));
    CascadeMux I__5648 (
            .O(N__41873),
            .I(N__41864));
    Span4Mux_v I__5647 (
            .O(N__41870),
            .I(N__41859));
    LocalMux I__5646 (
            .O(N__41867),
            .I(N__41859));
    InMux I__5645 (
            .O(N__41864),
            .I(N__41855));
    Span4Mux_h I__5644 (
            .O(N__41859),
            .I(N__41852));
    InMux I__5643 (
            .O(N__41858),
            .I(N__41849));
    LocalMux I__5642 (
            .O(N__41855),
            .I(\ppm_encoder_1.init_pulsesZ0Z_13 ));
    Odrv4 I__5641 (
            .O(N__41852),
            .I(\ppm_encoder_1.init_pulsesZ0Z_13 ));
    LocalMux I__5640 (
            .O(N__41849),
            .I(\ppm_encoder_1.init_pulsesZ0Z_13 ));
    CascadeMux I__5639 (
            .O(N__41842),
            .I(N__41839));
    InMux I__5638 (
            .O(N__41839),
            .I(N__41836));
    LocalMux I__5637 (
            .O(N__41836),
            .I(N__41833));
    Odrv12 I__5636 (
            .O(N__41833),
            .I(\ppm_encoder_1.un1_init_pulses_11_14 ));
    CascadeMux I__5635 (
            .O(N__41830),
            .I(N__41827));
    InMux I__5634 (
            .O(N__41827),
            .I(N__41824));
    LocalMux I__5633 (
            .O(N__41824),
            .I(\ppm_encoder_1.init_pulses_RNIOHJF3Z0Z_13 ));
    InMux I__5632 (
            .O(N__41821),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_12 ));
    InMux I__5631 (
            .O(N__41818),
            .I(N__41815));
    LocalMux I__5630 (
            .O(N__41815),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_14 ));
    InMux I__5629 (
            .O(N__41812),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_13 ));
    InMux I__5628 (
            .O(N__41809),
            .I(N__41806));
    LocalMux I__5627 (
            .O(N__41806),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_15 ));
    InMux I__5626 (
            .O(N__41803),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_14 ));
    InMux I__5625 (
            .O(N__41800),
            .I(bfn_8_3_0_));
    InMux I__5624 (
            .O(N__41797),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_16 ));
    InMux I__5623 (
            .O(N__41794),
            .I(N__41791));
    LocalMux I__5622 (
            .O(N__41791),
            .I(N__41783));
    InMux I__5621 (
            .O(N__41790),
            .I(N__41780));
    InMux I__5620 (
            .O(N__41789),
            .I(N__41777));
    InMux I__5619 (
            .O(N__41788),
            .I(N__41773));
    InMux I__5618 (
            .O(N__41787),
            .I(N__41766));
    InMux I__5617 (
            .O(N__41786),
            .I(N__41766));
    Span4Mux_v I__5616 (
            .O(N__41783),
            .I(N__41761));
    LocalMux I__5615 (
            .O(N__41780),
            .I(N__41761));
    LocalMux I__5614 (
            .O(N__41777),
            .I(N__41755));
    InMux I__5613 (
            .O(N__41776),
            .I(N__41752));
    LocalMux I__5612 (
            .O(N__41773),
            .I(N__41749));
    InMux I__5611 (
            .O(N__41772),
            .I(N__41744));
    InMux I__5610 (
            .O(N__41771),
            .I(N__41744));
    LocalMux I__5609 (
            .O(N__41766),
            .I(N__41741));
    Span4Mux_h I__5608 (
            .O(N__41761),
            .I(N__41738));
    InMux I__5607 (
            .O(N__41760),
            .I(N__41735));
    InMux I__5606 (
            .O(N__41759),
            .I(N__41732));
    InMux I__5605 (
            .O(N__41758),
            .I(N__41729));
    Span4Mux_h I__5604 (
            .O(N__41755),
            .I(N__41722));
    LocalMux I__5603 (
            .O(N__41752),
            .I(N__41722));
    Span4Mux_s2_v I__5602 (
            .O(N__41749),
            .I(N__41722));
    LocalMux I__5601 (
            .O(N__41744),
            .I(N__41717));
    Span4Mux_s1_v I__5600 (
            .O(N__41741),
            .I(N__41717));
    Odrv4 I__5599 (
            .O(N__41738),
            .I(\ppm_encoder_1.PPM_STATE_RNIMINSZ0Z_0 ));
    LocalMux I__5598 (
            .O(N__41735),
            .I(\ppm_encoder_1.PPM_STATE_RNIMINSZ0Z_0 ));
    LocalMux I__5597 (
            .O(N__41732),
            .I(\ppm_encoder_1.PPM_STATE_RNIMINSZ0Z_0 ));
    LocalMux I__5596 (
            .O(N__41729),
            .I(\ppm_encoder_1.PPM_STATE_RNIMINSZ0Z_0 ));
    Odrv4 I__5595 (
            .O(N__41722),
            .I(\ppm_encoder_1.PPM_STATE_RNIMINSZ0Z_0 ));
    Odrv4 I__5594 (
            .O(N__41717),
            .I(\ppm_encoder_1.PPM_STATE_RNIMINSZ0Z_0 ));
    InMux I__5593 (
            .O(N__41704),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_17 ));
    InMux I__5592 (
            .O(N__41701),
            .I(N__41698));
    LocalMux I__5591 (
            .O(N__41698),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_11 ));
    InMux I__5590 (
            .O(N__41695),
            .I(N__41692));
    LocalMux I__5589 (
            .O(N__41692),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_13 ));
    InMux I__5588 (
            .O(N__41689),
            .I(N__41686));
    LocalMux I__5587 (
            .O(N__41686),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_5 ));
    InMux I__5586 (
            .O(N__41683),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_4 ));
    InMux I__5585 (
            .O(N__41680),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_5 ));
    InMux I__5584 (
            .O(N__41677),
            .I(N__41674));
    LocalMux I__5583 (
            .O(N__41674),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_7 ));
    InMux I__5582 (
            .O(N__41671),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_6 ));
    InMux I__5581 (
            .O(N__41668),
            .I(N__41665));
    LocalMux I__5580 (
            .O(N__41665),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_8 ));
    InMux I__5579 (
            .O(N__41662),
            .I(bfn_8_2_0_));
    InMux I__5578 (
            .O(N__41659),
            .I(N__41656));
    LocalMux I__5577 (
            .O(N__41656),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_9 ));
    InMux I__5576 (
            .O(N__41653),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_8 ));
    InMux I__5575 (
            .O(N__41650),
            .I(N__41647));
    LocalMux I__5574 (
            .O(N__41647),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_10 ));
    InMux I__5573 (
            .O(N__41644),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_9 ));
    InMux I__5572 (
            .O(N__41641),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_10 ));
    InMux I__5571 (
            .O(N__41638),
            .I(N__41635));
    LocalMux I__5570 (
            .O(N__41635),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_12 ));
    InMux I__5569 (
            .O(N__41632),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_11 ));
    InMux I__5568 (
            .O(N__41629),
            .I(N__41624));
    CascadeMux I__5567 (
            .O(N__41628),
            .I(N__41620));
    InMux I__5566 (
            .O(N__41627),
            .I(N__41617));
    LocalMux I__5565 (
            .O(N__41624),
            .I(N__41614));
    InMux I__5564 (
            .O(N__41623),
            .I(N__41611));
    InMux I__5563 (
            .O(N__41620),
            .I(N__41608));
    LocalMux I__5562 (
            .O(N__41617),
            .I(N__41601));
    Span12Mux_v I__5561 (
            .O(N__41614),
            .I(N__41601));
    LocalMux I__5560 (
            .O(N__41611),
            .I(N__41601));
    LocalMux I__5559 (
            .O(N__41608),
            .I(\Commands_frame_decoder.countZ0Z_0 ));
    Odrv12 I__5558 (
            .O(N__41601),
            .I(\Commands_frame_decoder.countZ0Z_0 ));
    InMux I__5557 (
            .O(N__41596),
            .I(N__41593));
    LocalMux I__5556 (
            .O(N__41593),
            .I(N__41590));
    Span4Mux_v I__5555 (
            .O(N__41590),
            .I(N__41587));
    Odrv4 I__5554 (
            .O(N__41587),
            .I(\uart_pc.N_144_1 ));
    CascadeMux I__5553 (
            .O(N__41584),
            .I(N__41580));
    InMux I__5552 (
            .O(N__41583),
            .I(N__41574));
    InMux I__5551 (
            .O(N__41580),
            .I(N__41574));
    InMux I__5550 (
            .O(N__41579),
            .I(N__41568));
    LocalMux I__5549 (
            .O(N__41574),
            .I(N__41565));
    InMux I__5548 (
            .O(N__41573),
            .I(N__41558));
    InMux I__5547 (
            .O(N__41572),
            .I(N__41558));
    InMux I__5546 (
            .O(N__41571),
            .I(N__41558));
    LocalMux I__5545 (
            .O(N__41568),
            .I(\uart_pc.N_143 ));
    Odrv4 I__5544 (
            .O(N__41565),
            .I(\uart_pc.N_143 ));
    LocalMux I__5543 (
            .O(N__41558),
            .I(\uart_pc.N_143 ));
    CascadeMux I__5542 (
            .O(N__41551),
            .I(N__41548));
    InMux I__5541 (
            .O(N__41548),
            .I(N__41544));
    InMux I__5540 (
            .O(N__41547),
            .I(N__41541));
    LocalMux I__5539 (
            .O(N__41544),
            .I(N__41538));
    LocalMux I__5538 (
            .O(N__41541),
            .I(\Commands_frame_decoder.stateZ0Z_0 ));
    Odrv12 I__5537 (
            .O(N__41538),
            .I(\Commands_frame_decoder.stateZ0Z_0 ));
    CascadeMux I__5536 (
            .O(N__41533),
            .I(N__41530));
    InMux I__5535 (
            .O(N__41530),
            .I(N__41527));
    LocalMux I__5534 (
            .O(N__41527),
            .I(N__41524));
    Span4Mux_v I__5533 (
            .O(N__41524),
            .I(N__41521));
    Odrv4 I__5532 (
            .O(N__41521),
            .I(\Commands_frame_decoder.state_ns_0_a3_3_1 ));
    IoInMux I__5531 (
            .O(N__41518),
            .I(N__41515));
    LocalMux I__5530 (
            .O(N__41515),
            .I(N__41512));
    Span4Mux_s1_v I__5529 (
            .O(N__41512),
            .I(N__41509));
    Span4Mux_v I__5528 (
            .O(N__41509),
            .I(N__41506));
    Odrv4 I__5527 (
            .O(N__41506),
            .I(\pid_front.state_0_0 ));
    CascadeMux I__5526 (
            .O(N__41503),
            .I(N__41500));
    InMux I__5525 (
            .O(N__41500),
            .I(N__41497));
    LocalMux I__5524 (
            .O(N__41497),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5I0L2Z0Z_3 ));
    InMux I__5523 (
            .O(N__41494),
            .I(N__41491));
    LocalMux I__5522 (
            .O(N__41491),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_1 ));
    InMux I__5521 (
            .O(N__41488),
            .I(N__41485));
    LocalMux I__5520 (
            .O(N__41485),
            .I(N__41482));
    Span4Mux_h I__5519 (
            .O(N__41482),
            .I(N__41479));
    Odrv4 I__5518 (
            .O(N__41479),
            .I(\ppm_encoder_1.un1_init_pulses_11_1 ));
    InMux I__5517 (
            .O(N__41476),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_0 ));
    CascadeMux I__5516 (
            .O(N__41473),
            .I(N__41470));
    InMux I__5515 (
            .O(N__41470),
            .I(N__41467));
    LocalMux I__5514 (
            .O(N__41467),
            .I(N__41464));
    Span4Mux_s2_v I__5513 (
            .O(N__41464),
            .I(N__41461));
    Odrv4 I__5512 (
            .O(N__41461),
            .I(\ppm_encoder_1.init_pulses_RNIHGIP3Z0Z_2 ));
    InMux I__5511 (
            .O(N__41458),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_1 ));
    InMux I__5510 (
            .O(N__41455),
            .I(N__41452));
    LocalMux I__5509 (
            .O(N__41452),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_3 ));
    InMux I__5508 (
            .O(N__41449),
            .I(N__41446));
    LocalMux I__5507 (
            .O(N__41446),
            .I(N__41443));
    Span4Mux_v I__5506 (
            .O(N__41443),
            .I(N__41440));
    Odrv4 I__5505 (
            .O(N__41440),
            .I(\ppm_encoder_1.un1_init_pulses_11_3 ));
    InMux I__5504 (
            .O(N__41437),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_2 ));
    InMux I__5503 (
            .O(N__41434),
            .I(N__41431));
    LocalMux I__5502 (
            .O(N__41431),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_4 ));
    InMux I__5501 (
            .O(N__41428),
            .I(N__41425));
    LocalMux I__5500 (
            .O(N__41425),
            .I(N__41422));
    Span4Mux_v I__5499 (
            .O(N__41422),
            .I(N__41419));
    Odrv4 I__5498 (
            .O(N__41419),
            .I(\ppm_encoder_1.un1_init_pulses_11_4 ));
    InMux I__5497 (
            .O(N__41416),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_3 ));
    InMux I__5496 (
            .O(N__41413),
            .I(\uart_pc.un4_timer_Count_1_cry_2 ));
    InMux I__5495 (
            .O(N__41410),
            .I(\uart_pc.un4_timer_Count_1_cry_3 ));
    InMux I__5494 (
            .O(N__41407),
            .I(N__41404));
    LocalMux I__5493 (
            .O(N__41404),
            .I(\uart_pc.timer_Count_RNO_0Z0Z_4 ));
    InMux I__5492 (
            .O(N__41401),
            .I(N__41392));
    InMux I__5491 (
            .O(N__41400),
            .I(N__41379));
    InMux I__5490 (
            .O(N__41399),
            .I(N__41379));
    InMux I__5489 (
            .O(N__41398),
            .I(N__41379));
    InMux I__5488 (
            .O(N__41397),
            .I(N__41379));
    InMux I__5487 (
            .O(N__41396),
            .I(N__41379));
    InMux I__5486 (
            .O(N__41395),
            .I(N__41376));
    LocalMux I__5485 (
            .O(N__41392),
            .I(N__41373));
    InMux I__5484 (
            .O(N__41391),
            .I(N__41368));
    InMux I__5483 (
            .O(N__41390),
            .I(N__41368));
    LocalMux I__5482 (
            .O(N__41379),
            .I(N__41365));
    LocalMux I__5481 (
            .O(N__41376),
            .I(\uart_pc.timer_CountZ0Z_4 ));
    Odrv4 I__5480 (
            .O(N__41373),
            .I(\uart_pc.timer_CountZ0Z_4 ));
    LocalMux I__5479 (
            .O(N__41368),
            .I(\uart_pc.timer_CountZ0Z_4 ));
    Odrv12 I__5478 (
            .O(N__41365),
            .I(\uart_pc.timer_CountZ0Z_4 ));
    InMux I__5477 (
            .O(N__41356),
            .I(N__41353));
    LocalMux I__5476 (
            .O(N__41353),
            .I(\uart_pc.timer_Count_RNO_0Z0Z_3 ));
    CascadeMux I__5475 (
            .O(N__41350),
            .I(N__41343));
    InMux I__5474 (
            .O(N__41349),
            .I(N__41332));
    InMux I__5473 (
            .O(N__41348),
            .I(N__41332));
    InMux I__5472 (
            .O(N__41347),
            .I(N__41332));
    InMux I__5471 (
            .O(N__41346),
            .I(N__41332));
    InMux I__5470 (
            .O(N__41343),
            .I(N__41332));
    LocalMux I__5469 (
            .O(N__41332),
            .I(N__41326));
    InMux I__5468 (
            .O(N__41331),
            .I(N__41321));
    InMux I__5467 (
            .O(N__41330),
            .I(N__41321));
    InMux I__5466 (
            .O(N__41329),
            .I(N__41318));
    Span4Mux_v I__5465 (
            .O(N__41326),
            .I(N__41313));
    LocalMux I__5464 (
            .O(N__41321),
            .I(N__41313));
    LocalMux I__5463 (
            .O(N__41318),
            .I(\uart_pc.timer_CountZ1Z_3 ));
    Odrv4 I__5462 (
            .O(N__41313),
            .I(\uart_pc.timer_CountZ1Z_3 ));
    CascadeMux I__5461 (
            .O(N__41308),
            .I(N__41302));
    InMux I__5460 (
            .O(N__41307),
            .I(N__41299));
    InMux I__5459 (
            .O(N__41306),
            .I(N__41292));
    InMux I__5458 (
            .O(N__41305),
            .I(N__41292));
    InMux I__5457 (
            .O(N__41302),
            .I(N__41292));
    LocalMux I__5456 (
            .O(N__41299),
            .I(\uart_pc.timer_CountZ0Z_0 ));
    LocalMux I__5455 (
            .O(N__41292),
            .I(\uart_pc.timer_CountZ0Z_0 ));
    InMux I__5454 (
            .O(N__41287),
            .I(N__41280));
    CascadeMux I__5453 (
            .O(N__41286),
            .I(N__41277));
    CascadeMux I__5452 (
            .O(N__41285),
            .I(N__41274));
    CascadeMux I__5451 (
            .O(N__41284),
            .I(N__41271));
    CascadeMux I__5450 (
            .O(N__41283),
            .I(N__41268));
    LocalMux I__5449 (
            .O(N__41280),
            .I(N__41265));
    InMux I__5448 (
            .O(N__41277),
            .I(N__41262));
    InMux I__5447 (
            .O(N__41274),
            .I(N__41257));
    InMux I__5446 (
            .O(N__41271),
            .I(N__41257));
    InMux I__5445 (
            .O(N__41268),
            .I(N__41254));
    Span4Mux_v I__5444 (
            .O(N__41265),
            .I(N__41245));
    LocalMux I__5443 (
            .O(N__41262),
            .I(N__41245));
    LocalMux I__5442 (
            .O(N__41257),
            .I(N__41245));
    LocalMux I__5441 (
            .O(N__41254),
            .I(N__41245));
    Odrv4 I__5440 (
            .O(N__41245),
            .I(\uart_pc.timer_Count_0_sqmuxa ));
    CascadeMux I__5439 (
            .O(N__41242),
            .I(\uart_pc.timer_Count_RNO_0Z0Z_1_cascade_ ));
    InMux I__5438 (
            .O(N__41239),
            .I(N__41235));
    InMux I__5437 (
            .O(N__41238),
            .I(N__41232));
    LocalMux I__5436 (
            .O(N__41235),
            .I(\uart_pc.timer_CountZ1Z_1 ));
    LocalMux I__5435 (
            .O(N__41232),
            .I(\uart_pc.timer_CountZ1Z_1 ));
    InMux I__5434 (
            .O(N__41227),
            .I(N__41223));
    InMux I__5433 (
            .O(N__41226),
            .I(N__41220));
    LocalMux I__5432 (
            .O(N__41223),
            .I(N__41212));
    LocalMux I__5431 (
            .O(N__41220),
            .I(N__41212));
    InMux I__5430 (
            .O(N__41219),
            .I(N__41209));
    InMux I__5429 (
            .O(N__41218),
            .I(N__41204));
    InMux I__5428 (
            .O(N__41217),
            .I(N__41204));
    Odrv12 I__5427 (
            .O(N__41212),
            .I(\Commands_frame_decoder.stateZ0Z_14 ));
    LocalMux I__5426 (
            .O(N__41209),
            .I(\Commands_frame_decoder.stateZ0Z_14 ));
    LocalMux I__5425 (
            .O(N__41204),
            .I(\Commands_frame_decoder.stateZ0Z_14 ));
    CascadeMux I__5424 (
            .O(N__41197),
            .I(N__41194));
    InMux I__5423 (
            .O(N__41194),
            .I(N__41188));
    InMux I__5422 (
            .O(N__41193),
            .I(N__41188));
    LocalMux I__5421 (
            .O(N__41188),
            .I(\Commands_frame_decoder.stateZ0Z_2 ));
    CascadeMux I__5420 (
            .O(N__41185),
            .I(\uart_pc.state_srsts_0_0_0_cascade_ ));
    CascadeMux I__5419 (
            .O(N__41182),
            .I(N__41179));
    InMux I__5418 (
            .O(N__41179),
            .I(N__41176));
    LocalMux I__5417 (
            .O(N__41176),
            .I(N__41173));
    Span4Mux_h I__5416 (
            .O(N__41173),
            .I(N__41169));
    InMux I__5415 (
            .O(N__41172),
            .I(N__41166));
    Odrv4 I__5414 (
            .O(N__41169),
            .I(\uart_pc.stateZ0Z_0 ));
    LocalMux I__5413 (
            .O(N__41166),
            .I(\uart_pc.stateZ0Z_0 ));
    CascadeMux I__5412 (
            .O(N__41161),
            .I(\uart_pc.N_126_li_cascade_ ));
    CascadeMux I__5411 (
            .O(N__41158),
            .I(N__41153));
    CascadeMux I__5410 (
            .O(N__41157),
            .I(N__41150));
    InMux I__5409 (
            .O(N__41156),
            .I(N__41147));
    InMux I__5408 (
            .O(N__41153),
            .I(N__41142));
    InMux I__5407 (
            .O(N__41150),
            .I(N__41142));
    LocalMux I__5406 (
            .O(N__41147),
            .I(\uart_pc.timer_CountZ1Z_2 ));
    LocalMux I__5405 (
            .O(N__41142),
            .I(\uart_pc.timer_CountZ1Z_2 ));
    InMux I__5404 (
            .O(N__41137),
            .I(N__41134));
    LocalMux I__5403 (
            .O(N__41134),
            .I(\uart_pc.timer_Count_RNO_0Z0Z_2 ));
    InMux I__5402 (
            .O(N__41131),
            .I(\uart_pc.un4_timer_Count_1_cry_1 ));
    InMux I__5401 (
            .O(N__41128),
            .I(N__41125));
    LocalMux I__5400 (
            .O(N__41125),
            .I(N__41122));
    Odrv12 I__5399 (
            .O(N__41122),
            .I(\Commands_frame_decoder.count_1_sqmuxa ));
    CascadeMux I__5398 (
            .O(N__41119),
            .I(N__41113));
    InMux I__5397 (
            .O(N__41118),
            .I(N__41108));
    InMux I__5396 (
            .O(N__41117),
            .I(N__41108));
    InMux I__5395 (
            .O(N__41116),
            .I(N__41103));
    InMux I__5394 (
            .O(N__41113),
            .I(N__41103));
    LocalMux I__5393 (
            .O(N__41108),
            .I(\uart_pc.stateZ0Z_2 ));
    LocalMux I__5392 (
            .O(N__41103),
            .I(\uart_pc.stateZ0Z_2 ));
    InMux I__5391 (
            .O(N__41098),
            .I(N__41095));
    LocalMux I__5390 (
            .O(N__41095),
            .I(\uart_pc.N_145 ));
    InMux I__5389 (
            .O(N__41092),
            .I(N__41089));
    LocalMux I__5388 (
            .O(N__41089),
            .I(N__41086));
    Odrv12 I__5387 (
            .O(N__41086),
            .I(\Commands_frame_decoder.N_370_2 ));
    InMux I__5386 (
            .O(N__41083),
            .I(N__41080));
    LocalMux I__5385 (
            .O(N__41080),
            .I(N__41077));
    Odrv4 I__5384 (
            .O(N__41077),
            .I(\Commands_frame_decoder.N_371 ));
    CascadeMux I__5383 (
            .O(N__41074),
            .I(\Commands_frame_decoder.N_370_2_cascade_ ));
    CascadeMux I__5382 (
            .O(N__41071),
            .I(\Commands_frame_decoder.state_ns_i_0_0_cascade_ ));
    InMux I__5381 (
            .O(N__41068),
            .I(N__41065));
    LocalMux I__5380 (
            .O(N__41065),
            .I(N__41062));
    Odrv4 I__5379 (
            .O(N__41062),
            .I(\Commands_frame_decoder.N_372 ));
    CascadeMux I__5378 (
            .O(N__41059),
            .I(\Commands_frame_decoder.state_RNO_0Z0Z_14_cascade_ ));
    InMux I__5377 (
            .O(N__41056),
            .I(N__41050));
    InMux I__5376 (
            .O(N__41055),
            .I(N__41050));
    LocalMux I__5375 (
            .O(N__41050),
            .I(N__41047));
    Odrv4 I__5374 (
            .O(N__41047),
            .I(\Commands_frame_decoder.N_365_0 ));
    CascadeMux I__5373 (
            .O(N__41044),
            .I(\Commands_frame_decoder.N_365_0_cascade_ ));
    InMux I__5372 (
            .O(N__41041),
            .I(N__41038));
    LocalMux I__5371 (
            .O(N__41038),
            .I(\Commands_frame_decoder.WDT_RNITK4LZ0Z_8 ));
    InMux I__5370 (
            .O(N__41035),
            .I(N__41032));
    LocalMux I__5369 (
            .O(N__41032),
            .I(N__41029));
    Span4Mux_v I__5368 (
            .O(N__41029),
            .I(N__41026));
    Span4Mux_h I__5367 (
            .O(N__41026),
            .I(N__41023));
    Odrv4 I__5366 (
            .O(N__41023),
            .I(\pid_front.O_0_13 ));
    CascadeMux I__5365 (
            .O(N__41020),
            .I(N__41015));
    InMux I__5364 (
            .O(N__41019),
            .I(N__41012));
    InMux I__5363 (
            .O(N__41018),
            .I(N__41007));
    InMux I__5362 (
            .O(N__41015),
            .I(N__41007));
    LocalMux I__5361 (
            .O(N__41012),
            .I(N__41002));
    LocalMux I__5360 (
            .O(N__41007),
            .I(N__41002));
    Odrv4 I__5359 (
            .O(N__41002),
            .I(\uart_pc.stateZ0Z_1 ));
    CascadeMux I__5358 (
            .O(N__40999),
            .I(\uart_pc.state_srsts_i_0_2_cascade_ ));
    CascadeMux I__5357 (
            .O(N__40996),
            .I(\uart_pc.N_144_1_cascade_ ));
    CascadeMux I__5356 (
            .O(N__40993),
            .I(\Commands_frame_decoder.WDT_RNIHV6PZ0Z_11_cascade_ ));
    InMux I__5355 (
            .O(N__40990),
            .I(N__40987));
    LocalMux I__5354 (
            .O(N__40987),
            .I(\Commands_frame_decoder.WDT_RNIET8A1_0Z0Z_4 ));
    InMux I__5353 (
            .O(N__40984),
            .I(N__40981));
    LocalMux I__5352 (
            .O(N__40981),
            .I(\Commands_frame_decoder.WDT_RNI30853Z0Z_10 ));
    InMux I__5351 (
            .O(N__40978),
            .I(N__40969));
    InMux I__5350 (
            .O(N__40977),
            .I(N__40969));
    InMux I__5349 (
            .O(N__40976),
            .I(N__40969));
    LocalMux I__5348 (
            .O(N__40969),
            .I(\Commands_frame_decoder.preinitZ0 ));
    InMux I__5347 (
            .O(N__40966),
            .I(N__40963));
    LocalMux I__5346 (
            .O(N__40963),
            .I(\Commands_frame_decoder.WDT_RNI2VDI1Z0Z_10 ));
    InMux I__5345 (
            .O(N__40960),
            .I(N__40957));
    LocalMux I__5344 (
            .O(N__40957),
            .I(\Commands_frame_decoder.WDT_RNITK4L_0Z0Z_8 ));
    CascadeMux I__5343 (
            .O(N__40954),
            .I(\Commands_frame_decoder.WDT_RNIET8A1Z0Z_4_cascade_ ));
    InMux I__5342 (
            .O(N__40951),
            .I(N__40948));
    LocalMux I__5341 (
            .O(N__40948),
            .I(\Commands_frame_decoder.WDT_RNIHV6P_0Z0Z_11 ));
    CascadeMux I__5340 (
            .O(N__40945),
            .I(\Commands_frame_decoder.WDT8lt14_0_cascade_ ));
    InMux I__5339 (
            .O(N__40942),
            .I(N__40938));
    InMux I__5338 (
            .O(N__40941),
            .I(N__40935));
    LocalMux I__5337 (
            .O(N__40938),
            .I(N__40930));
    LocalMux I__5336 (
            .O(N__40935),
            .I(N__40930));
    Odrv4 I__5335 (
            .O(N__40930),
            .I(scaler_4_data_9));
    InMux I__5334 (
            .O(N__40927),
            .I(\scaler_4.un2_source_data_0_cry_4 ));
    InMux I__5333 (
            .O(N__40924),
            .I(\scaler_4.un2_source_data_0_cry_5 ));
    CascadeMux I__5332 (
            .O(N__40921),
            .I(N__40917));
    InMux I__5331 (
            .O(N__40920),
            .I(N__40914));
    InMux I__5330 (
            .O(N__40917),
            .I(N__40911));
    LocalMux I__5329 (
            .O(N__40914),
            .I(N__40908));
    LocalMux I__5328 (
            .O(N__40911),
            .I(N__40905));
    Odrv12 I__5327 (
            .O(N__40908),
            .I(scaler_4_data_11));
    Odrv4 I__5326 (
            .O(N__40905),
            .I(scaler_4_data_11));
    InMux I__5325 (
            .O(N__40900),
            .I(\scaler_4.un2_source_data_0_cry_6 ));
    InMux I__5324 (
            .O(N__40897),
            .I(\scaler_4.un2_source_data_0_cry_7 ));
    InMux I__5323 (
            .O(N__40894),
            .I(bfn_7_12_0_));
    InMux I__5322 (
            .O(N__40891),
            .I(\scaler_4.un2_source_data_0_cry_9 ));
    InMux I__5321 (
            .O(N__40888),
            .I(N__40885));
    LocalMux I__5320 (
            .O(N__40885),
            .I(N__40882));
    Odrv4 I__5319 (
            .O(N__40882),
            .I(scaler_4_data_14));
    CascadeMux I__5318 (
            .O(N__40879),
            .I(\Commands_frame_decoder.preinit_RNIHOVZ0Z81_cascade_ ));
    InMux I__5317 (
            .O(N__40876),
            .I(N__40873));
    LocalMux I__5316 (
            .O(N__40873),
            .I(\ppm_encoder_1.un1_rudder_cry_10_THRU_CO ));
    InMux I__5315 (
            .O(N__40870),
            .I(\ppm_encoder_1.un1_rudder_cry_10 ));
    InMux I__5314 (
            .O(N__40867),
            .I(\ppm_encoder_1.un1_rudder_cry_11 ));
    InMux I__5313 (
            .O(N__40864),
            .I(\ppm_encoder_1.un1_rudder_cry_12 ));
    InMux I__5312 (
            .O(N__40861),
            .I(bfn_7_10_0_));
    InMux I__5311 (
            .O(N__40858),
            .I(\scaler_4.un2_source_data_0_cry_1 ));
    InMux I__5310 (
            .O(N__40855),
            .I(N__40851));
    InMux I__5309 (
            .O(N__40854),
            .I(N__40848));
    LocalMux I__5308 (
            .O(N__40851),
            .I(N__40845));
    LocalMux I__5307 (
            .O(N__40848),
            .I(N__40842));
    Odrv4 I__5306 (
            .O(N__40845),
            .I(scaler_4_data_7));
    Odrv4 I__5305 (
            .O(N__40842),
            .I(scaler_4_data_7));
    InMux I__5304 (
            .O(N__40837),
            .I(\scaler_4.un2_source_data_0_cry_2 ));
    InMux I__5303 (
            .O(N__40834),
            .I(\scaler_4.un2_source_data_0_cry_3 ));
    InMux I__5302 (
            .O(N__40831),
            .I(N__40824));
    InMux I__5301 (
            .O(N__40830),
            .I(N__40824));
    InMux I__5300 (
            .O(N__40829),
            .I(N__40821));
    LocalMux I__5299 (
            .O(N__40824),
            .I(N__40818));
    LocalMux I__5298 (
            .O(N__40821),
            .I(\ppm_encoder_1.elevatorZ0Z_11 ));
    Odrv4 I__5297 (
            .O(N__40818),
            .I(\ppm_encoder_1.elevatorZ0Z_11 ));
    InMux I__5296 (
            .O(N__40813),
            .I(N__40810));
    LocalMux I__5295 (
            .O(N__40810),
            .I(N__40805));
    InMux I__5294 (
            .O(N__40809),
            .I(N__40802));
    CascadeMux I__5293 (
            .O(N__40808),
            .I(N__40799));
    Span4Mux_v I__5292 (
            .O(N__40805),
            .I(N__40796));
    LocalMux I__5291 (
            .O(N__40802),
            .I(N__40793));
    InMux I__5290 (
            .O(N__40799),
            .I(N__40790));
    Span4Mux_h I__5289 (
            .O(N__40796),
            .I(N__40787));
    Span4Mux_h I__5288 (
            .O(N__40793),
            .I(N__40784));
    LocalMux I__5287 (
            .O(N__40790),
            .I(\ppm_encoder_1.elevatorZ0Z_2 ));
    Odrv4 I__5286 (
            .O(N__40787),
            .I(\ppm_encoder_1.elevatorZ0Z_2 ));
    Odrv4 I__5285 (
            .O(N__40784),
            .I(\ppm_encoder_1.elevatorZ0Z_2 ));
    CascadeMux I__5284 (
            .O(N__40777),
            .I(N__40772));
    CascadeMux I__5283 (
            .O(N__40776),
            .I(N__40769));
    CascadeMux I__5282 (
            .O(N__40775),
            .I(N__40766));
    InMux I__5281 (
            .O(N__40772),
            .I(N__40763));
    InMux I__5280 (
            .O(N__40769),
            .I(N__40758));
    InMux I__5279 (
            .O(N__40766),
            .I(N__40758));
    LocalMux I__5278 (
            .O(N__40763),
            .I(N__40755));
    LocalMux I__5277 (
            .O(N__40758),
            .I(N__40752));
    Odrv4 I__5276 (
            .O(N__40755),
            .I(\ppm_encoder_1.rudderZ0Z_11 ));
    Odrv4 I__5275 (
            .O(N__40752),
            .I(\ppm_encoder_1.rudderZ0Z_11 ));
    InMux I__5274 (
            .O(N__40747),
            .I(N__40744));
    LocalMux I__5273 (
            .O(N__40744),
            .I(\ppm_encoder_1.un1_rudder_cry_6_THRU_CO ));
    InMux I__5272 (
            .O(N__40741),
            .I(\ppm_encoder_1.un1_rudder_cry_6 ));
    InMux I__5271 (
            .O(N__40738),
            .I(\ppm_encoder_1.un1_rudder_cry_7 ));
    InMux I__5270 (
            .O(N__40735),
            .I(N__40732));
    LocalMux I__5269 (
            .O(N__40732),
            .I(\ppm_encoder_1.un1_rudder_cry_8_THRU_CO ));
    InMux I__5268 (
            .O(N__40729),
            .I(\ppm_encoder_1.un1_rudder_cry_8 ));
    InMux I__5267 (
            .O(N__40726),
            .I(\ppm_encoder_1.un1_rudder_cry_9 ));
    InMux I__5266 (
            .O(N__40723),
            .I(N__40720));
    LocalMux I__5265 (
            .O(N__40720),
            .I(N__40717));
    Odrv4 I__5264 (
            .O(N__40717),
            .I(\ppm_encoder_1.un2_throttle_iv_0_0_4 ));
    CascadeMux I__5263 (
            .O(N__40714),
            .I(\ppm_encoder_1.un2_throttle_iv_0_2_10_cascade_ ));
    CascadeMux I__5262 (
            .O(N__40711),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_10_cascade_ ));
    InMux I__5261 (
            .O(N__40708),
            .I(N__40705));
    LocalMux I__5260 (
            .O(N__40705),
            .I(\ppm_encoder_1.N_458 ));
    InMux I__5259 (
            .O(N__40702),
            .I(N__40699));
    LocalMux I__5258 (
            .O(N__40699),
            .I(\ppm_encoder_1.un2_throttle_iv_0_1_10 ));
    InMux I__5257 (
            .O(N__40696),
            .I(N__40693));
    LocalMux I__5256 (
            .O(N__40693),
            .I(N__40689));
    InMux I__5255 (
            .O(N__40692),
            .I(N__40686));
    Span4Mux_h I__5254 (
            .O(N__40689),
            .I(N__40682));
    LocalMux I__5253 (
            .O(N__40686),
            .I(N__40679));
    InMux I__5252 (
            .O(N__40685),
            .I(N__40676));
    Span4Mux_v I__5251 (
            .O(N__40682),
            .I(N__40673));
    Span4Mux_h I__5250 (
            .O(N__40679),
            .I(N__40670));
    LocalMux I__5249 (
            .O(N__40676),
            .I(\ppm_encoder_1.elevatorZ0Z_1 ));
    Odrv4 I__5248 (
            .O(N__40673),
            .I(\ppm_encoder_1.elevatorZ0Z_1 ));
    Odrv4 I__5247 (
            .O(N__40670),
            .I(\ppm_encoder_1.elevatorZ0Z_1 ));
    InMux I__5246 (
            .O(N__40663),
            .I(N__40660));
    LocalMux I__5245 (
            .O(N__40660),
            .I(N__40657));
    Span4Mux_v I__5244 (
            .O(N__40657),
            .I(N__40654));
    Odrv4 I__5243 (
            .O(N__40654),
            .I(\uart_drone_sync.aux_0__0__0_0 ));
    CascadeMux I__5242 (
            .O(N__40651),
            .I(N__40646));
    CascadeMux I__5241 (
            .O(N__40650),
            .I(N__40643));
    InMux I__5240 (
            .O(N__40649),
            .I(N__40640));
    InMux I__5239 (
            .O(N__40646),
            .I(N__40637));
    InMux I__5238 (
            .O(N__40643),
            .I(N__40634));
    LocalMux I__5237 (
            .O(N__40640),
            .I(N__40631));
    LocalMux I__5236 (
            .O(N__40637),
            .I(N__40628));
    LocalMux I__5235 (
            .O(N__40634),
            .I(N__40623));
    Span4Mux_v I__5234 (
            .O(N__40631),
            .I(N__40623));
    Span4Mux_h I__5233 (
            .O(N__40628),
            .I(N__40620));
    Odrv4 I__5232 (
            .O(N__40623),
            .I(\ppm_encoder_1.throttleZ0Z_11 ));
    Odrv4 I__5231 (
            .O(N__40620),
            .I(\ppm_encoder_1.throttleZ0Z_11 ));
    InMux I__5230 (
            .O(N__40615),
            .I(N__40612));
    LocalMux I__5229 (
            .O(N__40612),
            .I(\ppm_encoder_1.un2_throttle_iv_0_1_11 ));
    CascadeMux I__5228 (
            .O(N__40609),
            .I(\ppm_encoder_1.un2_throttle_iv_0_0_11_cascade_ ));
    CascadeMux I__5227 (
            .O(N__40606),
            .I(\ppm_encoder_1.un2_throttle_iv_0_0_13_cascade_ ));
    InMux I__5226 (
            .O(N__40603),
            .I(N__40600));
    LocalMux I__5225 (
            .O(N__40600),
            .I(\ppm_encoder_1.N_516 ));
    InMux I__5224 (
            .O(N__40597),
            .I(N__40594));
    LocalMux I__5223 (
            .O(N__40594),
            .I(N__40591));
    Span4Mux_h I__5222 (
            .O(N__40591),
            .I(N__40588));
    Span4Mux_h I__5221 (
            .O(N__40588),
            .I(N__40585));
    Odrv4 I__5220 (
            .O(N__40585),
            .I(\ppm_encoder_1.N_440 ));
    CascadeMux I__5219 (
            .O(N__40582),
            .I(\ppm_encoder_1.N_516_cascade_ ));
    InMux I__5218 (
            .O(N__40579),
            .I(N__40576));
    LocalMux I__5217 (
            .O(N__40576),
            .I(uart_input_drone_c));
    InMux I__5216 (
            .O(N__40573),
            .I(N__40570));
    LocalMux I__5215 (
            .O(N__40570),
            .I(N__40567));
    Odrv4 I__5214 (
            .O(N__40567),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_13 ));
    InMux I__5213 (
            .O(N__40564),
            .I(N__40558));
    InMux I__5212 (
            .O(N__40563),
            .I(N__40558));
    LocalMux I__5211 (
            .O(N__40558),
            .I(N__40554));
    InMux I__5210 (
            .O(N__40557),
            .I(N__40551));
    Span4Mux_v I__5209 (
            .O(N__40554),
            .I(N__40546));
    LocalMux I__5208 (
            .O(N__40551),
            .I(N__40546));
    Span4Mux_h I__5207 (
            .O(N__40546),
            .I(N__40543));
    Span4Mux_v I__5206 (
            .O(N__40543),
            .I(N__40540));
    Span4Mux_v I__5205 (
            .O(N__40540),
            .I(N__40537));
    Odrv4 I__5204 (
            .O(N__40537),
            .I(\pid_alt.error_d_regZ0Z_15 ));
    InMux I__5203 (
            .O(N__40534),
            .I(N__40531));
    LocalMux I__5202 (
            .O(N__40531),
            .I(N__40527));
    InMux I__5201 (
            .O(N__40530),
            .I(N__40524));
    Span4Mux_h I__5200 (
            .O(N__40527),
            .I(N__40521));
    LocalMux I__5199 (
            .O(N__40524),
            .I(\pid_alt.error_d_reg_prevZ0Z_15 ));
    Odrv4 I__5198 (
            .O(N__40521),
            .I(\pid_alt.error_d_reg_prevZ0Z_15 ));
    CEMux I__5197 (
            .O(N__40516),
            .I(N__40450));
    CEMux I__5196 (
            .O(N__40515),
            .I(N__40450));
    CEMux I__5195 (
            .O(N__40514),
            .I(N__40450));
    CEMux I__5194 (
            .O(N__40513),
            .I(N__40450));
    CEMux I__5193 (
            .O(N__40512),
            .I(N__40450));
    CEMux I__5192 (
            .O(N__40511),
            .I(N__40450));
    CEMux I__5191 (
            .O(N__40510),
            .I(N__40450));
    CEMux I__5190 (
            .O(N__40509),
            .I(N__40450));
    CEMux I__5189 (
            .O(N__40508),
            .I(N__40450));
    CEMux I__5188 (
            .O(N__40507),
            .I(N__40450));
    CEMux I__5187 (
            .O(N__40506),
            .I(N__40450));
    CEMux I__5186 (
            .O(N__40505),
            .I(N__40450));
    CEMux I__5185 (
            .O(N__40504),
            .I(N__40450));
    CEMux I__5184 (
            .O(N__40503),
            .I(N__40450));
    CEMux I__5183 (
            .O(N__40502),
            .I(N__40450));
    CEMux I__5182 (
            .O(N__40501),
            .I(N__40450));
    CEMux I__5181 (
            .O(N__40500),
            .I(N__40450));
    CEMux I__5180 (
            .O(N__40499),
            .I(N__40450));
    CEMux I__5179 (
            .O(N__40498),
            .I(N__40450));
    CEMux I__5178 (
            .O(N__40497),
            .I(N__40450));
    CEMux I__5177 (
            .O(N__40496),
            .I(N__40450));
    CEMux I__5176 (
            .O(N__40495),
            .I(N__40450));
    GlobalMux I__5175 (
            .O(N__40450),
            .I(N__40447));
    gio2CtrlBuf I__5174 (
            .O(N__40447),
            .I(\pid_alt.state_0_g_0 ));
    InMux I__5173 (
            .O(N__40444),
            .I(N__40441));
    LocalMux I__5172 (
            .O(N__40441),
            .I(N__40438));
    Odrv4 I__5171 (
            .O(N__40438),
            .I(\pid_alt.N_111 ));
    CascadeMux I__5170 (
            .O(N__40435),
            .I(\pid_alt.un1_reset_1_0_i_cascade_ ));
    CascadeMux I__5169 (
            .O(N__40432),
            .I(N__40429));
    InMux I__5168 (
            .O(N__40429),
            .I(N__40426));
    LocalMux I__5167 (
            .O(N__40426),
            .I(N__40423));
    Odrv4 I__5166 (
            .O(N__40423),
            .I(alt_command_7));
    CascadeMux I__5165 (
            .O(N__40420),
            .I(N__40417));
    InMux I__5164 (
            .O(N__40417),
            .I(N__40412));
    CascadeMux I__5163 (
            .O(N__40416),
            .I(N__40408));
    InMux I__5162 (
            .O(N__40415),
            .I(N__40405));
    LocalMux I__5161 (
            .O(N__40412),
            .I(N__40402));
    InMux I__5160 (
            .O(N__40411),
            .I(N__40399));
    InMux I__5159 (
            .O(N__40408),
            .I(N__40396));
    LocalMux I__5158 (
            .O(N__40405),
            .I(N__40391));
    Span4Mux_s1_v I__5157 (
            .O(N__40402),
            .I(N__40391));
    LocalMux I__5156 (
            .O(N__40399),
            .I(N__40386));
    LocalMux I__5155 (
            .O(N__40396),
            .I(N__40386));
    Odrv4 I__5154 (
            .O(N__40391),
            .I(\ppm_encoder_1.init_pulsesZ0Z_1 ));
    Odrv12 I__5153 (
            .O(N__40386),
            .I(\ppm_encoder_1.init_pulsesZ0Z_1 ));
    CascadeMux I__5152 (
            .O(N__40381),
            .I(N__40377));
    CascadeMux I__5151 (
            .O(N__40380),
            .I(N__40374));
    InMux I__5150 (
            .O(N__40377),
            .I(N__40366));
    InMux I__5149 (
            .O(N__40374),
            .I(N__40366));
    InMux I__5148 (
            .O(N__40373),
            .I(N__40366));
    LocalMux I__5147 (
            .O(N__40366),
            .I(\Commands_frame_decoder.source_CH1data8 ));
    InMux I__5146 (
            .O(N__40363),
            .I(N__40359));
    InMux I__5145 (
            .O(N__40362),
            .I(N__40356));
    LocalMux I__5144 (
            .O(N__40359),
            .I(N__40353));
    LocalMux I__5143 (
            .O(N__40356),
            .I(alt_command_2));
    Odrv4 I__5142 (
            .O(N__40353),
            .I(alt_command_2));
    CascadeMux I__5141 (
            .O(N__40348),
            .I(\Commands_frame_decoder.state_ns_i_a2_0_2_0_cascade_ ));
    CascadeMux I__5140 (
            .O(N__40345),
            .I(N__40342));
    InMux I__5139 (
            .O(N__40342),
            .I(N__40339));
    LocalMux I__5138 (
            .O(N__40339),
            .I(alt_command_4));
    CascadeMux I__5137 (
            .O(N__40336),
            .I(N__40333));
    InMux I__5136 (
            .O(N__40333),
            .I(N__40330));
    LocalMux I__5135 (
            .O(N__40330),
            .I(alt_command_5));
    CascadeMux I__5134 (
            .O(N__40327),
            .I(N__40324));
    InMux I__5133 (
            .O(N__40324),
            .I(N__40321));
    LocalMux I__5132 (
            .O(N__40321),
            .I(alt_command_6));
    InMux I__5131 (
            .O(N__40318),
            .I(N__40315));
    LocalMux I__5130 (
            .O(N__40315),
            .I(N__40312));
    Span4Mux_v I__5129 (
            .O(N__40312),
            .I(N__40309));
    Span4Mux_h I__5128 (
            .O(N__40309),
            .I(N__40306));
    Odrv4 I__5127 (
            .O(N__40306),
            .I(alt_kp_2));
    InMux I__5126 (
            .O(N__40303),
            .I(N__40300));
    LocalMux I__5125 (
            .O(N__40300),
            .I(drone_altitude_i_8));
    InMux I__5124 (
            .O(N__40297),
            .I(N__40293));
    InMux I__5123 (
            .O(N__40296),
            .I(N__40290));
    LocalMux I__5122 (
            .O(N__40293),
            .I(N__40287));
    LocalMux I__5121 (
            .O(N__40290),
            .I(N__40284));
    Span4Mux_v I__5120 (
            .O(N__40287),
            .I(N__40281));
    Span4Mux_v I__5119 (
            .O(N__40284),
            .I(N__40278));
    Span4Mux_v I__5118 (
            .O(N__40281),
            .I(N__40275));
    Span4Mux_h I__5117 (
            .O(N__40278),
            .I(N__40272));
    Odrv4 I__5116 (
            .O(N__40275),
            .I(\pid_alt.error_p_regZ0Z_15 ));
    Odrv4 I__5115 (
            .O(N__40272),
            .I(\pid_alt.error_p_regZ0Z_15 ));
    InMux I__5114 (
            .O(N__40267),
            .I(N__40264));
    LocalMux I__5113 (
            .O(N__40264),
            .I(N__40260));
    InMux I__5112 (
            .O(N__40263),
            .I(N__40257));
    Span4Mux_v I__5111 (
            .O(N__40260),
            .I(N__40252));
    LocalMux I__5110 (
            .O(N__40257),
            .I(N__40252));
    Span4Mux_h I__5109 (
            .O(N__40252),
            .I(N__40249));
    Odrv4 I__5108 (
            .O(N__40249),
            .I(\pid_alt.error_d_reg_prev_esr_RNISPHMZ0Z_15 ));
    InMux I__5107 (
            .O(N__40246),
            .I(N__40243));
    LocalMux I__5106 (
            .O(N__40243),
            .I(N__40240));
    Span4Mux_h I__5105 (
            .O(N__40240),
            .I(N__40237));
    Span4Mux_v I__5104 (
            .O(N__40237),
            .I(N__40234));
    Span4Mux_v I__5103 (
            .O(N__40234),
            .I(N__40231));
    Span4Mux_v I__5102 (
            .O(N__40231),
            .I(N__40228));
    Odrv4 I__5101 (
            .O(N__40228),
            .I(uart_input_pc_c));
    InMux I__5100 (
            .O(N__40225),
            .I(N__40222));
    LocalMux I__5099 (
            .O(N__40222),
            .I(\uart_pc_sync.aux_0__0_Z0Z_0 ));
    InMux I__5098 (
            .O(N__40219),
            .I(N__40213));
    InMux I__5097 (
            .O(N__40218),
            .I(N__40208));
    InMux I__5096 (
            .O(N__40217),
            .I(N__40208));
    InMux I__5095 (
            .O(N__40216),
            .I(N__40205));
    LocalMux I__5094 (
            .O(N__40213),
            .I(N__40200));
    LocalMux I__5093 (
            .O(N__40208),
            .I(N__40200));
    LocalMux I__5092 (
            .O(N__40205),
            .I(N__40197));
    Odrv4 I__5091 (
            .O(N__40200),
            .I(\pid_alt.pid_preregZ0Z_12 ));
    Odrv4 I__5090 (
            .O(N__40197),
            .I(\pid_alt.pid_preregZ0Z_12 ));
    InMux I__5089 (
            .O(N__40192),
            .I(N__40188));
    CascadeMux I__5088 (
            .O(N__40191),
            .I(N__40185));
    LocalMux I__5087 (
            .O(N__40188),
            .I(N__40182));
    InMux I__5086 (
            .O(N__40185),
            .I(N__40179));
    Span4Mux_v I__5085 (
            .O(N__40182),
            .I(N__40176));
    LocalMux I__5084 (
            .O(N__40179),
            .I(\pid_alt.pid_preregZ0Z_5 ));
    Odrv4 I__5083 (
            .O(N__40176),
            .I(\pid_alt.pid_preregZ0Z_5 ));
    InMux I__5082 (
            .O(N__40171),
            .I(N__40167));
    InMux I__5081 (
            .O(N__40170),
            .I(N__40164));
    LocalMux I__5080 (
            .O(N__40167),
            .I(N__40157));
    LocalMux I__5079 (
            .O(N__40164),
            .I(N__40157));
    InMux I__5078 (
            .O(N__40163),
            .I(N__40152));
    InMux I__5077 (
            .O(N__40162),
            .I(N__40152));
    Sp12to4 I__5076 (
            .O(N__40157),
            .I(N__40147));
    LocalMux I__5075 (
            .O(N__40152),
            .I(N__40147));
    Odrv12 I__5074 (
            .O(N__40147),
            .I(\pid_alt.N_154 ));
    CEMux I__5073 (
            .O(N__40144),
            .I(N__40141));
    LocalMux I__5072 (
            .O(N__40141),
            .I(N__40138));
    Span12Mux_s10_v I__5071 (
            .O(N__40138),
            .I(N__40135));
    Odrv12 I__5070 (
            .O(N__40135),
            .I(\pid_alt.state_1_0_0 ));
    CascadeMux I__5069 (
            .O(N__40132),
            .I(\Commands_frame_decoder.source_CH1data8_cascade_ ));
    CascadeMux I__5068 (
            .O(N__40129),
            .I(N__40125));
    InMux I__5067 (
            .O(N__40128),
            .I(N__40122));
    InMux I__5066 (
            .O(N__40125),
            .I(N__40119));
    LocalMux I__5065 (
            .O(N__40122),
            .I(alt_command_1));
    LocalMux I__5064 (
            .O(N__40119),
            .I(alt_command_1));
    CascadeMux I__5063 (
            .O(N__40114),
            .I(N__40111));
    InMux I__5062 (
            .O(N__40111),
            .I(N__40108));
    LocalMux I__5061 (
            .O(N__40108),
            .I(\Commands_frame_decoder.source_CH1data8lto7Z0Z_2 ));
    InMux I__5060 (
            .O(N__40105),
            .I(N__40101));
    InMux I__5059 (
            .O(N__40104),
            .I(N__40098));
    LocalMux I__5058 (
            .O(N__40101),
            .I(alt_command_3));
    LocalMux I__5057 (
            .O(N__40098),
            .I(alt_command_3));
    CascadeMux I__5056 (
            .O(N__40093),
            .I(N__40089));
    InMux I__5055 (
            .O(N__40092),
            .I(N__40086));
    InMux I__5054 (
            .O(N__40089),
            .I(N__40083));
    LocalMux I__5053 (
            .O(N__40086),
            .I(alt_command_0));
    LocalMux I__5052 (
            .O(N__40083),
            .I(alt_command_0));
    CascadeMux I__5051 (
            .O(N__40078),
            .I(N__40074));
    CascadeMux I__5050 (
            .O(N__40077),
            .I(N__40071));
    InMux I__5049 (
            .O(N__40074),
            .I(N__40068));
    InMux I__5048 (
            .O(N__40071),
            .I(N__40065));
    LocalMux I__5047 (
            .O(N__40068),
            .I(N__40062));
    LocalMux I__5046 (
            .O(N__40065),
            .I(\pid_alt.error_d_reg_prev_esr_RNIUI2T2Z0Z_6 ));
    Odrv4 I__5045 (
            .O(N__40062),
            .I(\pid_alt.error_d_reg_prev_esr_RNIUI2T2Z0Z_6 ));
    InMux I__5044 (
            .O(N__40057),
            .I(N__40048));
    InMux I__5043 (
            .O(N__40056),
            .I(N__40048));
    InMux I__5042 (
            .O(N__40055),
            .I(N__40048));
    LocalMux I__5041 (
            .O(N__40048),
            .I(N__40045));
    Span4Mux_h I__5040 (
            .O(N__40045),
            .I(N__40042));
    Span4Mux_v I__5039 (
            .O(N__40042),
            .I(N__40039));
    Span4Mux_v I__5038 (
            .O(N__40039),
            .I(N__40036));
    Odrv4 I__5037 (
            .O(N__40036),
            .I(\pid_alt.error_d_regZ0Z_7 ));
    CascadeMux I__5036 (
            .O(N__40033),
            .I(N__40030));
    InMux I__5035 (
            .O(N__40030),
            .I(N__40024));
    InMux I__5034 (
            .O(N__40029),
            .I(N__40024));
    LocalMux I__5033 (
            .O(N__40024),
            .I(\pid_alt.error_d_reg_prevZ0Z_7 ));
    InMux I__5032 (
            .O(N__40021),
            .I(N__40015));
    InMux I__5031 (
            .O(N__40020),
            .I(N__40015));
    LocalMux I__5030 (
            .O(N__40015),
            .I(N__40012));
    Span4Mux_h I__5029 (
            .O(N__40012),
            .I(N__40009));
    Span4Mux_v I__5028 (
            .O(N__40009),
            .I(N__40006));
    Span4Mux_h I__5027 (
            .O(N__40006),
            .I(N__40003));
    Odrv4 I__5026 (
            .O(N__40003),
            .I(\pid_alt.error_p_regZ0Z_7 ));
    InMux I__5025 (
            .O(N__40000),
            .I(N__39997));
    LocalMux I__5024 (
            .O(N__39997),
            .I(\pid_alt.error_d_reg_prev_esr_RNIF2611_0Z0Z_7 ));
    InMux I__5023 (
            .O(N__39994),
            .I(N__39990));
    CascadeMux I__5022 (
            .O(N__39993),
            .I(N__39987));
    LocalMux I__5021 (
            .O(N__39990),
            .I(N__39984));
    InMux I__5020 (
            .O(N__39987),
            .I(N__39981));
    Odrv4 I__5019 (
            .O(N__39984),
            .I(\pid_alt.error_d_reg_prev_esr_RNIL81T2Z0Z_5 ));
    LocalMux I__5018 (
            .O(N__39981),
            .I(\pid_alt.error_d_reg_prev_esr_RNIL81T2Z0Z_5 ));
    InMux I__5017 (
            .O(N__39976),
            .I(N__39970));
    InMux I__5016 (
            .O(N__39975),
            .I(N__39970));
    LocalMux I__5015 (
            .O(N__39970),
            .I(N__39967));
    Odrv12 I__5014 (
            .O(N__39967),
            .I(\pid_alt.error_d_reg_prev_esr_RNICV511Z0Z_6 ));
    CascadeMux I__5013 (
            .O(N__39964),
            .I(\pid_alt.error_d_reg_prev_esr_RNIF2611_0Z0Z_7_cascade_ ));
    InMux I__5012 (
            .O(N__39961),
            .I(N__39958));
    LocalMux I__5011 (
            .O(N__39958),
            .I(N__39953));
    InMux I__5010 (
            .O(N__39957),
            .I(N__39948));
    InMux I__5009 (
            .O(N__39956),
            .I(N__39948));
    Span4Mux_h I__5008 (
            .O(N__39953),
            .I(N__39945));
    LocalMux I__5007 (
            .O(N__39948),
            .I(N__39942));
    Span4Mux_v I__5006 (
            .O(N__39945),
            .I(N__39939));
    Span4Mux_h I__5005 (
            .O(N__39942),
            .I(N__39936));
    Odrv4 I__5004 (
            .O(N__39939),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ ));
    Odrv4 I__5003 (
            .O(N__39936),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ ));
    InMux I__5002 (
            .O(N__39931),
            .I(N__39928));
    LocalMux I__5001 (
            .O(N__39928),
            .I(N__39925));
    Odrv4 I__5000 (
            .O(N__39925),
            .I(\pid_alt.error_d_reg_prev_esr_RNIJR3Q5Z0Z_6 ));
    InMux I__4999 (
            .O(N__39922),
            .I(N__39919));
    LocalMux I__4998 (
            .O(N__39919),
            .I(N__39916));
    Span4Mux_h I__4997 (
            .O(N__39916),
            .I(N__39913));
    Span4Mux_h I__4996 (
            .O(N__39913),
            .I(N__39910));
    Odrv4 I__4995 (
            .O(N__39910),
            .I(\pid_front.O_0_21 ));
    InMux I__4994 (
            .O(N__39907),
            .I(N__39904));
    LocalMux I__4993 (
            .O(N__39904),
            .I(N__39901));
    Odrv12 I__4992 (
            .O(N__39901),
            .I(\pid_front.O_0_7 ));
    InMux I__4991 (
            .O(N__39898),
            .I(N__39895));
    LocalMux I__4990 (
            .O(N__39895),
            .I(N__39892));
    Span12Mux_v I__4989 (
            .O(N__39892),
            .I(N__39889));
    Odrv12 I__4988 (
            .O(N__39889),
            .I(\pid_front.O_0_11 ));
    InMux I__4987 (
            .O(N__39886),
            .I(N__39883));
    LocalMux I__4986 (
            .O(N__39883),
            .I(N__39880));
    Span4Mux_h I__4985 (
            .O(N__39880),
            .I(N__39877));
    Span4Mux_h I__4984 (
            .O(N__39877),
            .I(N__39874));
    Odrv4 I__4983 (
            .O(N__39874),
            .I(\pid_front.O_0_12 ));
    InMux I__4982 (
            .O(N__39871),
            .I(N__39862));
    InMux I__4981 (
            .O(N__39870),
            .I(N__39862));
    InMux I__4980 (
            .O(N__39869),
            .I(N__39859));
    InMux I__4979 (
            .O(N__39868),
            .I(N__39854));
    InMux I__4978 (
            .O(N__39867),
            .I(N__39854));
    LocalMux I__4977 (
            .O(N__39862),
            .I(\pid_alt.pid_preregZ0Z_4 ));
    LocalMux I__4976 (
            .O(N__39859),
            .I(\pid_alt.pid_preregZ0Z_4 ));
    LocalMux I__4975 (
            .O(N__39854),
            .I(\pid_alt.pid_preregZ0Z_4 ));
    CascadeMux I__4974 (
            .O(N__39847),
            .I(\pid_alt.source_pid_9_0_0_4_cascade_ ));
    InMux I__4973 (
            .O(N__39844),
            .I(N__39840));
    InMux I__4972 (
            .O(N__39843),
            .I(N__39837));
    LocalMux I__4971 (
            .O(N__39840),
            .I(N__39834));
    LocalMux I__4970 (
            .O(N__39837),
            .I(N__39831));
    Span4Mux_v I__4969 (
            .O(N__39834),
            .I(N__39826));
    Span4Mux_h I__4968 (
            .O(N__39831),
            .I(N__39826));
    Odrv4 I__4967 (
            .O(N__39826),
            .I(throttle_order_4));
    InMux I__4966 (
            .O(N__39823),
            .I(N__39817));
    InMux I__4965 (
            .O(N__39822),
            .I(N__39817));
    LocalMux I__4964 (
            .O(N__39817),
            .I(N__39814));
    Span4Mux_h I__4963 (
            .O(N__39814),
            .I(N__39811));
    Odrv4 I__4962 (
            .O(N__39811),
            .I(\pid_alt.N_52 ));
    InMux I__4961 (
            .O(N__39808),
            .I(N__39805));
    LocalMux I__4960 (
            .O(N__39805),
            .I(N__39801));
    InMux I__4959 (
            .O(N__39804),
            .I(N__39798));
    Span4Mux_h I__4958 (
            .O(N__39801),
            .I(N__39793));
    LocalMux I__4957 (
            .O(N__39798),
            .I(N__39793));
    Span4Mux_v I__4956 (
            .O(N__39793),
            .I(N__39790));
    Odrv4 I__4955 (
            .O(N__39790),
            .I(throttle_order_5));
    CascadeMux I__4954 (
            .O(N__39787),
            .I(N__39782));
    CascadeMux I__4953 (
            .O(N__39786),
            .I(N__39777));
    CascadeMux I__4952 (
            .O(N__39785),
            .I(N__39773));
    InMux I__4951 (
            .O(N__39782),
            .I(N__39769));
    InMux I__4950 (
            .O(N__39781),
            .I(N__39755));
    InMux I__4949 (
            .O(N__39780),
            .I(N__39755));
    InMux I__4948 (
            .O(N__39777),
            .I(N__39755));
    InMux I__4947 (
            .O(N__39776),
            .I(N__39755));
    InMux I__4946 (
            .O(N__39773),
            .I(N__39755));
    InMux I__4945 (
            .O(N__39772),
            .I(N__39752));
    LocalMux I__4944 (
            .O(N__39769),
            .I(N__39749));
    InMux I__4943 (
            .O(N__39768),
            .I(N__39742));
    InMux I__4942 (
            .O(N__39767),
            .I(N__39742));
    InMux I__4941 (
            .O(N__39766),
            .I(N__39742));
    LocalMux I__4940 (
            .O(N__39755),
            .I(N__39739));
    LocalMux I__4939 (
            .O(N__39752),
            .I(N__39736));
    Span4Mux_v I__4938 (
            .O(N__39749),
            .I(N__39727));
    LocalMux I__4937 (
            .O(N__39742),
            .I(N__39727));
    Span4Mux_h I__4936 (
            .O(N__39739),
            .I(N__39727));
    Span4Mux_h I__4935 (
            .O(N__39736),
            .I(N__39727));
    Odrv4 I__4934 (
            .O(N__39727),
            .I(\pid_alt.pid_preregZ0Z_24 ));
    CascadeMux I__4933 (
            .O(N__39724),
            .I(N__39719));
    InMux I__4932 (
            .O(N__39723),
            .I(N__39716));
    InMux I__4931 (
            .O(N__39722),
            .I(N__39711));
    InMux I__4930 (
            .O(N__39719),
            .I(N__39708));
    LocalMux I__4929 (
            .O(N__39716),
            .I(N__39704));
    InMux I__4928 (
            .O(N__39715),
            .I(N__39699));
    InMux I__4927 (
            .O(N__39714),
            .I(N__39699));
    LocalMux I__4926 (
            .O(N__39711),
            .I(N__39694));
    LocalMux I__4925 (
            .O(N__39708),
            .I(N__39694));
    InMux I__4924 (
            .O(N__39707),
            .I(N__39691));
    Span4Mux_h I__4923 (
            .O(N__39704),
            .I(N__39686));
    LocalMux I__4922 (
            .O(N__39699),
            .I(N__39686));
    Span4Mux_h I__4921 (
            .O(N__39694),
            .I(N__39683));
    LocalMux I__4920 (
            .O(N__39691),
            .I(\pid_alt.pid_preregZ0Z_13 ));
    Odrv4 I__4919 (
            .O(N__39686),
            .I(\pid_alt.pid_preregZ0Z_13 ));
    Odrv4 I__4918 (
            .O(N__39683),
            .I(\pid_alt.pid_preregZ0Z_13 ));
    InMux I__4917 (
            .O(N__39676),
            .I(N__39670));
    InMux I__4916 (
            .O(N__39675),
            .I(N__39656));
    InMux I__4915 (
            .O(N__39674),
            .I(N__39656));
    InMux I__4914 (
            .O(N__39673),
            .I(N__39656));
    LocalMux I__4913 (
            .O(N__39670),
            .I(N__39653));
    InMux I__4912 (
            .O(N__39669),
            .I(N__39642));
    InMux I__4911 (
            .O(N__39668),
            .I(N__39642));
    InMux I__4910 (
            .O(N__39667),
            .I(N__39642));
    InMux I__4909 (
            .O(N__39666),
            .I(N__39642));
    InMux I__4908 (
            .O(N__39665),
            .I(N__39642));
    InMux I__4907 (
            .O(N__39664),
            .I(N__39637));
    InMux I__4906 (
            .O(N__39663),
            .I(N__39637));
    LocalMux I__4905 (
            .O(N__39656),
            .I(\pid_alt.N_539 ));
    Odrv4 I__4904 (
            .O(N__39653),
            .I(\pid_alt.N_539 ));
    LocalMux I__4903 (
            .O(N__39642),
            .I(\pid_alt.N_539 ));
    LocalMux I__4902 (
            .O(N__39637),
            .I(\pid_alt.N_539 ));
    InMux I__4901 (
            .O(N__39628),
            .I(N__39624));
    InMux I__4900 (
            .O(N__39627),
            .I(N__39621));
    LocalMux I__4899 (
            .O(N__39624),
            .I(N__39618));
    LocalMux I__4898 (
            .O(N__39621),
            .I(N__39615));
    Sp12to4 I__4897 (
            .O(N__39618),
            .I(N__39612));
    Span4Mux_h I__4896 (
            .O(N__39615),
            .I(N__39609));
    Odrv12 I__4895 (
            .O(N__39612),
            .I(throttle_order_13));
    Odrv4 I__4894 (
            .O(N__39609),
            .I(throttle_order_13));
    CEMux I__4893 (
            .O(N__39604),
            .I(N__39601));
    LocalMux I__4892 (
            .O(N__39601),
            .I(N__39598));
    Span4Mux_v I__4891 (
            .O(N__39598),
            .I(N__39595));
    Span4Mux_h I__4890 (
            .O(N__39595),
            .I(N__39590));
    CEMux I__4889 (
            .O(N__39594),
            .I(N__39587));
    CEMux I__4888 (
            .O(N__39593),
            .I(N__39584));
    Span4Mux_s2_h I__4887 (
            .O(N__39590),
            .I(N__39579));
    LocalMux I__4886 (
            .O(N__39587),
            .I(N__39579));
    LocalMux I__4885 (
            .O(N__39584),
            .I(N__39576));
    Span4Mux_h I__4884 (
            .O(N__39579),
            .I(N__39573));
    Odrv12 I__4883 (
            .O(N__39576),
            .I(\pid_alt.N_72_i_1 ));
    Odrv4 I__4882 (
            .O(N__39573),
            .I(\pid_alt.N_72_i_1 ));
    SRMux I__4881 (
            .O(N__39568),
            .I(N__39563));
    SRMux I__4880 (
            .O(N__39567),
            .I(N__39560));
    SRMux I__4879 (
            .O(N__39566),
            .I(N__39557));
    LocalMux I__4878 (
            .O(N__39563),
            .I(N__39553));
    LocalMux I__4877 (
            .O(N__39560),
            .I(N__39550));
    LocalMux I__4876 (
            .O(N__39557),
            .I(N__39547));
    SRMux I__4875 (
            .O(N__39556),
            .I(N__39544));
    Span4Mux_h I__4874 (
            .O(N__39553),
            .I(N__39541));
    Span4Mux_v I__4873 (
            .O(N__39550),
            .I(N__39538));
    Span4Mux_h I__4872 (
            .O(N__39547),
            .I(N__39535));
    LocalMux I__4871 (
            .O(N__39544),
            .I(N__39532));
    Odrv4 I__4870 (
            .O(N__39541),
            .I(\pid_alt.un1_reset_0_i ));
    Odrv4 I__4869 (
            .O(N__39538),
            .I(\pid_alt.un1_reset_0_i ));
    Odrv4 I__4868 (
            .O(N__39535),
            .I(\pid_alt.un1_reset_0_i ));
    Odrv12 I__4867 (
            .O(N__39532),
            .I(\pid_alt.un1_reset_0_i ));
    InMux I__4866 (
            .O(N__39523),
            .I(N__39520));
    LocalMux I__4865 (
            .O(N__39520),
            .I(\pid_alt.error_d_reg_prev_esr_RNI5G6Q5Z0Z_7 ));
    InMux I__4864 (
            .O(N__39517),
            .I(N__39513));
    InMux I__4863 (
            .O(N__39516),
            .I(N__39510));
    LocalMux I__4862 (
            .O(N__39513),
            .I(N__39507));
    LocalMux I__4861 (
            .O(N__39510),
            .I(N__39504));
    Span4Mux_v I__4860 (
            .O(N__39507),
            .I(N__39501));
    Span4Mux_h I__4859 (
            .O(N__39504),
            .I(N__39498));
    Span4Mux_v I__4858 (
            .O(N__39501),
            .I(N__39495));
    Span4Mux_v I__4857 (
            .O(N__39498),
            .I(N__39490));
    Span4Mux_h I__4856 (
            .O(N__39495),
            .I(N__39490));
    Odrv4 I__4855 (
            .O(N__39490),
            .I(\pid_alt.error_p_regZ0Z_8 ));
    InMux I__4854 (
            .O(N__39487),
            .I(N__39483));
    InMux I__4853 (
            .O(N__39486),
            .I(N__39480));
    LocalMux I__4852 (
            .O(N__39483),
            .I(N__39477));
    LocalMux I__4851 (
            .O(N__39480),
            .I(\pid_alt.error_d_reg_prevZ0Z_8 ));
    Odrv4 I__4850 (
            .O(N__39477),
            .I(\pid_alt.error_d_reg_prevZ0Z_8 ));
    InMux I__4849 (
            .O(N__39472),
            .I(N__39466));
    InMux I__4848 (
            .O(N__39471),
            .I(N__39466));
    LocalMux I__4847 (
            .O(N__39466),
            .I(N__39462));
    InMux I__4846 (
            .O(N__39465),
            .I(N__39459));
    Span4Mux_v I__4845 (
            .O(N__39462),
            .I(N__39454));
    LocalMux I__4844 (
            .O(N__39459),
            .I(N__39454));
    Span4Mux_v I__4843 (
            .O(N__39454),
            .I(N__39451));
    Span4Mux_h I__4842 (
            .O(N__39451),
            .I(N__39448));
    Span4Mux_v I__4841 (
            .O(N__39448),
            .I(N__39445));
    Odrv4 I__4840 (
            .O(N__39445),
            .I(\pid_alt.error_d_regZ0Z_8 ));
    InMux I__4839 (
            .O(N__39442),
            .I(N__39439));
    LocalMux I__4838 (
            .O(N__39439),
            .I(\pid_alt.error_d_reg_prev_esr_RNII5611_0Z0Z_8 ));
    CascadeMux I__4837 (
            .O(N__39436),
            .I(\pid_alt.error_d_reg_prev_esr_RNII5611_0Z0Z_8_cascade_ ));
    InMux I__4836 (
            .O(N__39433),
            .I(N__39428));
    InMux I__4835 (
            .O(N__39432),
            .I(N__39423));
    InMux I__4834 (
            .O(N__39431),
            .I(N__39423));
    LocalMux I__4833 (
            .O(N__39428),
            .I(N__39420));
    LocalMux I__4832 (
            .O(N__39423),
            .I(N__39417));
    Span4Mux_v I__4831 (
            .O(N__39420),
            .I(N__39414));
    Span4Mux_h I__4830 (
            .O(N__39417),
            .I(N__39411));
    Odrv4 I__4829 (
            .O(N__39414),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ ));
    Odrv4 I__4828 (
            .O(N__39411),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ ));
    CascadeMux I__4827 (
            .O(N__39406),
            .I(N__39403));
    InMux I__4826 (
            .O(N__39403),
            .I(N__39399));
    CascadeMux I__4825 (
            .O(N__39402),
            .I(N__39396));
    LocalMux I__4824 (
            .O(N__39399),
            .I(N__39393));
    InMux I__4823 (
            .O(N__39396),
            .I(N__39390));
    Odrv4 I__4822 (
            .O(N__39393),
            .I(\pid_alt.error_d_reg_prev_esr_RNI7T3T2Z0Z_7 ));
    LocalMux I__4821 (
            .O(N__39390),
            .I(\pid_alt.error_d_reg_prev_esr_RNI7T3T2Z0Z_7 ));
    InMux I__4820 (
            .O(N__39385),
            .I(N__39379));
    InMux I__4819 (
            .O(N__39384),
            .I(N__39379));
    LocalMux I__4818 (
            .O(N__39379),
            .I(\pid_alt.error_d_reg_prev_esr_RNIF2611Z0Z_7 ));
    CascadeMux I__4817 (
            .O(N__39376),
            .I(\pid_alt.un1_reset_0_i_cascade_ ));
    InMux I__4816 (
            .O(N__39373),
            .I(N__39366));
    InMux I__4815 (
            .O(N__39372),
            .I(N__39366));
    InMux I__4814 (
            .O(N__39371),
            .I(N__39363));
    LocalMux I__4813 (
            .O(N__39366),
            .I(N__39360));
    LocalMux I__4812 (
            .O(N__39363),
            .I(N__39357));
    Odrv4 I__4811 (
            .O(N__39360),
            .I(\pid_alt.pid_preregZ0Z_8 ));
    Odrv4 I__4810 (
            .O(N__39357),
            .I(\pid_alt.pid_preregZ0Z_8 ));
    InMux I__4809 (
            .O(N__39352),
            .I(N__39345));
    InMux I__4808 (
            .O(N__39351),
            .I(N__39345));
    InMux I__4807 (
            .O(N__39350),
            .I(N__39342));
    LocalMux I__4806 (
            .O(N__39345),
            .I(N__39339));
    LocalMux I__4805 (
            .O(N__39342),
            .I(N__39336));
    Odrv4 I__4804 (
            .O(N__39339),
            .I(\pid_alt.pid_preregZ0Z_7 ));
    Odrv4 I__4803 (
            .O(N__39336),
            .I(\pid_alt.pid_preregZ0Z_7 ));
    CascadeMux I__4802 (
            .O(N__39331),
            .I(N__39326));
    CascadeMux I__4801 (
            .O(N__39330),
            .I(N__39323));
    InMux I__4800 (
            .O(N__39329),
            .I(N__39318));
    InMux I__4799 (
            .O(N__39326),
            .I(N__39318));
    InMux I__4798 (
            .O(N__39323),
            .I(N__39315));
    LocalMux I__4797 (
            .O(N__39318),
            .I(N__39312));
    LocalMux I__4796 (
            .O(N__39315),
            .I(N__39309));
    Odrv4 I__4795 (
            .O(N__39312),
            .I(\pid_alt.pid_preregZ0Z_9 ));
    Odrv4 I__4794 (
            .O(N__39309),
            .I(\pid_alt.pid_preregZ0Z_9 ));
    InMux I__4793 (
            .O(N__39304),
            .I(N__39298));
    InMux I__4792 (
            .O(N__39303),
            .I(N__39298));
    LocalMux I__4791 (
            .O(N__39298),
            .I(N__39294));
    InMux I__4790 (
            .O(N__39297),
            .I(N__39291));
    Odrv4 I__4789 (
            .O(N__39294),
            .I(\pid_alt.pid_preregZ0Z_6 ));
    LocalMux I__4788 (
            .O(N__39291),
            .I(\pid_alt.pid_preregZ0Z_6 ));
    InMux I__4787 (
            .O(N__39286),
            .I(N__39279));
    InMux I__4786 (
            .O(N__39285),
            .I(N__39279));
    InMux I__4785 (
            .O(N__39284),
            .I(N__39276));
    LocalMux I__4784 (
            .O(N__39279),
            .I(N__39271));
    LocalMux I__4783 (
            .O(N__39276),
            .I(N__39271));
    Odrv4 I__4782 (
            .O(N__39271),
            .I(\pid_alt.pid_preregZ0Z_11 ));
    CascadeMux I__4781 (
            .O(N__39268),
            .I(\pid_alt.source_pid_1_sqmuxa_0_o2_3_cascade_ ));
    InMux I__4780 (
            .O(N__39265),
            .I(N__39258));
    InMux I__4779 (
            .O(N__39264),
            .I(N__39258));
    InMux I__4778 (
            .O(N__39263),
            .I(N__39255));
    LocalMux I__4777 (
            .O(N__39258),
            .I(N__39252));
    LocalMux I__4776 (
            .O(N__39255),
            .I(N__39249));
    Odrv4 I__4775 (
            .O(N__39252),
            .I(\pid_alt.pid_preregZ0Z_10 ));
    Odrv4 I__4774 (
            .O(N__39249),
            .I(\pid_alt.pid_preregZ0Z_10 ));
    InMux I__4773 (
            .O(N__39244),
            .I(N__39240));
    InMux I__4772 (
            .O(N__39243),
            .I(N__39237));
    LocalMux I__4771 (
            .O(N__39240),
            .I(\pid_alt.N_51 ));
    LocalMux I__4770 (
            .O(N__39237),
            .I(\pid_alt.N_51 ));
    CascadeMux I__4769 (
            .O(N__39232),
            .I(N__39229));
    InMux I__4768 (
            .O(N__39229),
            .I(N__39223));
    InMux I__4767 (
            .O(N__39228),
            .I(N__39223));
    LocalMux I__4766 (
            .O(N__39223),
            .I(\pid_alt.source_pid_1_sqmuxa_0_a2_0_2 ));
    InMux I__4765 (
            .O(N__39220),
            .I(N__39217));
    LocalMux I__4764 (
            .O(N__39217),
            .I(\pid_alt.source_pid_1_sqmuxa_0_a2_1_5 ));
    InMux I__4763 (
            .O(N__39214),
            .I(N__39211));
    LocalMux I__4762 (
            .O(N__39211),
            .I(\pid_alt.source_pid_1_sqmuxa_0_a2_1_7 ));
    InMux I__4761 (
            .O(N__39208),
            .I(N__39205));
    LocalMux I__4760 (
            .O(N__39205),
            .I(N__39202));
    Span4Mux_h I__4759 (
            .O(N__39202),
            .I(N__39199));
    Odrv4 I__4758 (
            .O(N__39199),
            .I(\pid_alt.pid_preregZ0Z_22 ));
    InMux I__4757 (
            .O(N__39196),
            .I(N__39193));
    LocalMux I__4756 (
            .O(N__39193),
            .I(N__39190));
    Odrv4 I__4755 (
            .O(N__39190),
            .I(\pid_alt.pid_preregZ0Z_19 ));
    CascadeMux I__4754 (
            .O(N__39187),
            .I(N__39184));
    InMux I__4753 (
            .O(N__39184),
            .I(N__39181));
    LocalMux I__4752 (
            .O(N__39181),
            .I(N__39178));
    Span4Mux_h I__4751 (
            .O(N__39178),
            .I(N__39175));
    Odrv4 I__4750 (
            .O(N__39175),
            .I(\pid_alt.pid_preregZ0Z_20 ));
    InMux I__4749 (
            .O(N__39172),
            .I(N__39169));
    LocalMux I__4748 (
            .O(N__39169),
            .I(N__39166));
    Odrv4 I__4747 (
            .O(N__39166),
            .I(\pid_alt.pid_preregZ0Z_17 ));
    InMux I__4746 (
            .O(N__39163),
            .I(N__39160));
    LocalMux I__4745 (
            .O(N__39160),
            .I(N__39157));
    Odrv4 I__4744 (
            .O(N__39157),
            .I(\pid_alt.pid_preregZ0Z_23 ));
    InMux I__4743 (
            .O(N__39154),
            .I(N__39151));
    LocalMux I__4742 (
            .O(N__39151),
            .I(N__39148));
    Odrv4 I__4741 (
            .O(N__39148),
            .I(\pid_alt.pid_preregZ0Z_18 ));
    CascadeMux I__4740 (
            .O(N__39145),
            .I(N__39142));
    InMux I__4739 (
            .O(N__39142),
            .I(N__39139));
    LocalMux I__4738 (
            .O(N__39139),
            .I(N__39136));
    Span4Mux_h I__4737 (
            .O(N__39136),
            .I(N__39133));
    Odrv4 I__4736 (
            .O(N__39133),
            .I(\pid_alt.pid_preregZ0Z_21 ));
    InMux I__4735 (
            .O(N__39130),
            .I(N__39127));
    LocalMux I__4734 (
            .O(N__39127),
            .I(N__39124));
    Odrv4 I__4733 (
            .O(N__39124),
            .I(\pid_alt.pid_preregZ0Z_15 ));
    InMux I__4732 (
            .O(N__39121),
            .I(N__39118));
    LocalMux I__4731 (
            .O(N__39118),
            .I(N__39115));
    Span4Mux_h I__4730 (
            .O(N__39115),
            .I(N__39112));
    Odrv4 I__4729 (
            .O(N__39112),
            .I(\pid_alt.pid_preregZ0Z_16 ));
    InMux I__4728 (
            .O(N__39109),
            .I(N__39106));
    LocalMux I__4727 (
            .O(N__39106),
            .I(\pid_alt.pid_preregZ0Z_14 ));
    CascadeMux I__4726 (
            .O(N__39103),
            .I(\pid_alt.source_pid_1_sqmuxa_0_a2_2_5_cascade_ ));
    InMux I__4725 (
            .O(N__39100),
            .I(N__39097));
    LocalMux I__4724 (
            .O(N__39097),
            .I(\pid_alt.source_pid_1_sqmuxa_0_a2_2_6 ));
    CascadeMux I__4723 (
            .O(N__39094),
            .I(\pid_alt.N_539_cascade_ ));
    CascadeMux I__4722 (
            .O(N__39091),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_9_cascade_ ));
    InMux I__4721 (
            .O(N__39088),
            .I(N__39085));
    LocalMux I__4720 (
            .O(N__39085),
            .I(\ppm_encoder_1.N_454 ));
    InMux I__4719 (
            .O(N__39082),
            .I(N__39079));
    LocalMux I__4718 (
            .O(N__39079),
            .I(\ppm_encoder_1.un2_throttle_iv_0_1_9 ));
    CascadeMux I__4717 (
            .O(N__39076),
            .I(N__39072));
    CascadeMux I__4716 (
            .O(N__39075),
            .I(N__39069));
    InMux I__4715 (
            .O(N__39072),
            .I(N__39066));
    InMux I__4714 (
            .O(N__39069),
            .I(N__39063));
    LocalMux I__4713 (
            .O(N__39066),
            .I(\ppm_encoder_1.throttleZ0Z_13 ));
    LocalMux I__4712 (
            .O(N__39063),
            .I(\ppm_encoder_1.throttleZ0Z_13 ));
    CascadeMux I__4711 (
            .O(N__39058),
            .I(\pid_alt.source_pid_1_sqmuxa_0_a2_0_3_cascade_ ));
    CascadeMux I__4710 (
            .O(N__39055),
            .I(\pid_alt.N_57_cascade_ ));
    CascadeMux I__4709 (
            .O(N__39052),
            .I(\pid_alt.un1_reset_1_cascade_ ));
    InMux I__4708 (
            .O(N__39049),
            .I(N__39046));
    LocalMux I__4707 (
            .O(N__39046),
            .I(\ppm_encoder_1.un2_throttle_iv_0_1_8 ));
    CascadeMux I__4706 (
            .O(N__39043),
            .I(N__39038));
    InMux I__4705 (
            .O(N__39042),
            .I(N__39035));
    InMux I__4704 (
            .O(N__39041),
            .I(N__39032));
    InMux I__4703 (
            .O(N__39038),
            .I(N__39029));
    LocalMux I__4702 (
            .O(N__39035),
            .I(\ppm_encoder_1.throttleZ0Z_4 ));
    LocalMux I__4701 (
            .O(N__39032),
            .I(\ppm_encoder_1.throttleZ0Z_4 ));
    LocalMux I__4700 (
            .O(N__39029),
            .I(\ppm_encoder_1.throttleZ0Z_4 ));
    InMux I__4699 (
            .O(N__39022),
            .I(N__39019));
    LocalMux I__4698 (
            .O(N__39019),
            .I(\ppm_encoder_1.un2_throttle_iv_0_1_4 ));
    CascadeMux I__4697 (
            .O(N__39016),
            .I(\ppm_encoder_1.N_260_i_cascade_ ));
    CascadeMux I__4696 (
            .O(N__39013),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_4_cascade_ ));
    CascadeMux I__4695 (
            .O(N__39010),
            .I(\ppm_encoder_1.un2_throttle_iv_0_2_9_cascade_ ));
    CascadeMux I__4694 (
            .O(N__39007),
            .I(\ppm_encoder_1.N_303_cascade_ ));
    InMux I__4693 (
            .O(N__39004),
            .I(N__39001));
    LocalMux I__4692 (
            .O(N__39001),
            .I(\ppm_encoder_1.un2_throttle_iv_0_2_2 ));
    CascadeMux I__4691 (
            .O(N__38998),
            .I(\ppm_encoder_1.N_448_cascade_ ));
    CascadeMux I__4690 (
            .O(N__38995),
            .I(N__38991));
    InMux I__4689 (
            .O(N__38994),
            .I(N__38983));
    InMux I__4688 (
            .O(N__38991),
            .I(N__38983));
    InMux I__4687 (
            .O(N__38990),
            .I(N__38983));
    LocalMux I__4686 (
            .O(N__38983),
            .I(\ppm_encoder_1.elevatorZ0Z_12 ));
    CascadeMux I__4685 (
            .O(N__38980),
            .I(\ppm_encoder_1.un2_throttle_iv_0_2_3_cascade_ ));
    InMux I__4684 (
            .O(N__38977),
            .I(N__38974));
    LocalMux I__4683 (
            .O(N__38974),
            .I(\ppm_encoder_1.un2_throttle_iv_0_1_3 ));
    CascadeMux I__4682 (
            .O(N__38971),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_3_cascade_ ));
    CascadeMux I__4681 (
            .O(N__38968),
            .I(\ppm_encoder_1.aileron_RNI7E8E1Z0Z_1_cascade_ ));
    CascadeMux I__4680 (
            .O(N__38965),
            .I(\ppm_encoder_1.un2_throttle_iv_0_1_1_cascade_ ));
    InMux I__4679 (
            .O(N__38962),
            .I(N__38959));
    LocalMux I__4678 (
            .O(N__38959),
            .I(\ppm_encoder_1.un2_throttle_iv_0_0_1 ));
    CascadeMux I__4677 (
            .O(N__38956),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_1_cascade_ ));
    InMux I__4676 (
            .O(N__38953),
            .I(N__38944));
    InMux I__4675 (
            .O(N__38952),
            .I(N__38941));
    InMux I__4674 (
            .O(N__38951),
            .I(N__38938));
    InMux I__4673 (
            .O(N__38950),
            .I(N__38933));
    InMux I__4672 (
            .O(N__38949),
            .I(N__38933));
    InMux I__4671 (
            .O(N__38948),
            .I(N__38928));
    InMux I__4670 (
            .O(N__38947),
            .I(N__38928));
    LocalMux I__4669 (
            .O(N__38944),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ));
    LocalMux I__4668 (
            .O(N__38941),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ));
    LocalMux I__4667 (
            .O(N__38938),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ));
    LocalMux I__4666 (
            .O(N__38933),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ));
    LocalMux I__4665 (
            .O(N__38928),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ));
    InMux I__4664 (
            .O(N__38917),
            .I(N__38911));
    InMux I__4663 (
            .O(N__38916),
            .I(N__38904));
    InMux I__4662 (
            .O(N__38915),
            .I(N__38904));
    InMux I__4661 (
            .O(N__38914),
            .I(N__38904));
    LocalMux I__4660 (
            .O(N__38911),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1 ));
    LocalMux I__4659 (
            .O(N__38904),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1 ));
    InMux I__4658 (
            .O(N__38899),
            .I(N__38893));
    InMux I__4657 (
            .O(N__38898),
            .I(N__38886));
    InMux I__4656 (
            .O(N__38897),
            .I(N__38886));
    InMux I__4655 (
            .O(N__38896),
            .I(N__38886));
    LocalMux I__4654 (
            .O(N__38893),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ));
    LocalMux I__4653 (
            .O(N__38886),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ));
    CascadeMux I__4652 (
            .O(N__38881),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI6LFQZ0Z_0_cascade_ ));
    InMux I__4651 (
            .O(N__38878),
            .I(N__38875));
    LocalMux I__4650 (
            .O(N__38875),
            .I(N__38872));
    Odrv4 I__4649 (
            .O(N__38872),
            .I(\ppm_encoder_1.PPM_STATE_fastZ0Z_0 ));
    CascadeMux I__4648 (
            .O(N__38869),
            .I(\ppm_encoder_1.PPM_STATE_fast_RNICIABZ0Z_0_cascade_ ));
    CascadeMux I__4647 (
            .O(N__38866),
            .I(N__38862));
    InMux I__4646 (
            .O(N__38865),
            .I(N__38858));
    InMux I__4645 (
            .O(N__38862),
            .I(N__38855));
    InMux I__4644 (
            .O(N__38861),
            .I(N__38852));
    LocalMux I__4643 (
            .O(N__38858),
            .I(N__38849));
    LocalMux I__4642 (
            .O(N__38855),
            .I(N__38846));
    LocalMux I__4641 (
            .O(N__38852),
            .I(N__38843));
    Span4Mux_v I__4640 (
            .O(N__38849),
            .I(N__38840));
    Span4Mux_h I__4639 (
            .O(N__38846),
            .I(N__38837));
    Odrv4 I__4638 (
            .O(N__38843),
            .I(\pid_alt.error_i_acumm_esr_RNIQMD91Z0Z_1 ));
    Odrv4 I__4637 (
            .O(N__38840),
            .I(\pid_alt.error_i_acumm_esr_RNIQMD91Z0Z_1 ));
    Odrv4 I__4636 (
            .O(N__38837),
            .I(\pid_alt.error_i_acumm_esr_RNIQMD91Z0Z_1 ));
    CascadeMux I__4635 (
            .O(N__38830),
            .I(N__38827));
    InMux I__4634 (
            .O(N__38827),
            .I(N__38824));
    LocalMux I__4633 (
            .O(N__38824),
            .I(N__38820));
    InMux I__4632 (
            .O(N__38823),
            .I(N__38817));
    Odrv12 I__4631 (
            .O(N__38820),
            .I(\pid_alt.error_i_acumm_preregZ0Z_1 ));
    LocalMux I__4630 (
            .O(N__38817),
            .I(\pid_alt.error_i_acumm_preregZ0Z_1 ));
    CascadeMux I__4629 (
            .O(N__38812),
            .I(\pid_alt.m21_e_0_cascade_ ));
    InMux I__4628 (
            .O(N__38809),
            .I(N__38795));
    InMux I__4627 (
            .O(N__38808),
            .I(N__38795));
    InMux I__4626 (
            .O(N__38807),
            .I(N__38795));
    InMux I__4625 (
            .O(N__38806),
            .I(N__38795));
    InMux I__4624 (
            .O(N__38805),
            .I(N__38792));
    InMux I__4623 (
            .O(N__38804),
            .I(N__38789));
    LocalMux I__4622 (
            .O(N__38795),
            .I(\pid_alt.error_i_acumm7lto4 ));
    LocalMux I__4621 (
            .O(N__38792),
            .I(\pid_alt.error_i_acumm7lto4 ));
    LocalMux I__4620 (
            .O(N__38789),
            .I(\pid_alt.error_i_acumm7lto4 ));
    InMux I__4619 (
            .O(N__38782),
            .I(N__38779));
    LocalMux I__4618 (
            .O(N__38779),
            .I(\pid_alt.m21_e_9 ));
    InMux I__4617 (
            .O(N__38776),
            .I(N__38773));
    LocalMux I__4616 (
            .O(N__38773),
            .I(N__38769));
    CascadeMux I__4615 (
            .O(N__38772),
            .I(N__38766));
    Span4Mux_h I__4614 (
            .O(N__38769),
            .I(N__38763));
    InMux I__4613 (
            .O(N__38766),
            .I(N__38760));
    Span4Mux_v I__4612 (
            .O(N__38763),
            .I(N__38757));
    LocalMux I__4611 (
            .O(N__38760),
            .I(N__38754));
    Span4Mux_v I__4610 (
            .O(N__38757),
            .I(N__38751));
    Span4Mux_v I__4609 (
            .O(N__38754),
            .I(N__38748));
    Odrv4 I__4608 (
            .O(N__38751),
            .I(\pid_alt.error_i_regZ0Z_0 ));
    Odrv4 I__4607 (
            .O(N__38748),
            .I(\pid_alt.error_i_regZ0Z_0 ));
    InMux I__4606 (
            .O(N__38743),
            .I(N__38739));
    InMux I__4605 (
            .O(N__38742),
            .I(N__38736));
    LocalMux I__4604 (
            .O(N__38739),
            .I(N__38733));
    LocalMux I__4603 (
            .O(N__38736),
            .I(N__38730));
    Odrv4 I__4602 (
            .O(N__38733),
            .I(\pid_alt.error_i_acummZ0Z_0 ));
    Odrv12 I__4601 (
            .O(N__38730),
            .I(\pid_alt.error_i_acummZ0Z_0 ));
    InMux I__4600 (
            .O(N__38725),
            .I(N__38722));
    LocalMux I__4599 (
            .O(N__38722),
            .I(N__38718));
    InMux I__4598 (
            .O(N__38721),
            .I(N__38715));
    Odrv4 I__4597 (
            .O(N__38718),
            .I(\pid_alt.error_i_acumm_preregZ0Z_0 ));
    LocalMux I__4596 (
            .O(N__38715),
            .I(\pid_alt.error_i_acumm_preregZ0Z_0 ));
    CascadeMux I__4595 (
            .O(N__38710),
            .I(N__38707));
    InMux I__4594 (
            .O(N__38707),
            .I(N__38704));
    LocalMux I__4593 (
            .O(N__38704),
            .I(N__38701));
    Span4Mux_h I__4592 (
            .O(N__38701),
            .I(N__38696));
    InMux I__4591 (
            .O(N__38700),
            .I(N__38691));
    InMux I__4590 (
            .O(N__38699),
            .I(N__38691));
    Odrv4 I__4589 (
            .O(N__38696),
            .I(\pid_alt.error_i_acumm_preregZ0Z_7 ));
    LocalMux I__4588 (
            .O(N__38691),
            .I(\pid_alt.error_i_acumm_preregZ0Z_7 ));
    InMux I__4587 (
            .O(N__38686),
            .I(N__38683));
    LocalMux I__4586 (
            .O(N__38683),
            .I(N__38679));
    InMux I__4585 (
            .O(N__38682),
            .I(N__38676));
    Span4Mux_h I__4584 (
            .O(N__38679),
            .I(N__38672));
    LocalMux I__4583 (
            .O(N__38676),
            .I(N__38669));
    InMux I__4582 (
            .O(N__38675),
            .I(N__38666));
    Odrv4 I__4581 (
            .O(N__38672),
            .I(\pid_alt.error_i_acumm_preregZ0Z_6 ));
    Odrv12 I__4580 (
            .O(N__38669),
            .I(\pid_alt.error_i_acumm_preregZ0Z_6 ));
    LocalMux I__4579 (
            .O(N__38666),
            .I(\pid_alt.error_i_acumm_preregZ0Z_6 ));
    InMux I__4578 (
            .O(N__38659),
            .I(N__38652));
    InMux I__4577 (
            .O(N__38658),
            .I(N__38652));
    InMux I__4576 (
            .O(N__38657),
            .I(N__38649));
    LocalMux I__4575 (
            .O(N__38652),
            .I(N__38646));
    LocalMux I__4574 (
            .O(N__38649),
            .I(\pid_alt.m35_e_2 ));
    Odrv4 I__4573 (
            .O(N__38646),
            .I(\pid_alt.m35_e_2 ));
    InMux I__4572 (
            .O(N__38641),
            .I(N__38638));
    LocalMux I__4571 (
            .O(N__38638),
            .I(N__38635));
    Span4Mux_h I__4570 (
            .O(N__38635),
            .I(N__38630));
    InMux I__4569 (
            .O(N__38634),
            .I(N__38625));
    InMux I__4568 (
            .O(N__38633),
            .I(N__38625));
    Span4Mux_v I__4567 (
            .O(N__38630),
            .I(N__38620));
    LocalMux I__4566 (
            .O(N__38625),
            .I(N__38620));
    Odrv4 I__4565 (
            .O(N__38620),
            .I(\pid_alt.error_i_reg_esr_RNIT8KA1Z0Z_5 ));
    CascadeMux I__4564 (
            .O(N__38617),
            .I(N__38612));
    CascadeMux I__4563 (
            .O(N__38616),
            .I(N__38609));
    CascadeMux I__4562 (
            .O(N__38615),
            .I(N__38605));
    InMux I__4561 (
            .O(N__38612),
            .I(N__38602));
    InMux I__4560 (
            .O(N__38609),
            .I(N__38599));
    CascadeMux I__4559 (
            .O(N__38608),
            .I(N__38596));
    InMux I__4558 (
            .O(N__38605),
            .I(N__38593));
    LocalMux I__4557 (
            .O(N__38602),
            .I(N__38590));
    LocalMux I__4556 (
            .O(N__38599),
            .I(N__38587));
    InMux I__4555 (
            .O(N__38596),
            .I(N__38584));
    LocalMux I__4554 (
            .O(N__38593),
            .I(N__38581));
    Span4Mux_v I__4553 (
            .O(N__38590),
            .I(N__38571));
    Span4Mux_v I__4552 (
            .O(N__38587),
            .I(N__38571));
    LocalMux I__4551 (
            .O(N__38584),
            .I(N__38571));
    Span4Mux_v I__4550 (
            .O(N__38581),
            .I(N__38571));
    InMux I__4549 (
            .O(N__38580),
            .I(N__38568));
    Odrv4 I__4548 (
            .O(N__38571),
            .I(\pid_alt.error_i_acumm7lto5 ));
    LocalMux I__4547 (
            .O(N__38568),
            .I(\pid_alt.error_i_acumm7lto5 ));
    InMux I__4546 (
            .O(N__38563),
            .I(N__38560));
    LocalMux I__4545 (
            .O(N__38560),
            .I(N__38557));
    Span12Mux_v I__4544 (
            .O(N__38557),
            .I(N__38554));
    Odrv12 I__4543 (
            .O(N__38554),
            .I(\pid_front.O_0_20 ));
    InMux I__4542 (
            .O(N__38551),
            .I(N__38548));
    LocalMux I__4541 (
            .O(N__38548),
            .I(N__38545));
    Span4Mux_v I__4540 (
            .O(N__38545),
            .I(N__38540));
    InMux I__4539 (
            .O(N__38544),
            .I(N__38537));
    InMux I__4538 (
            .O(N__38543),
            .I(N__38534));
    Span4Mux_v I__4537 (
            .O(N__38540),
            .I(N__38529));
    LocalMux I__4536 (
            .O(N__38537),
            .I(N__38529));
    LocalMux I__4535 (
            .O(N__38534),
            .I(N__38526));
    Span4Mux_h I__4534 (
            .O(N__38529),
            .I(N__38523));
    Span4Mux_h I__4533 (
            .O(N__38526),
            .I(N__38520));
    Span4Mux_v I__4532 (
            .O(N__38523),
            .I(N__38517));
    Span4Mux_v I__4531 (
            .O(N__38520),
            .I(N__38514));
    Odrv4 I__4530 (
            .O(N__38517),
            .I(\pid_alt.error_7 ));
    Odrv4 I__4529 (
            .O(N__38514),
            .I(\pid_alt.error_7 ));
    InMux I__4528 (
            .O(N__38509),
            .I(\pid_alt.error_cry_6 ));
    InMux I__4527 (
            .O(N__38506),
            .I(N__38501));
    InMux I__4526 (
            .O(N__38505),
            .I(N__38498));
    InMux I__4525 (
            .O(N__38504),
            .I(N__38495));
    LocalMux I__4524 (
            .O(N__38501),
            .I(N__38492));
    LocalMux I__4523 (
            .O(N__38498),
            .I(N__38489));
    LocalMux I__4522 (
            .O(N__38495),
            .I(N__38486));
    Span4Mux_v I__4521 (
            .O(N__38492),
            .I(N__38483));
    Span4Mux_v I__4520 (
            .O(N__38489),
            .I(N__38480));
    Span12Mux_s4_h I__4519 (
            .O(N__38486),
            .I(N__38477));
    Span4Mux_h I__4518 (
            .O(N__38483),
            .I(N__38474));
    Span4Mux_h I__4517 (
            .O(N__38480),
            .I(N__38471));
    Odrv12 I__4516 (
            .O(N__38477),
            .I(\pid_alt.error_8 ));
    Odrv4 I__4515 (
            .O(N__38474),
            .I(\pid_alt.error_8 ));
    Odrv4 I__4514 (
            .O(N__38471),
            .I(\pid_alt.error_8 ));
    InMux I__4513 (
            .O(N__38464),
            .I(bfn_4_19_0_));
    InMux I__4512 (
            .O(N__38461),
            .I(N__38458));
    LocalMux I__4511 (
            .O(N__38458),
            .I(N__38455));
    Span4Mux_v I__4510 (
            .O(N__38455),
            .I(N__38450));
    InMux I__4509 (
            .O(N__38454),
            .I(N__38447));
    InMux I__4508 (
            .O(N__38453),
            .I(N__38444));
    Span4Mux_v I__4507 (
            .O(N__38450),
            .I(N__38439));
    LocalMux I__4506 (
            .O(N__38447),
            .I(N__38439));
    LocalMux I__4505 (
            .O(N__38444),
            .I(N__38436));
    Span4Mux_h I__4504 (
            .O(N__38439),
            .I(N__38433));
    Span4Mux_h I__4503 (
            .O(N__38436),
            .I(N__38430));
    Span4Mux_v I__4502 (
            .O(N__38433),
            .I(N__38427));
    Span4Mux_v I__4501 (
            .O(N__38430),
            .I(N__38424));
    Odrv4 I__4500 (
            .O(N__38427),
            .I(\pid_alt.error_9 ));
    Odrv4 I__4499 (
            .O(N__38424),
            .I(\pid_alt.error_9 ));
    InMux I__4498 (
            .O(N__38419),
            .I(\pid_alt.error_cry_8 ));
    InMux I__4497 (
            .O(N__38416),
            .I(N__38413));
    LocalMux I__4496 (
            .O(N__38413),
            .I(N__38410));
    Span4Mux_s1_h I__4495 (
            .O(N__38410),
            .I(N__38405));
    InMux I__4494 (
            .O(N__38409),
            .I(N__38402));
    InMux I__4493 (
            .O(N__38408),
            .I(N__38399));
    Span4Mux_v I__4492 (
            .O(N__38405),
            .I(N__38394));
    LocalMux I__4491 (
            .O(N__38402),
            .I(N__38394));
    LocalMux I__4490 (
            .O(N__38399),
            .I(N__38391));
    Span4Mux_v I__4489 (
            .O(N__38394),
            .I(N__38388));
    Span4Mux_v I__4488 (
            .O(N__38391),
            .I(N__38385));
    Span4Mux_h I__4487 (
            .O(N__38388),
            .I(N__38382));
    Span4Mux_h I__4486 (
            .O(N__38385),
            .I(N__38379));
    Odrv4 I__4485 (
            .O(N__38382),
            .I(\pid_alt.error_10 ));
    Odrv4 I__4484 (
            .O(N__38379),
            .I(\pid_alt.error_10 ));
    InMux I__4483 (
            .O(N__38374),
            .I(\pid_alt.error_cry_9 ));
    InMux I__4482 (
            .O(N__38371),
            .I(N__38368));
    LocalMux I__4481 (
            .O(N__38368),
            .I(N__38363));
    InMux I__4480 (
            .O(N__38367),
            .I(N__38360));
    InMux I__4479 (
            .O(N__38366),
            .I(N__38357));
    Span4Mux_h I__4478 (
            .O(N__38363),
            .I(N__38354));
    LocalMux I__4477 (
            .O(N__38360),
            .I(N__38351));
    LocalMux I__4476 (
            .O(N__38357),
            .I(N__38348));
    Span4Mux_v I__4475 (
            .O(N__38354),
            .I(N__38345));
    Span4Mux_v I__4474 (
            .O(N__38351),
            .I(N__38342));
    Span4Mux_v I__4473 (
            .O(N__38348),
            .I(N__38339));
    Span4Mux_v I__4472 (
            .O(N__38345),
            .I(N__38334));
    Span4Mux_h I__4471 (
            .O(N__38342),
            .I(N__38334));
    Span4Mux_h I__4470 (
            .O(N__38339),
            .I(N__38331));
    Odrv4 I__4469 (
            .O(N__38334),
            .I(\pid_alt.error_11 ));
    Odrv4 I__4468 (
            .O(N__38331),
            .I(\pid_alt.error_11 ));
    InMux I__4467 (
            .O(N__38326),
            .I(\pid_alt.error_cry_10 ));
    InMux I__4466 (
            .O(N__38323),
            .I(N__38320));
    LocalMux I__4465 (
            .O(N__38320),
            .I(N__38315));
    InMux I__4464 (
            .O(N__38319),
            .I(N__38312));
    InMux I__4463 (
            .O(N__38318),
            .I(N__38309));
    Span4Mux_h I__4462 (
            .O(N__38315),
            .I(N__38306));
    LocalMux I__4461 (
            .O(N__38312),
            .I(N__38303));
    LocalMux I__4460 (
            .O(N__38309),
            .I(N__38300));
    Span4Mux_v I__4459 (
            .O(N__38306),
            .I(N__38297));
    Span4Mux_v I__4458 (
            .O(N__38303),
            .I(N__38294));
    Span4Mux_v I__4457 (
            .O(N__38300),
            .I(N__38291));
    Span4Mux_v I__4456 (
            .O(N__38297),
            .I(N__38286));
    Span4Mux_h I__4455 (
            .O(N__38294),
            .I(N__38286));
    Span4Mux_h I__4454 (
            .O(N__38291),
            .I(N__38283));
    Odrv4 I__4453 (
            .O(N__38286),
            .I(\pid_alt.error_12 ));
    Odrv4 I__4452 (
            .O(N__38283),
            .I(\pid_alt.error_12 ));
    InMux I__4451 (
            .O(N__38278),
            .I(\pid_alt.error_cry_11 ));
    InMux I__4450 (
            .O(N__38275),
            .I(N__38272));
    LocalMux I__4449 (
            .O(N__38272),
            .I(N__38267));
    InMux I__4448 (
            .O(N__38271),
            .I(N__38264));
    InMux I__4447 (
            .O(N__38270),
            .I(N__38261));
    Span4Mux_h I__4446 (
            .O(N__38267),
            .I(N__38258));
    LocalMux I__4445 (
            .O(N__38264),
            .I(N__38255));
    LocalMux I__4444 (
            .O(N__38261),
            .I(N__38252));
    Span4Mux_v I__4443 (
            .O(N__38258),
            .I(N__38249));
    Span4Mux_v I__4442 (
            .O(N__38255),
            .I(N__38246));
    Span4Mux_v I__4441 (
            .O(N__38252),
            .I(N__38243));
    Span4Mux_v I__4440 (
            .O(N__38249),
            .I(N__38238));
    Span4Mux_h I__4439 (
            .O(N__38246),
            .I(N__38238));
    Span4Mux_h I__4438 (
            .O(N__38243),
            .I(N__38235));
    Odrv4 I__4437 (
            .O(N__38238),
            .I(\pid_alt.error_13 ));
    Odrv4 I__4436 (
            .O(N__38235),
            .I(\pid_alt.error_13 ));
    InMux I__4435 (
            .O(N__38230),
            .I(\pid_alt.error_cry_12 ));
    InMux I__4434 (
            .O(N__38227),
            .I(N__38223));
    InMux I__4433 (
            .O(N__38226),
            .I(N__38219));
    LocalMux I__4432 (
            .O(N__38223),
            .I(N__38216));
    InMux I__4431 (
            .O(N__38222),
            .I(N__38213));
    LocalMux I__4430 (
            .O(N__38219),
            .I(N__38210));
    Span4Mux_h I__4429 (
            .O(N__38216),
            .I(N__38207));
    LocalMux I__4428 (
            .O(N__38213),
            .I(N__38204));
    Span12Mux_s2_h I__4427 (
            .O(N__38210),
            .I(N__38201));
    Span4Mux_v I__4426 (
            .O(N__38207),
            .I(N__38198));
    Span12Mux_s4_h I__4425 (
            .O(N__38204),
            .I(N__38195));
    Span12Mux_v I__4424 (
            .O(N__38201),
            .I(N__38192));
    Odrv4 I__4423 (
            .O(N__38198),
            .I(\pid_alt.error_14 ));
    Odrv12 I__4422 (
            .O(N__38195),
            .I(\pid_alt.error_14 ));
    Odrv12 I__4421 (
            .O(N__38192),
            .I(\pid_alt.error_14 ));
    InMux I__4420 (
            .O(N__38185),
            .I(\pid_alt.error_cry_13 ));
    InMux I__4419 (
            .O(N__38182),
            .I(\pid_alt.error_cry_14 ));
    InMux I__4418 (
            .O(N__38179),
            .I(N__38176));
    LocalMux I__4417 (
            .O(N__38176),
            .I(N__38173));
    Span4Mux_v I__4416 (
            .O(N__38173),
            .I(N__38168));
    InMux I__4415 (
            .O(N__38172),
            .I(N__38165));
    InMux I__4414 (
            .O(N__38171),
            .I(N__38162));
    Span4Mux_v I__4413 (
            .O(N__38168),
            .I(N__38157));
    LocalMux I__4412 (
            .O(N__38165),
            .I(N__38157));
    LocalMux I__4411 (
            .O(N__38162),
            .I(N__38154));
    Span4Mux_h I__4410 (
            .O(N__38157),
            .I(N__38151));
    Span4Mux_v I__4409 (
            .O(N__38154),
            .I(N__38148));
    Span4Mux_v I__4408 (
            .O(N__38151),
            .I(N__38145));
    Span4Mux_h I__4407 (
            .O(N__38148),
            .I(N__38142));
    Odrv4 I__4406 (
            .O(N__38145),
            .I(\pid_alt.error_15 ));
    Odrv4 I__4405 (
            .O(N__38142),
            .I(\pid_alt.error_15 ));
    CascadeMux I__4404 (
            .O(N__38137),
            .I(N__38134));
    InMux I__4403 (
            .O(N__38134),
            .I(N__38131));
    LocalMux I__4402 (
            .O(N__38131),
            .I(N__38127));
    InMux I__4401 (
            .O(N__38130),
            .I(N__38124));
    Span4Mux_h I__4400 (
            .O(N__38127),
            .I(N__38120));
    LocalMux I__4399 (
            .O(N__38124),
            .I(N__38117));
    InMux I__4398 (
            .O(N__38123),
            .I(N__38114));
    Odrv4 I__4397 (
            .O(N__38120),
            .I(\pid_alt.error_i_acumm_preregZ0Z_9 ));
    Odrv4 I__4396 (
            .O(N__38117),
            .I(\pid_alt.error_i_acumm_preregZ0Z_9 ));
    LocalMux I__4395 (
            .O(N__38114),
            .I(\pid_alt.error_i_acumm_preregZ0Z_9 ));
    InMux I__4394 (
            .O(N__38107),
            .I(N__38102));
    InMux I__4393 (
            .O(N__38106),
            .I(N__38099));
    InMux I__4392 (
            .O(N__38105),
            .I(N__38096));
    LocalMux I__4391 (
            .O(N__38102),
            .I(N__38093));
    LocalMux I__4390 (
            .O(N__38099),
            .I(N__38086));
    LocalMux I__4389 (
            .O(N__38096),
            .I(N__38086));
    Span4Mux_h I__4388 (
            .O(N__38093),
            .I(N__38086));
    Odrv4 I__4387 (
            .O(N__38086),
            .I(\pid_alt.error_i_acumm_preregZ0Z_8 ));
    CascadeMux I__4386 (
            .O(N__38083),
            .I(N__38078));
    CascadeMux I__4385 (
            .O(N__38082),
            .I(N__38075));
    InMux I__4384 (
            .O(N__38081),
            .I(N__38072));
    InMux I__4383 (
            .O(N__38078),
            .I(N__38069));
    InMux I__4382 (
            .O(N__38075),
            .I(N__38066));
    LocalMux I__4381 (
            .O(N__38072),
            .I(N__38061));
    LocalMux I__4380 (
            .O(N__38069),
            .I(N__38061));
    LocalMux I__4379 (
            .O(N__38066),
            .I(N__38058));
    Span4Mux_v I__4378 (
            .O(N__38061),
            .I(N__38055));
    Span4Mux_h I__4377 (
            .O(N__38058),
            .I(N__38052));
    Odrv4 I__4376 (
            .O(N__38055),
            .I(\pid_alt.error_i_acumm_preregZ0Z_11 ));
    Odrv4 I__4375 (
            .O(N__38052),
            .I(\pid_alt.error_i_acumm_preregZ0Z_11 ));
    InMux I__4374 (
            .O(N__38047),
            .I(N__38044));
    LocalMux I__4373 (
            .O(N__38044),
            .I(N__38041));
    Odrv4 I__4372 (
            .O(N__38041),
            .I(\pid_alt.m21_e_8 ));
    InMux I__4371 (
            .O(N__38038),
            .I(N__38035));
    LocalMux I__4370 (
            .O(N__38035),
            .I(N__38031));
    InMux I__4369 (
            .O(N__38034),
            .I(N__38028));
    Span4Mux_v I__4368 (
            .O(N__38031),
            .I(N__38022));
    LocalMux I__4367 (
            .O(N__38028),
            .I(N__38022));
    InMux I__4366 (
            .O(N__38027),
            .I(N__38019));
    Span4Mux_v I__4365 (
            .O(N__38022),
            .I(N__38016));
    LocalMux I__4364 (
            .O(N__38019),
            .I(N__38013));
    Span4Mux_v I__4363 (
            .O(N__38016),
            .I(N__38010));
    Span4Mux_v I__4362 (
            .O(N__38013),
            .I(N__38007));
    Span4Mux_h I__4361 (
            .O(N__38010),
            .I(N__38002));
    Span4Mux_h I__4360 (
            .O(N__38007),
            .I(N__38002));
    Span4Mux_v I__4359 (
            .O(N__38002),
            .I(N__37999));
    Odrv4 I__4358 (
            .O(N__37999),
            .I(\pid_alt.error_1 ));
    InMux I__4357 (
            .O(N__37996),
            .I(\pid_alt.error_cry_0 ));
    InMux I__4356 (
            .O(N__37993),
            .I(N__37990));
    LocalMux I__4355 (
            .O(N__37990),
            .I(N__37985));
    InMux I__4354 (
            .O(N__37989),
            .I(N__37982));
    InMux I__4353 (
            .O(N__37988),
            .I(N__37979));
    Span4Mux_v I__4352 (
            .O(N__37985),
            .I(N__37974));
    LocalMux I__4351 (
            .O(N__37982),
            .I(N__37974));
    LocalMux I__4350 (
            .O(N__37979),
            .I(N__37971));
    Span4Mux_v I__4349 (
            .O(N__37974),
            .I(N__37968));
    Span4Mux_v I__4348 (
            .O(N__37971),
            .I(N__37965));
    Span4Mux_h I__4347 (
            .O(N__37968),
            .I(N__37962));
    Span4Mux_h I__4346 (
            .O(N__37965),
            .I(N__37959));
    Odrv4 I__4345 (
            .O(N__37962),
            .I(\pid_alt.error_2 ));
    Odrv4 I__4344 (
            .O(N__37959),
            .I(\pid_alt.error_2 ));
    InMux I__4343 (
            .O(N__37954),
            .I(\pid_alt.error_cry_1 ));
    InMux I__4342 (
            .O(N__37951),
            .I(N__37948));
    LocalMux I__4341 (
            .O(N__37948),
            .I(N__37943));
    InMux I__4340 (
            .O(N__37947),
            .I(N__37940));
    InMux I__4339 (
            .O(N__37946),
            .I(N__37937));
    Span4Mux_h I__4338 (
            .O(N__37943),
            .I(N__37934));
    LocalMux I__4337 (
            .O(N__37940),
            .I(N__37931));
    LocalMux I__4336 (
            .O(N__37937),
            .I(N__37928));
    Span4Mux_v I__4335 (
            .O(N__37934),
            .I(N__37925));
    Span4Mux_v I__4334 (
            .O(N__37931),
            .I(N__37922));
    Span4Mux_v I__4333 (
            .O(N__37928),
            .I(N__37919));
    Span4Mux_v I__4332 (
            .O(N__37925),
            .I(N__37914));
    Span4Mux_h I__4331 (
            .O(N__37922),
            .I(N__37914));
    Span4Mux_h I__4330 (
            .O(N__37919),
            .I(N__37911));
    Odrv4 I__4329 (
            .O(N__37914),
            .I(\pid_alt.error_3 ));
    Odrv4 I__4328 (
            .O(N__37911),
            .I(\pid_alt.error_3 ));
    InMux I__4327 (
            .O(N__37906),
            .I(\pid_alt.error_cry_2 ));
    InMux I__4326 (
            .O(N__37903),
            .I(N__37900));
    LocalMux I__4325 (
            .O(N__37900),
            .I(N__37897));
    Span4Mux_v I__4324 (
            .O(N__37897),
            .I(N__37892));
    InMux I__4323 (
            .O(N__37896),
            .I(N__37889));
    InMux I__4322 (
            .O(N__37895),
            .I(N__37886));
    Span4Mux_v I__4321 (
            .O(N__37892),
            .I(N__37883));
    LocalMux I__4320 (
            .O(N__37889),
            .I(N__37880));
    LocalMux I__4319 (
            .O(N__37886),
            .I(N__37877));
    Span4Mux_h I__4318 (
            .O(N__37883),
            .I(N__37872));
    Span4Mux_h I__4317 (
            .O(N__37880),
            .I(N__37872));
    Span4Mux_v I__4316 (
            .O(N__37877),
            .I(N__37869));
    Span4Mux_v I__4315 (
            .O(N__37872),
            .I(N__37866));
    Span4Mux_h I__4314 (
            .O(N__37869),
            .I(N__37863));
    Odrv4 I__4313 (
            .O(N__37866),
            .I(\pid_alt.error_4 ));
    Odrv4 I__4312 (
            .O(N__37863),
            .I(\pid_alt.error_4 ));
    InMux I__4311 (
            .O(N__37858),
            .I(\pid_alt.error_cry_3 ));
    InMux I__4310 (
            .O(N__37855),
            .I(N__37852));
    LocalMux I__4309 (
            .O(N__37852),
            .I(N__37849));
    Span4Mux_v I__4308 (
            .O(N__37849),
            .I(N__37844));
    InMux I__4307 (
            .O(N__37848),
            .I(N__37841));
    InMux I__4306 (
            .O(N__37847),
            .I(N__37838));
    Span4Mux_v I__4305 (
            .O(N__37844),
            .I(N__37833));
    LocalMux I__4304 (
            .O(N__37841),
            .I(N__37833));
    LocalMux I__4303 (
            .O(N__37838),
            .I(N__37830));
    Span4Mux_h I__4302 (
            .O(N__37833),
            .I(N__37827));
    Span4Mux_v I__4301 (
            .O(N__37830),
            .I(N__37824));
    Span4Mux_v I__4300 (
            .O(N__37827),
            .I(N__37821));
    Span4Mux_h I__4299 (
            .O(N__37824),
            .I(N__37818));
    Odrv4 I__4298 (
            .O(N__37821),
            .I(\pid_alt.error_5 ));
    Odrv4 I__4297 (
            .O(N__37818),
            .I(\pid_alt.error_5 ));
    InMux I__4296 (
            .O(N__37813),
            .I(\pid_alt.error_cry_4 ));
    InMux I__4295 (
            .O(N__37810),
            .I(N__37807));
    LocalMux I__4294 (
            .O(N__37807),
            .I(N__37803));
    InMux I__4293 (
            .O(N__37806),
            .I(N__37799));
    Span4Mux_v I__4292 (
            .O(N__37803),
            .I(N__37796));
    InMux I__4291 (
            .O(N__37802),
            .I(N__37793));
    LocalMux I__4290 (
            .O(N__37799),
            .I(N__37790));
    Span4Mux_h I__4289 (
            .O(N__37796),
            .I(N__37787));
    LocalMux I__4288 (
            .O(N__37793),
            .I(N__37784));
    Span4Mux_h I__4287 (
            .O(N__37790),
            .I(N__37781));
    Sp12to4 I__4286 (
            .O(N__37787),
            .I(N__37776));
    Span12Mux_s4_h I__4285 (
            .O(N__37784),
            .I(N__37776));
    Span4Mux_v I__4284 (
            .O(N__37781),
            .I(N__37773));
    Odrv12 I__4283 (
            .O(N__37776),
            .I(\pid_alt.error_6 ));
    Odrv4 I__4282 (
            .O(N__37773),
            .I(\pid_alt.error_6 ));
    InMux I__4281 (
            .O(N__37768),
            .I(\pid_alt.error_cry_5 ));
    InMux I__4280 (
            .O(N__37765),
            .I(N__37760));
    InMux I__4279 (
            .O(N__37764),
            .I(N__37755));
    InMux I__4278 (
            .O(N__37763),
            .I(N__37755));
    LocalMux I__4277 (
            .O(N__37760),
            .I(N__37752));
    LocalMux I__4276 (
            .O(N__37755),
            .I(N__37749));
    Odrv4 I__4275 (
            .O(N__37752),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ ));
    Odrv4 I__4274 (
            .O(N__37749),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ ));
    InMux I__4273 (
            .O(N__37744),
            .I(N__37741));
    LocalMux I__4272 (
            .O(N__37741),
            .I(N__37738));
    Span4Mux_v I__4271 (
            .O(N__37738),
            .I(N__37733));
    InMux I__4270 (
            .O(N__37737),
            .I(N__37728));
    InMux I__4269 (
            .O(N__37736),
            .I(N__37728));
    Odrv4 I__4268 (
            .O(N__37733),
            .I(\pid_alt.error_i_reg_esr_RNIBKPJZ0Z_19 ));
    LocalMux I__4267 (
            .O(N__37728),
            .I(\pid_alt.error_i_reg_esr_RNIBKPJZ0Z_19 ));
    InMux I__4266 (
            .O(N__37723),
            .I(N__37720));
    LocalMux I__4265 (
            .O(N__37720),
            .I(N__37717));
    Span4Mux_v I__4264 (
            .O(N__37717),
            .I(N__37714));
    Odrv4 I__4263 (
            .O(N__37714),
            .I(\pid_alt.error_i_acumm_preregZ0Z_19 ));
    InMux I__4262 (
            .O(N__37711),
            .I(N__37708));
    LocalMux I__4261 (
            .O(N__37708),
            .I(N__37705));
    Odrv4 I__4260 (
            .O(N__37705),
            .I(\pid_alt.error_d_reg_prev_esr_RNIN49Q5Z0Z_8 ));
    InMux I__4259 (
            .O(N__37702),
            .I(N__37699));
    LocalMux I__4258 (
            .O(N__37699),
            .I(N__37695));
    InMux I__4257 (
            .O(N__37698),
            .I(N__37692));
    Span4Mux_h I__4256 (
            .O(N__37695),
            .I(N__37689));
    LocalMux I__4255 (
            .O(N__37692),
            .I(N__37686));
    Span4Mux_v I__4254 (
            .O(N__37689),
            .I(N__37683));
    Odrv12 I__4253 (
            .O(N__37686),
            .I(\pid_alt.error_p_regZ0Z_9 ));
    Odrv4 I__4252 (
            .O(N__37683),
            .I(\pid_alt.error_p_regZ0Z_9 ));
    InMux I__4251 (
            .O(N__37678),
            .I(N__37675));
    LocalMux I__4250 (
            .O(N__37675),
            .I(\pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9 ));
    CascadeMux I__4249 (
            .O(N__37672),
            .I(\pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9_cascade_ ));
    InMux I__4248 (
            .O(N__37669),
            .I(N__37665));
    CascadeMux I__4247 (
            .O(N__37668),
            .I(N__37662));
    LocalMux I__4246 (
            .O(N__37665),
            .I(N__37659));
    InMux I__4245 (
            .O(N__37662),
            .I(N__37656));
    Span4Mux_v I__4244 (
            .O(N__37659),
            .I(N__37653));
    LocalMux I__4243 (
            .O(N__37656),
            .I(N__37650));
    Odrv4 I__4242 (
            .O(N__37653),
            .I(\pid_alt.error_d_reg_prev_esr_RNIG75T2Z0Z_8 ));
    Odrv4 I__4241 (
            .O(N__37650),
            .I(\pid_alt.error_d_reg_prev_esr_RNIG75T2Z0Z_8 ));
    InMux I__4240 (
            .O(N__37645),
            .I(N__37639));
    InMux I__4239 (
            .O(N__37644),
            .I(N__37639));
    LocalMux I__4238 (
            .O(N__37639),
            .I(\pid_alt.error_d_reg_prev_esr_RNII5611Z0Z_8 ));
    InMux I__4237 (
            .O(N__37636),
            .I(N__37631));
    InMux I__4236 (
            .O(N__37635),
            .I(N__37626));
    InMux I__4235 (
            .O(N__37634),
            .I(N__37626));
    LocalMux I__4234 (
            .O(N__37631),
            .I(N__37623));
    LocalMux I__4233 (
            .O(N__37626),
            .I(N__37620));
    Span12Mux_v I__4232 (
            .O(N__37623),
            .I(N__37615));
    Span12Mux_h I__4231 (
            .O(N__37620),
            .I(N__37615));
    Odrv12 I__4230 (
            .O(N__37615),
            .I(\pid_alt.error_d_regZ0Z_9 ));
    InMux I__4229 (
            .O(N__37612),
            .I(N__37609));
    LocalMux I__4228 (
            .O(N__37609),
            .I(N__37606));
    Span4Mux_v I__4227 (
            .O(N__37606),
            .I(N__37602));
    InMux I__4226 (
            .O(N__37605),
            .I(N__37599));
    Odrv4 I__4225 (
            .O(N__37602),
            .I(\pid_alt.error_d_reg_prevZ0Z_9 ));
    LocalMux I__4224 (
            .O(N__37599),
            .I(\pid_alt.error_d_reg_prevZ0Z_9 ));
    InMux I__4223 (
            .O(N__37594),
            .I(N__37585));
    InMux I__4222 (
            .O(N__37593),
            .I(N__37585));
    InMux I__4221 (
            .O(N__37592),
            .I(N__37585));
    LocalMux I__4220 (
            .O(N__37585),
            .I(N__37582));
    Odrv4 I__4219 (
            .O(N__37582),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_8_c_RNI9POQ ));
    InMux I__4218 (
            .O(N__37579),
            .I(N__37576));
    LocalMux I__4217 (
            .O(N__37576),
            .I(N__37573));
    Span4Mux_h I__4216 (
            .O(N__37573),
            .I(N__37570));
    Odrv4 I__4215 (
            .O(N__37570),
            .I(\pid_alt.error_d_reg_prev_esr_RNIOVN14Z0Z_17 ));
    CascadeMux I__4214 (
            .O(N__37567),
            .I(N__37563));
    InMux I__4213 (
            .O(N__37566),
            .I(N__37560));
    InMux I__4212 (
            .O(N__37563),
            .I(N__37557));
    LocalMux I__4211 (
            .O(N__37560),
            .I(N__37554));
    LocalMux I__4210 (
            .O(N__37557),
            .I(N__37551));
    Span4Mux_v I__4209 (
            .O(N__37554),
            .I(N__37548));
    Span4Mux_h I__4208 (
            .O(N__37551),
            .I(N__37545));
    Odrv4 I__4207 (
            .O(N__37548),
            .I(\pid_alt.error_d_reg_prev_esr_RNI8BR02Z0Z_16 ));
    Odrv4 I__4206 (
            .O(N__37545),
            .I(\pid_alt.error_d_reg_prev_esr_RNI8BR02Z0Z_16 ));
    InMux I__4205 (
            .O(N__37540),
            .I(\pid_alt.un1_pid_prereg_0_cry_17 ));
    InMux I__4204 (
            .O(N__37537),
            .I(N__37534));
    LocalMux I__4203 (
            .O(N__37534),
            .I(N__37531));
    Odrv4 I__4202 (
            .O(N__37531),
            .I(\pid_alt.error_d_reg_prev_esr_RNI8IQ14Z0Z_18 ));
    CascadeMux I__4201 (
            .O(N__37528),
            .I(N__37525));
    InMux I__4200 (
            .O(N__37525),
            .I(N__37522));
    LocalMux I__4199 (
            .O(N__37522),
            .I(N__37518));
    InMux I__4198 (
            .O(N__37521),
            .I(N__37515));
    Span4Mux_h I__4197 (
            .O(N__37518),
            .I(N__37512));
    LocalMux I__4196 (
            .O(N__37515),
            .I(\pid_alt.error_d_reg_prev_esr_RNIGKS02Z0Z_17 ));
    Odrv4 I__4195 (
            .O(N__37512),
            .I(\pid_alt.error_d_reg_prev_esr_RNIGKS02Z0Z_17 ));
    InMux I__4194 (
            .O(N__37507),
            .I(\pid_alt.un1_pid_prereg_0_cry_18 ));
    InMux I__4193 (
            .O(N__37504),
            .I(N__37501));
    LocalMux I__4192 (
            .O(N__37501),
            .I(N__37498));
    Odrv4 I__4191 (
            .O(N__37498),
            .I(\pid_alt.error_d_reg_prev_esr_RNIK3024Z0Z_19 ));
    CascadeMux I__4190 (
            .O(N__37495),
            .I(N__37492));
    InMux I__4189 (
            .O(N__37492),
            .I(N__37488));
    InMux I__4188 (
            .O(N__37491),
            .I(N__37485));
    LocalMux I__4187 (
            .O(N__37488),
            .I(N__37482));
    LocalMux I__4186 (
            .O(N__37485),
            .I(\pid_alt.error_d_reg_prev_esr_RNIOTT02Z0Z_18 ));
    Odrv4 I__4185 (
            .O(N__37482),
            .I(\pid_alt.error_d_reg_prev_esr_RNIOTT02Z0Z_18 ));
    InMux I__4184 (
            .O(N__37477),
            .I(\pid_alt.un1_pid_prereg_0_cry_19 ));
    InMux I__4183 (
            .O(N__37474),
            .I(N__37471));
    LocalMux I__4182 (
            .O(N__37471),
            .I(N__37468));
    Span4Mux_h I__4181 (
            .O(N__37468),
            .I(N__37465));
    Odrv4 I__4180 (
            .O(N__37465),
            .I(\pid_alt.error_d_reg_prev_esr_RNICG9B1_0Z0Z_20 ));
    CascadeMux I__4179 (
            .O(N__37462),
            .I(N__37459));
    InMux I__4178 (
            .O(N__37459),
            .I(N__37456));
    LocalMux I__4177 (
            .O(N__37456),
            .I(N__37453));
    Odrv4 I__4176 (
            .O(N__37453),
            .I(\pid_alt.error_d_reg_prev_esr_RNIS5212Z0Z_19 ));
    InMux I__4175 (
            .O(N__37450),
            .I(\pid_alt.un1_pid_prereg_0_cry_20 ));
    InMux I__4174 (
            .O(N__37447),
            .I(N__37444));
    LocalMux I__4173 (
            .O(N__37444),
            .I(N__37441));
    Span4Mux_h I__4172 (
            .O(N__37441),
            .I(N__37438));
    Odrv4 I__4171 (
            .O(N__37438),
            .I(\pid_alt.error_d_reg_prev_esr_RNICG9B1_1Z0Z_20 ));
    InMux I__4170 (
            .O(N__37435),
            .I(\pid_alt.un1_pid_prereg_0_cry_21 ));
    CascadeMux I__4169 (
            .O(N__37432),
            .I(N__37428));
    InMux I__4168 (
            .O(N__37431),
            .I(N__37425));
    InMux I__4167 (
            .O(N__37428),
            .I(N__37422));
    LocalMux I__4166 (
            .O(N__37425),
            .I(N__37419));
    LocalMux I__4165 (
            .O(N__37422),
            .I(N__37416));
    Span4Mux_h I__4164 (
            .O(N__37419),
            .I(N__37413));
    Span4Mux_h I__4163 (
            .O(N__37416),
            .I(N__37410));
    Odrv4 I__4162 (
            .O(N__37413),
            .I(\pid_alt.error_d_reg_prev_esr_RNICG9B1Z0Z_20 ));
    Odrv4 I__4161 (
            .O(N__37410),
            .I(\pid_alt.error_d_reg_prev_esr_RNICG9B1Z0Z_20 ));
    CascadeMux I__4160 (
            .O(N__37405),
            .I(N__37402));
    InMux I__4159 (
            .O(N__37402),
            .I(N__37399));
    LocalMux I__4158 (
            .O(N__37399),
            .I(N__37396));
    Span12Mux_h I__4157 (
            .O(N__37396),
            .I(N__37393));
    Odrv12 I__4156 (
            .O(N__37393),
            .I(\pid_alt.error_d_reg_prev_esr_RNICG9B1_2Z0Z_20 ));
    InMux I__4155 (
            .O(N__37390),
            .I(bfn_4_16_0_));
    InMux I__4154 (
            .O(N__37387),
            .I(N__37384));
    LocalMux I__4153 (
            .O(N__37384),
            .I(N__37381));
    Span4Mux_h I__4152 (
            .O(N__37381),
            .I(N__37378));
    Odrv4 I__4151 (
            .O(N__37378),
            .I(\pid_alt.un1_pid_prereg_0_axb_24 ));
    InMux I__4150 (
            .O(N__37375),
            .I(\pid_alt.un1_pid_prereg_0_cry_23 ));
    InMux I__4149 (
            .O(N__37372),
            .I(N__37369));
    LocalMux I__4148 (
            .O(N__37369),
            .I(N__37366));
    Span4Mux_h I__4147 (
            .O(N__37366),
            .I(N__37361));
    InMux I__4146 (
            .O(N__37365),
            .I(N__37356));
    InMux I__4145 (
            .O(N__37364),
            .I(N__37356));
    Odrv4 I__4144 (
            .O(N__37361),
            .I(\pid_alt.error_i_reg_esr_RNI15KJZ0Z_14 ));
    LocalMux I__4143 (
            .O(N__37356),
            .I(\pid_alt.error_i_reg_esr_RNI15KJZ0Z_14 ));
    InMux I__4142 (
            .O(N__37351),
            .I(N__37345));
    InMux I__4141 (
            .O(N__37350),
            .I(N__37345));
    LocalMux I__4140 (
            .O(N__37345),
            .I(N__37342));
    Span4Mux_v I__4139 (
            .O(N__37342),
            .I(N__37339));
    Odrv4 I__4138 (
            .O(N__37339),
            .I(\pid_alt.error_i_acumm_preregZ0Z_14 ));
    InMux I__4137 (
            .O(N__37336),
            .I(N__37333));
    LocalMux I__4136 (
            .O(N__37333),
            .I(N__37330));
    Span4Mux_h I__4135 (
            .O(N__37330),
            .I(N__37327));
    Odrv4 I__4134 (
            .O(N__37327),
            .I(\pid_alt.error_d_reg_prev_esr_RNICI045Z0Z_9 ));
    InMux I__4133 (
            .O(N__37324),
            .I(\pid_alt.un1_pid_prereg_0_cry_9 ));
    InMux I__4132 (
            .O(N__37321),
            .I(N__37318));
    LocalMux I__4131 (
            .O(N__37318),
            .I(N__37315));
    Span4Mux_v I__4130 (
            .O(N__37315),
            .I(N__37312));
    Odrv4 I__4129 (
            .O(N__37312),
            .I(\pid_alt.error_d_reg_prev_esr_RNITPKD4Z0Z_10 ));
    CascadeMux I__4128 (
            .O(N__37309),
            .I(N__37306));
    InMux I__4127 (
            .O(N__37306),
            .I(N__37303));
    LocalMux I__4126 (
            .O(N__37303),
            .I(N__37300));
    Span4Mux_h I__4125 (
            .O(N__37300),
            .I(N__37296));
    InMux I__4124 (
            .O(N__37299),
            .I(N__37293));
    Span4Mux_v I__4123 (
            .O(N__37296),
            .I(N__37290));
    LocalMux I__4122 (
            .O(N__37293),
            .I(\pid_alt.error_d_reg_prev_esr_RNISAR62Z0Z_9 ));
    Odrv4 I__4121 (
            .O(N__37290),
            .I(\pid_alt.error_d_reg_prev_esr_RNISAR62Z0Z_9 ));
    InMux I__4120 (
            .O(N__37285),
            .I(\pid_alt.un1_pid_prereg_0_cry_10 ));
    InMux I__4119 (
            .O(N__37282),
            .I(N__37279));
    LocalMux I__4118 (
            .O(N__37279),
            .I(\pid_alt.error_d_reg_prev_esr_RNIB8KD4Z0Z_11 ));
    CascadeMux I__4117 (
            .O(N__37276),
            .I(N__37272));
    InMux I__4116 (
            .O(N__37275),
            .I(N__37269));
    InMux I__4115 (
            .O(N__37272),
            .I(N__37266));
    LocalMux I__4114 (
            .O(N__37269),
            .I(N__37263));
    LocalMux I__4113 (
            .O(N__37266),
            .I(N__37260));
    Span4Mux_v I__4112 (
            .O(N__37263),
            .I(N__37257));
    Span4Mux_h I__4111 (
            .O(N__37260),
            .I(N__37254));
    Odrv4 I__4110 (
            .O(N__37257),
            .I(\pid_alt.error_d_reg_prev_esr_RNI1FP62Z0Z_10 ));
    Odrv4 I__4109 (
            .O(N__37254),
            .I(\pid_alt.error_d_reg_prev_esr_RNI1FP62Z0Z_10 ));
    InMux I__4108 (
            .O(N__37249),
            .I(\pid_alt.un1_pid_prereg_0_cry_11 ));
    InMux I__4107 (
            .O(N__37246),
            .I(N__37243));
    LocalMux I__4106 (
            .O(N__37243),
            .I(\pid_alt.error_d_reg_prev_esr_RNI64JA4Z0Z_12 ));
    CascadeMux I__4105 (
            .O(N__37240),
            .I(N__37236));
    CascadeMux I__4104 (
            .O(N__37239),
            .I(N__37233));
    InMux I__4103 (
            .O(N__37236),
            .I(N__37230));
    InMux I__4102 (
            .O(N__37233),
            .I(N__37227));
    LocalMux I__4101 (
            .O(N__37230),
            .I(\pid_alt.error_d_reg_prev_esr_RNIAPQ62Z0Z_11 ));
    LocalMux I__4100 (
            .O(N__37227),
            .I(\pid_alt.error_d_reg_prev_esr_RNIAPQ62Z0Z_11 ));
    InMux I__4099 (
            .O(N__37222),
            .I(\pid_alt.un1_pid_prereg_0_cry_12 ));
    InMux I__4098 (
            .O(N__37219),
            .I(N__37216));
    LocalMux I__4097 (
            .O(N__37216),
            .I(N__37213));
    Odrv4 I__4096 (
            .O(N__37213),
            .I(\pid_alt.error_d_reg_prev_esr_RNICQF44Z0Z_13 ));
    CascadeMux I__4095 (
            .O(N__37210),
            .I(N__37206));
    InMux I__4094 (
            .O(N__37209),
            .I(N__37203));
    InMux I__4093 (
            .O(N__37206),
            .I(N__37200));
    LocalMux I__4092 (
            .O(N__37203),
            .I(\pid_alt.error_d_reg_prev_esr_RNISAO32Z0Z_12 ));
    LocalMux I__4091 (
            .O(N__37200),
            .I(\pid_alt.error_d_reg_prev_esr_RNISAO32Z0Z_12 ));
    InMux I__4090 (
            .O(N__37195),
            .I(\pid_alt.un1_pid_prereg_0_cry_13 ));
    InMux I__4089 (
            .O(N__37192),
            .I(N__37189));
    LocalMux I__4088 (
            .O(N__37189),
            .I(N__37186));
    Odrv4 I__4087 (
            .O(N__37186),
            .I(\pid_alt.error_d_reg_prev_esr_RNI88G14Z0Z_14 ));
    CascadeMux I__4086 (
            .O(N__37183),
            .I(N__37179));
    CascadeMux I__4085 (
            .O(N__37182),
            .I(N__37176));
    InMux I__4084 (
            .O(N__37179),
            .I(N__37173));
    InMux I__4083 (
            .O(N__37176),
            .I(N__37170));
    LocalMux I__4082 (
            .O(N__37173),
            .I(\pid_alt.error_d_reg_prev_esr_RNIGFN02Z0Z_13 ));
    LocalMux I__4081 (
            .O(N__37170),
            .I(\pid_alt.error_d_reg_prev_esr_RNIGFN02Z0Z_13 ));
    InMux I__4080 (
            .O(N__37165),
            .I(bfn_4_15_0_));
    InMux I__4079 (
            .O(N__37162),
            .I(N__37159));
    LocalMux I__4078 (
            .O(N__37159),
            .I(N__37156));
    Span4Mux_h I__4077 (
            .O(N__37156),
            .I(N__37153));
    Odrv4 I__4076 (
            .O(N__37153),
            .I(\pid_alt.error_d_reg_prev_esr_RNIOQI14Z0Z_15 ));
    CascadeMux I__4075 (
            .O(N__37150),
            .I(N__37147));
    InMux I__4074 (
            .O(N__37147),
            .I(N__37144));
    LocalMux I__4073 (
            .O(N__37144),
            .I(N__37140));
    CascadeMux I__4072 (
            .O(N__37143),
            .I(N__37137));
    Span4Mux_v I__4071 (
            .O(N__37140),
            .I(N__37134));
    InMux I__4070 (
            .O(N__37137),
            .I(N__37131));
    Odrv4 I__4069 (
            .O(N__37134),
            .I(\pid_alt.error_d_reg_prev_esr_RNIOOO02Z0Z_14 ));
    LocalMux I__4068 (
            .O(N__37131),
            .I(\pid_alt.error_d_reg_prev_esr_RNIOOO02Z0Z_14 ));
    InMux I__4067 (
            .O(N__37126),
            .I(\pid_alt.un1_pid_prereg_0_cry_15 ));
    InMux I__4066 (
            .O(N__37123),
            .I(N__37119));
    CascadeMux I__4065 (
            .O(N__37122),
            .I(N__37116));
    LocalMux I__4064 (
            .O(N__37119),
            .I(N__37113));
    InMux I__4063 (
            .O(N__37116),
            .I(N__37110));
    Span4Mux_h I__4062 (
            .O(N__37113),
            .I(N__37107));
    LocalMux I__4061 (
            .O(N__37110),
            .I(\pid_alt.error_d_reg_prev_esr_RNI02Q02Z0Z_15 ));
    Odrv4 I__4060 (
            .O(N__37107),
            .I(\pid_alt.error_d_reg_prev_esr_RNI02Q02Z0Z_15 ));
    CascadeMux I__4059 (
            .O(N__37102),
            .I(N__37099));
    InMux I__4058 (
            .O(N__37099),
            .I(N__37096));
    LocalMux I__4057 (
            .O(N__37096),
            .I(N__37093));
    Span4Mux_h I__4056 (
            .O(N__37093),
            .I(N__37090));
    Odrv4 I__4055 (
            .O(N__37090),
            .I(\pid_alt.error_d_reg_prev_esr_RNI8DL14Z0Z_16 ));
    InMux I__4054 (
            .O(N__37087),
            .I(\pid_alt.un1_pid_prereg_0_cry_16 ));
    InMux I__4053 (
            .O(N__37084),
            .I(N__37081));
    LocalMux I__4052 (
            .O(N__37081),
            .I(N__37078));
    Odrv4 I__4051 (
            .O(N__37078),
            .I(\pid_alt.error_d_reg_prev_esr_RNIF0465Z0Z_1 ));
    CascadeMux I__4050 (
            .O(N__37075),
            .I(N__37072));
    InMux I__4049 (
            .O(N__37072),
            .I(N__37067));
    InMux I__4048 (
            .O(N__37071),
            .I(N__37064));
    InMux I__4047 (
            .O(N__37070),
            .I(N__37061));
    LocalMux I__4046 (
            .O(N__37067),
            .I(N__37058));
    LocalMux I__4045 (
            .O(N__37064),
            .I(N__37055));
    LocalMux I__4044 (
            .O(N__37061),
            .I(N__37052));
    Span4Mux_h I__4043 (
            .O(N__37058),
            .I(N__37049));
    Odrv4 I__4042 (
            .O(N__37055),
            .I(\pid_alt.error_i_acumm_esr_RNITQE91Z0Z_2 ));
    Odrv4 I__4041 (
            .O(N__37052),
            .I(\pid_alt.error_i_acumm_esr_RNITQE91Z0Z_2 ));
    Odrv4 I__4040 (
            .O(N__37049),
            .I(\pid_alt.error_i_acumm_esr_RNITQE91Z0Z_2 ));
    InMux I__4039 (
            .O(N__37042),
            .I(N__37038));
    InMux I__4038 (
            .O(N__37041),
            .I(N__37035));
    LocalMux I__4037 (
            .O(N__37038),
            .I(\pid_alt.pid_preregZ0Z_2 ));
    LocalMux I__4036 (
            .O(N__37035),
            .I(\pid_alt.pid_preregZ0Z_2 ));
    InMux I__4035 (
            .O(N__37030),
            .I(\pid_alt.un1_pid_prereg_0_cry_1 ));
    InMux I__4034 (
            .O(N__37027),
            .I(N__37024));
    LocalMux I__4033 (
            .O(N__37024),
            .I(\pid_alt.error_d_reg_prev_esr_RNILDG87Z0Z_2 ));
    CascadeMux I__4032 (
            .O(N__37021),
            .I(N__37017));
    CascadeMux I__4031 (
            .O(N__37020),
            .I(N__37014));
    InMux I__4030 (
            .O(N__37017),
            .I(N__37010));
    InMux I__4029 (
            .O(N__37014),
            .I(N__37007));
    InMux I__4028 (
            .O(N__37013),
            .I(N__37004));
    LocalMux I__4027 (
            .O(N__37010),
            .I(N__37001));
    LocalMux I__4026 (
            .O(N__37007),
            .I(N__36998));
    LocalMux I__4025 (
            .O(N__37004),
            .I(N__36995));
    Span4Mux_h I__4024 (
            .O(N__37001),
            .I(N__36992));
    Odrv4 I__4023 (
            .O(N__36998),
            .I(\pid_alt.error_i_acumm_esr_RNI0VF91Z0Z_3 ));
    Odrv4 I__4022 (
            .O(N__36995),
            .I(\pid_alt.error_i_acumm_esr_RNI0VF91Z0Z_3 ));
    Odrv4 I__4021 (
            .O(N__36992),
            .I(\pid_alt.error_i_acumm_esr_RNI0VF91Z0Z_3 ));
    CascadeMux I__4020 (
            .O(N__36985),
            .I(N__36981));
    CascadeMux I__4019 (
            .O(N__36984),
            .I(N__36978));
    InMux I__4018 (
            .O(N__36981),
            .I(N__36975));
    InMux I__4017 (
            .O(N__36978),
            .I(N__36972));
    LocalMux I__4016 (
            .O(N__36975),
            .I(\pid_alt.pid_preregZ0Z_3 ));
    LocalMux I__4015 (
            .O(N__36972),
            .I(\pid_alt.pid_preregZ0Z_3 ));
    InMux I__4014 (
            .O(N__36967),
            .I(\pid_alt.un1_pid_prereg_0_cry_2 ));
    CascadeMux I__4013 (
            .O(N__36964),
            .I(N__36961));
    InMux I__4012 (
            .O(N__36961),
            .I(N__36958));
    LocalMux I__4011 (
            .O(N__36958),
            .I(N__36954));
    InMux I__4010 (
            .O(N__36957),
            .I(N__36951));
    Odrv4 I__4009 (
            .O(N__36954),
            .I(\pid_alt.error_d_reg_prev_esr_RNILE0V5Z0Z_2 ));
    LocalMux I__4008 (
            .O(N__36951),
            .I(\pid_alt.error_d_reg_prev_esr_RNILE0V5Z0Z_2 ));
    CascadeMux I__4007 (
            .O(N__36946),
            .I(N__36943));
    InMux I__4006 (
            .O(N__36943),
            .I(N__36940));
    LocalMux I__4005 (
            .O(N__36940),
            .I(\pid_alt.error_d_reg_prev_esr_RNI11TA9Z0Z_3 ));
    InMux I__4004 (
            .O(N__36937),
            .I(\pid_alt.un1_pid_prereg_0_cry_3 ));
    InMux I__4003 (
            .O(N__36934),
            .I(N__36931));
    LocalMux I__4002 (
            .O(N__36931),
            .I(\pid_alt.error_d_reg_prev_esr_RNIOGSO6Z0Z_4 ));
    CascadeMux I__4001 (
            .O(N__36928),
            .I(N__36924));
    InMux I__4000 (
            .O(N__36927),
            .I(N__36921));
    InMux I__3999 (
            .O(N__36924),
            .I(N__36918));
    LocalMux I__3998 (
            .O(N__36921),
            .I(\pid_alt.error_d_reg_prev_esr_RNICISB3Z0Z_3 ));
    LocalMux I__3997 (
            .O(N__36918),
            .I(\pid_alt.error_d_reg_prev_esr_RNICISB3Z0Z_3 ));
    InMux I__3996 (
            .O(N__36913),
            .I(\pid_alt.un1_pid_prereg_0_cry_4 ));
    InMux I__3995 (
            .O(N__36910),
            .I(N__36907));
    LocalMux I__3994 (
            .O(N__36907),
            .I(\pid_alt.error_d_reg_prev_esr_RNI171A6Z0Z_5 ));
    CascadeMux I__3993 (
            .O(N__36904),
            .I(N__36900));
    CascadeMux I__3992 (
            .O(N__36903),
            .I(N__36897));
    InMux I__3991 (
            .O(N__36900),
            .I(N__36894));
    InMux I__3990 (
            .O(N__36897),
            .I(N__36891));
    LocalMux I__3989 (
            .O(N__36894),
            .I(\pid_alt.error_d_reg_prev_esr_RNICUVC3Z0Z_4 ));
    LocalMux I__3988 (
            .O(N__36891),
            .I(\pid_alt.error_d_reg_prev_esr_RNICUVC3Z0Z_4 ));
    InMux I__3987 (
            .O(N__36886),
            .I(\pid_alt.un1_pid_prereg_0_cry_5 ));
    InMux I__3986 (
            .O(N__36883),
            .I(bfn_4_14_0_));
    InMux I__3985 (
            .O(N__36880),
            .I(\pid_alt.un1_pid_prereg_0_cry_7 ));
    InMux I__3984 (
            .O(N__36877),
            .I(\pid_alt.un1_pid_prereg_0_cry_8 ));
    CascadeMux I__3983 (
            .O(N__36874),
            .I(\pid_alt.N_54_cascade_ ));
    InMux I__3982 (
            .O(N__36871),
            .I(N__36867));
    InMux I__3981 (
            .O(N__36870),
            .I(N__36864));
    LocalMux I__3980 (
            .O(N__36867),
            .I(N__36861));
    LocalMux I__3979 (
            .O(N__36864),
            .I(N__36858));
    Odrv12 I__3978 (
            .O(N__36861),
            .I(throttle_order_1));
    Odrv4 I__3977 (
            .O(N__36858),
            .I(throttle_order_1));
    CascadeMux I__3976 (
            .O(N__36853),
            .I(N__36850));
    InMux I__3975 (
            .O(N__36850),
            .I(N__36847));
    LocalMux I__3974 (
            .O(N__36847),
            .I(N__36843));
    InMux I__3973 (
            .O(N__36846),
            .I(N__36840));
    Span4Mux_v I__3972 (
            .O(N__36843),
            .I(N__36835));
    LocalMux I__3971 (
            .O(N__36840),
            .I(N__36835));
    Odrv4 I__3970 (
            .O(N__36835),
            .I(throttle_order_2));
    CascadeMux I__3969 (
            .O(N__36832),
            .I(N__36828));
    InMux I__3968 (
            .O(N__36831),
            .I(N__36820));
    InMux I__3967 (
            .O(N__36828),
            .I(N__36820));
    InMux I__3966 (
            .O(N__36827),
            .I(N__36820));
    LocalMux I__3965 (
            .O(N__36820),
            .I(\pid_alt.N_54 ));
    InMux I__3964 (
            .O(N__36817),
            .I(N__36813));
    InMux I__3963 (
            .O(N__36816),
            .I(N__36810));
    LocalMux I__3962 (
            .O(N__36813),
            .I(N__36805));
    LocalMux I__3961 (
            .O(N__36810),
            .I(N__36805));
    Odrv12 I__3960 (
            .O(N__36805),
            .I(throttle_order_3));
    CascadeMux I__3959 (
            .O(N__36802),
            .I(N__36799));
    InMux I__3958 (
            .O(N__36799),
            .I(N__36796));
    LocalMux I__3957 (
            .O(N__36796),
            .I(N__36792));
    InMux I__3956 (
            .O(N__36795),
            .I(N__36789));
    Span4Mux_v I__3955 (
            .O(N__36792),
            .I(N__36786));
    LocalMux I__3954 (
            .O(N__36789),
            .I(N__36783));
    Span4Mux_h I__3953 (
            .O(N__36786),
            .I(N__36778));
    Span4Mux_v I__3952 (
            .O(N__36783),
            .I(N__36778));
    Odrv4 I__3951 (
            .O(N__36778),
            .I(\pid_alt.error_d_reg_prev_i_0 ));
    InMux I__3950 (
            .O(N__36775),
            .I(N__36772));
    LocalMux I__3949 (
            .O(N__36772),
            .I(N__36769));
    Span4Mux_v I__3948 (
            .O(N__36769),
            .I(N__36766));
    Odrv4 I__3947 (
            .O(N__36766),
            .I(\pid_alt.error_p_reg_esr_RNI3SMI1Z0Z_0 ));
    CascadeMux I__3946 (
            .O(N__36763),
            .I(N__36759));
    InMux I__3945 (
            .O(N__36762),
            .I(N__36756));
    InMux I__3944 (
            .O(N__36759),
            .I(N__36753));
    LocalMux I__3943 (
            .O(N__36756),
            .I(N__36750));
    LocalMux I__3942 (
            .O(N__36753),
            .I(N__36747));
    Span4Mux_s2_h I__3941 (
            .O(N__36750),
            .I(N__36744));
    Span4Mux_v I__3940 (
            .O(N__36747),
            .I(N__36741));
    Odrv4 I__3939 (
            .O(N__36744),
            .I(\pid_alt.un1_pid_prereg_0 ));
    Odrv4 I__3938 (
            .O(N__36741),
            .I(\pid_alt.un1_pid_prereg_0 ));
    InMux I__3937 (
            .O(N__36736),
            .I(N__36730));
    InMux I__3936 (
            .O(N__36735),
            .I(N__36730));
    LocalMux I__3935 (
            .O(N__36730),
            .I(\pid_alt.pid_preregZ0Z_0 ));
    InMux I__3934 (
            .O(N__36727),
            .I(\pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CO ));
    InMux I__3933 (
            .O(N__36724),
            .I(N__36721));
    LocalMux I__3932 (
            .O(N__36721),
            .I(N__36718));
    Span4Mux_h I__3931 (
            .O(N__36718),
            .I(N__36715));
    Odrv4 I__3930 (
            .O(N__36715),
            .I(\pid_alt.error_d_reg_prev_esr_RNIFPN33Z0Z_1 ));
    InMux I__3929 (
            .O(N__36712),
            .I(N__36706));
    InMux I__3928 (
            .O(N__36711),
            .I(N__36706));
    LocalMux I__3927 (
            .O(N__36706),
            .I(\pid_alt.pid_preregZ0Z_1 ));
    InMux I__3926 (
            .O(N__36703),
            .I(\pid_alt.un1_pid_prereg_0_cry_0 ));
    CascadeMux I__3925 (
            .O(N__36700),
            .I(\pid_alt.source_pid_1_sqmuxa_0_a2_1_4_cascade_ ));
    InMux I__3924 (
            .O(N__36697),
            .I(N__36693));
    InMux I__3923 (
            .O(N__36696),
            .I(N__36689));
    LocalMux I__3922 (
            .O(N__36693),
            .I(N__36686));
    InMux I__3921 (
            .O(N__36692),
            .I(N__36683));
    LocalMux I__3920 (
            .O(N__36689),
            .I(throttle_order_11));
    Odrv4 I__3919 (
            .O(N__36686),
            .I(throttle_order_11));
    LocalMux I__3918 (
            .O(N__36683),
            .I(throttle_order_11));
    CascadeMux I__3917 (
            .O(N__36676),
            .I(N__36672));
    InMux I__3916 (
            .O(N__36675),
            .I(N__36668));
    InMux I__3915 (
            .O(N__36672),
            .I(N__36665));
    InMux I__3914 (
            .O(N__36671),
            .I(N__36662));
    LocalMux I__3913 (
            .O(N__36668),
            .I(N__36659));
    LocalMux I__3912 (
            .O(N__36665),
            .I(N__36656));
    LocalMux I__3911 (
            .O(N__36662),
            .I(throttle_order_6));
    Odrv12 I__3910 (
            .O(N__36659),
            .I(throttle_order_6));
    Odrv4 I__3909 (
            .O(N__36656),
            .I(throttle_order_6));
    CascadeMux I__3908 (
            .O(N__36649),
            .I(N__36645));
    CascadeMux I__3907 (
            .O(N__36648),
            .I(N__36639));
    InMux I__3906 (
            .O(N__36645),
            .I(N__36625));
    InMux I__3905 (
            .O(N__36644),
            .I(N__36625));
    InMux I__3904 (
            .O(N__36643),
            .I(N__36625));
    InMux I__3903 (
            .O(N__36642),
            .I(N__36625));
    InMux I__3902 (
            .O(N__36639),
            .I(N__36625));
    InMux I__3901 (
            .O(N__36638),
            .I(N__36625));
    LocalMux I__3900 (
            .O(N__36625),
            .I(\pid_alt.source_pid_9_0_tz_6 ));
    CascadeMux I__3899 (
            .O(N__36622),
            .I(\pid_alt.N_52_cascade_ ));
    InMux I__3898 (
            .O(N__36619),
            .I(\ppm_encoder_1.un1_throttle_cry_6 ));
    InMux I__3897 (
            .O(N__36616),
            .I(bfn_4_10_0_));
    InMux I__3896 (
            .O(N__36613),
            .I(\ppm_encoder_1.un1_throttle_cry_8 ));
    InMux I__3895 (
            .O(N__36610),
            .I(N__36607));
    LocalMux I__3894 (
            .O(N__36607),
            .I(N__36604));
    Odrv4 I__3893 (
            .O(N__36604),
            .I(\ppm_encoder_1.un1_throttle_cry_9_THRU_CO ));
    InMux I__3892 (
            .O(N__36601),
            .I(\ppm_encoder_1.un1_throttle_cry_9 ));
    InMux I__3891 (
            .O(N__36598),
            .I(N__36595));
    LocalMux I__3890 (
            .O(N__36595),
            .I(N__36592));
    Odrv4 I__3889 (
            .O(N__36592),
            .I(\ppm_encoder_1.un1_throttle_cry_10_THRU_CO ));
    InMux I__3888 (
            .O(N__36589),
            .I(\ppm_encoder_1.un1_throttle_cry_10 ));
    InMux I__3887 (
            .O(N__36586),
            .I(\ppm_encoder_1.un1_throttle_cry_11 ));
    InMux I__3886 (
            .O(N__36583),
            .I(N__36580));
    LocalMux I__3885 (
            .O(N__36580),
            .I(N__36577));
    Odrv4 I__3884 (
            .O(N__36577),
            .I(\ppm_encoder_1.un1_throttle_cry_12_THRU_CO ));
    InMux I__3883 (
            .O(N__36574),
            .I(\ppm_encoder_1.un1_throttle_cry_12 ));
    InMux I__3882 (
            .O(N__36571),
            .I(\ppm_encoder_1.un1_throttle_cry_13 ));
    CascadeMux I__3881 (
            .O(N__36568),
            .I(N__36564));
    InMux I__3880 (
            .O(N__36567),
            .I(N__36561));
    InMux I__3879 (
            .O(N__36564),
            .I(N__36557));
    LocalMux I__3878 (
            .O(N__36561),
            .I(N__36554));
    InMux I__3877 (
            .O(N__36560),
            .I(N__36551));
    LocalMux I__3876 (
            .O(N__36557),
            .I(throttle_order_10));
    Odrv12 I__3875 (
            .O(N__36554),
            .I(throttle_order_10));
    LocalMux I__3874 (
            .O(N__36551),
            .I(throttle_order_10));
    CascadeMux I__3873 (
            .O(N__36544),
            .I(N__36541));
    InMux I__3872 (
            .O(N__36541),
            .I(N__36537));
    InMux I__3871 (
            .O(N__36540),
            .I(N__36534));
    LocalMux I__3870 (
            .O(N__36537),
            .I(N__36531));
    LocalMux I__3869 (
            .O(N__36534),
            .I(\ppm_encoder_1.throttleZ0Z_5 ));
    Odrv12 I__3868 (
            .O(N__36531),
            .I(\ppm_encoder_1.throttleZ0Z_5 ));
    InMux I__3867 (
            .O(N__36526),
            .I(N__36523));
    LocalMux I__3866 (
            .O(N__36523),
            .I(\ppm_encoder_1.un1_throttle_cry_0_THRU_CO ));
    InMux I__3865 (
            .O(N__36520),
            .I(\ppm_encoder_1.un1_throttle_cry_0 ));
    InMux I__3864 (
            .O(N__36517),
            .I(N__36514));
    LocalMux I__3863 (
            .O(N__36514),
            .I(N__36511));
    Odrv4 I__3862 (
            .O(N__36511),
            .I(\ppm_encoder_1.un1_throttle_cry_1_THRU_CO ));
    InMux I__3861 (
            .O(N__36508),
            .I(\ppm_encoder_1.un1_throttle_cry_1 ));
    InMux I__3860 (
            .O(N__36505),
            .I(N__36502));
    LocalMux I__3859 (
            .O(N__36502),
            .I(N__36499));
    Odrv4 I__3858 (
            .O(N__36499),
            .I(\ppm_encoder_1.un1_throttle_cry_2_THRU_CO ));
    InMux I__3857 (
            .O(N__36496),
            .I(\ppm_encoder_1.un1_throttle_cry_2 ));
    InMux I__3856 (
            .O(N__36493),
            .I(N__36490));
    LocalMux I__3855 (
            .O(N__36490),
            .I(N__36487));
    Odrv4 I__3854 (
            .O(N__36487),
            .I(\ppm_encoder_1.un1_throttle_cry_3_THRU_CO ));
    InMux I__3853 (
            .O(N__36484),
            .I(\ppm_encoder_1.un1_throttle_cry_3 ));
    InMux I__3852 (
            .O(N__36481),
            .I(N__36478));
    LocalMux I__3851 (
            .O(N__36478),
            .I(\ppm_encoder_1.un1_throttle_cry_4_THRU_CO ));
    InMux I__3850 (
            .O(N__36475),
            .I(\ppm_encoder_1.un1_throttle_cry_4 ));
    CascadeMux I__3849 (
            .O(N__36472),
            .I(N__36469));
    InMux I__3848 (
            .O(N__36469),
            .I(N__36466));
    LocalMux I__3847 (
            .O(N__36466),
            .I(N__36463));
    Span4Mux_h I__3846 (
            .O(N__36463),
            .I(N__36460));
    Odrv4 I__3845 (
            .O(N__36460),
            .I(\ppm_encoder_1.un1_throttle_cry_5_THRU_CO ));
    InMux I__3844 (
            .O(N__36457),
            .I(\ppm_encoder_1.un1_throttle_cry_5 ));
    InMux I__3843 (
            .O(N__36454),
            .I(N__36451));
    LocalMux I__3842 (
            .O(N__36451),
            .I(N__36446));
    InMux I__3841 (
            .O(N__36450),
            .I(N__36443));
    InMux I__3840 (
            .O(N__36449),
            .I(N__36440));
    Span4Mux_s3_v I__3839 (
            .O(N__36446),
            .I(N__36435));
    LocalMux I__3838 (
            .O(N__36443),
            .I(N__36435));
    LocalMux I__3837 (
            .O(N__36440),
            .I(\ppm_encoder_1.throttleZ0Z_2 ));
    Odrv4 I__3836 (
            .O(N__36435),
            .I(\ppm_encoder_1.throttleZ0Z_2 ));
    InMux I__3835 (
            .O(N__36430),
            .I(N__36426));
    InMux I__3834 (
            .O(N__36429),
            .I(N__36423));
    LocalMux I__3833 (
            .O(N__36426),
            .I(N__36420));
    LocalMux I__3832 (
            .O(N__36423),
            .I(\ppm_encoder_1.aileronZ0Z_5 ));
    Odrv12 I__3831 (
            .O(N__36420),
            .I(\ppm_encoder_1.aileronZ0Z_5 ));
    CascadeMux I__3830 (
            .O(N__36415),
            .I(N__36411));
    InMux I__3829 (
            .O(N__36414),
            .I(N__36405));
    InMux I__3828 (
            .O(N__36411),
            .I(N__36405));
    CascadeMux I__3827 (
            .O(N__36410),
            .I(N__36402));
    LocalMux I__3826 (
            .O(N__36405),
            .I(N__36399));
    InMux I__3825 (
            .O(N__36402),
            .I(N__36396));
    Span4Mux_h I__3824 (
            .O(N__36399),
            .I(N__36393));
    LocalMux I__3823 (
            .O(N__36396),
            .I(\ppm_encoder_1.throttleZ0Z_1 ));
    Odrv4 I__3822 (
            .O(N__36393),
            .I(\ppm_encoder_1.throttleZ0Z_1 ));
    CascadeMux I__3821 (
            .O(N__36388),
            .I(\ppm_encoder_1.N_264_i_i_cascade_ ));
    CascadeMux I__3820 (
            .O(N__36385),
            .I(\ppm_encoder_1.N_465_cascade_ ));
    CascadeMux I__3819 (
            .O(N__36382),
            .I(\ppm_encoder_1.un2_throttle_iv_0_2_8_cascade_ ));
    InMux I__3818 (
            .O(N__36379),
            .I(N__36376));
    LocalMux I__3817 (
            .O(N__36376),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_8 ));
    CascadeMux I__3816 (
            .O(N__36373),
            .I(N__36370));
    InMux I__3815 (
            .O(N__36370),
            .I(N__36367));
    LocalMux I__3814 (
            .O(N__36367),
            .I(N__36364));
    Odrv4 I__3813 (
            .O(N__36364),
            .I(\ppm_encoder_1.rudderZ0Z_5 ));
    CascadeMux I__3812 (
            .O(N__36361),
            .I(\ppm_encoder_1.N_507_cascade_ ));
    CascadeMux I__3811 (
            .O(N__36358),
            .I(\ppm_encoder_1.un2_throttle_iv_0_1_2_cascade_ ));
    CascadeMux I__3810 (
            .O(N__36355),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_2_cascade_ ));
    InMux I__3809 (
            .O(N__36352),
            .I(N__36349));
    LocalMux I__3808 (
            .O(N__36349),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_5 ));
    CascadeMux I__3807 (
            .O(N__36346),
            .I(\ppm_encoder_1.N_513_cascade_ ));
    InMux I__3806 (
            .O(N__36343),
            .I(N__36340));
    LocalMux I__3805 (
            .O(N__36340),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_2 ));
    CascadeMux I__3804 (
            .O(N__36337),
            .I(\ppm_encoder_1.un2_throttle_0_0_2_5_cascade_ ));
    InMux I__3803 (
            .O(N__36334),
            .I(N__36331));
    LocalMux I__3802 (
            .O(N__36331),
            .I(\ppm_encoder_1.un2_throttle_iv_0_0_5 ));
    InMux I__3801 (
            .O(N__36328),
            .I(N__36325));
    LocalMux I__3800 (
            .O(N__36325),
            .I(N__36322));
    Odrv4 I__3799 (
            .O(N__36322),
            .I(\ppm_encoder_1.pulses2count_9_0_1_1 ));
    InMux I__3798 (
            .O(N__36319),
            .I(N__36316));
    LocalMux I__3797 (
            .O(N__36316),
            .I(N__36313));
    Span4Mux_s3_h I__3796 (
            .O(N__36313),
            .I(N__36310));
    Odrv4 I__3795 (
            .O(N__36310),
            .I(alt_kp_5));
    InMux I__3794 (
            .O(N__36307),
            .I(N__36304));
    LocalMux I__3793 (
            .O(N__36304),
            .I(N__36301));
    Span4Mux_s3_h I__3792 (
            .O(N__36301),
            .I(N__36298));
    Odrv4 I__3791 (
            .O(N__36298),
            .I(alt_kp_7));
    InMux I__3790 (
            .O(N__36295),
            .I(N__36292));
    LocalMux I__3789 (
            .O(N__36292),
            .I(N__36289));
    Span4Mux_h I__3788 (
            .O(N__36289),
            .I(N__36286));
    Odrv4 I__3787 (
            .O(N__36286),
            .I(alt_kp_0));
    CascadeMux I__3786 (
            .O(N__36283),
            .I(\ppm_encoder_1.pulses2count_9_i_3_1_2_cascade_ ));
    InMux I__3785 (
            .O(N__36280),
            .I(N__36277));
    LocalMux I__3784 (
            .O(N__36277),
            .I(\ppm_encoder_1.pulses2count_9_0_0_1 ));
    CascadeMux I__3783 (
            .O(N__36274),
            .I(\pid_alt.N_9_0_cascade_ ));
    InMux I__3782 (
            .O(N__36271),
            .I(N__36268));
    LocalMux I__3781 (
            .O(N__36268),
            .I(\pid_alt.m21_e_10 ));
    InMux I__3780 (
            .O(N__36265),
            .I(N__36262));
    LocalMux I__3779 (
            .O(N__36262),
            .I(N__36259));
    Span4Mux_v I__3778 (
            .O(N__36259),
            .I(N__36256));
    Odrv4 I__3777 (
            .O(N__36256),
            .I(\pid_alt.error_i_acumm_preregZ0Z_18 ));
    CascadeMux I__3776 (
            .O(N__36253),
            .I(N__36250));
    InMux I__3775 (
            .O(N__36250),
            .I(N__36247));
    LocalMux I__3774 (
            .O(N__36247),
            .I(N__36244));
    Span4Mux_v I__3773 (
            .O(N__36244),
            .I(N__36241));
    Odrv4 I__3772 (
            .O(N__36241),
            .I(\pid_alt.error_i_acumm_preregZ0Z_16 ));
    InMux I__3771 (
            .O(N__36238),
            .I(N__36232));
    InMux I__3770 (
            .O(N__36237),
            .I(N__36232));
    LocalMux I__3769 (
            .O(N__36232),
            .I(\pid_alt.m7_e_4 ));
    InMux I__3768 (
            .O(N__36229),
            .I(N__36226));
    LocalMux I__3767 (
            .O(N__36226),
            .I(N__36221));
    InMux I__3766 (
            .O(N__36225),
            .I(N__36216));
    InMux I__3765 (
            .O(N__36224),
            .I(N__36216));
    Span4Mux_v I__3764 (
            .O(N__36221),
            .I(N__36213));
    LocalMux I__3763 (
            .O(N__36216),
            .I(N__36210));
    Odrv4 I__3762 (
            .O(N__36213),
            .I(\pid_alt.error_i_acumm_esr_RNI33H91Z0Z_4 ));
    Odrv4 I__3761 (
            .O(N__36210),
            .I(\pid_alt.error_i_acumm_esr_RNI33H91Z0Z_4 ));
    InMux I__3760 (
            .O(N__36205),
            .I(N__36202));
    LocalMux I__3759 (
            .O(N__36202),
            .I(N__36199));
    Span4Mux_v I__3758 (
            .O(N__36199),
            .I(N__36194));
    InMux I__3757 (
            .O(N__36198),
            .I(N__36189));
    InMux I__3756 (
            .O(N__36197),
            .I(N__36189));
    Odrv4 I__3755 (
            .O(N__36194),
            .I(\pid_alt.error_i_reg_esr_RNI7ENJZ0Z_17 ));
    LocalMux I__3754 (
            .O(N__36189),
            .I(\pid_alt.error_i_reg_esr_RNI7ENJZ0Z_17 ));
    CascadeMux I__3753 (
            .O(N__36184),
            .I(N__36181));
    InMux I__3752 (
            .O(N__36181),
            .I(N__36175));
    InMux I__3751 (
            .O(N__36180),
            .I(N__36175));
    LocalMux I__3750 (
            .O(N__36175),
            .I(\pid_alt.error_i_acumm_preregZ0Z_17 ));
    InMux I__3749 (
            .O(N__36172),
            .I(N__36169));
    LocalMux I__3748 (
            .O(N__36169),
            .I(N__36166));
    Span4Mux_v I__3747 (
            .O(N__36166),
            .I(N__36161));
    InMux I__3746 (
            .O(N__36165),
            .I(N__36156));
    InMux I__3745 (
            .O(N__36164),
            .I(N__36156));
    Odrv4 I__3744 (
            .O(N__36161),
            .I(\pid_alt.error_i_reg_esr_RNI38LJZ0Z_15 ));
    LocalMux I__3743 (
            .O(N__36156),
            .I(\pid_alt.error_i_reg_esr_RNI38LJZ0Z_15 ));
    InMux I__3742 (
            .O(N__36151),
            .I(N__36145));
    InMux I__3741 (
            .O(N__36150),
            .I(N__36145));
    LocalMux I__3740 (
            .O(N__36145),
            .I(\pid_alt.error_i_acumm_preregZ0Z_15 ));
    InMux I__3739 (
            .O(N__36142),
            .I(N__36139));
    LocalMux I__3738 (
            .O(N__36139),
            .I(N__36134));
    InMux I__3737 (
            .O(N__36138),
            .I(N__36129));
    InMux I__3736 (
            .O(N__36137),
            .I(N__36129));
    Odrv4 I__3735 (
            .O(N__36134),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ ));
    LocalMux I__3734 (
            .O(N__36129),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ ));
    InMux I__3733 (
            .O(N__36124),
            .I(N__36121));
    LocalMux I__3732 (
            .O(N__36121),
            .I(\pid_alt.error_i_acumm_preregZ0Z_20 ));
    InMux I__3731 (
            .O(N__36118),
            .I(N__36115));
    LocalMux I__3730 (
            .O(N__36115),
            .I(N__36110));
    InMux I__3729 (
            .O(N__36114),
            .I(N__36105));
    InMux I__3728 (
            .O(N__36113),
            .I(N__36105));
    Span4Mux_v I__3727 (
            .O(N__36110),
            .I(N__36100));
    LocalMux I__3726 (
            .O(N__36105),
            .I(N__36100));
    Odrv4 I__3725 (
            .O(N__36100),
            .I(\pid_alt.error_i_acumm_esr_RNIJ6LMZ0Z_13 ));
    InMux I__3724 (
            .O(N__36097),
            .I(N__36092));
    InMux I__3723 (
            .O(N__36096),
            .I(N__36087));
    InMux I__3722 (
            .O(N__36095),
            .I(N__36087));
    LocalMux I__3721 (
            .O(N__36092),
            .I(\pid_alt.error_i_acumm_preregZ0Z_10 ));
    LocalMux I__3720 (
            .O(N__36087),
            .I(\pid_alt.error_i_acumm_preregZ0Z_10 ));
    CascadeMux I__3719 (
            .O(N__36082),
            .I(\pid_alt.m21_e_2_cascade_ ));
    InMux I__3718 (
            .O(N__36079),
            .I(N__36076));
    LocalMux I__3717 (
            .O(N__36076),
            .I(N__36072));
    InMux I__3716 (
            .O(N__36075),
            .I(N__36069));
    Odrv4 I__3715 (
            .O(N__36072),
            .I(\pid_alt.error_i_acumm_preregZ0Z_2 ));
    LocalMux I__3714 (
            .O(N__36069),
            .I(\pid_alt.error_i_acumm_preregZ0Z_2 ));
    CascadeMux I__3713 (
            .O(N__36064),
            .I(N__36061));
    InMux I__3712 (
            .O(N__36061),
            .I(N__36057));
    InMux I__3711 (
            .O(N__36060),
            .I(N__36054));
    LocalMux I__3710 (
            .O(N__36057),
            .I(\pid_alt.error_i_acumm_preregZ0Z_3 ));
    LocalMux I__3709 (
            .O(N__36054),
            .I(\pid_alt.error_i_acumm_preregZ0Z_3 ));
    CascadeMux I__3708 (
            .O(N__36049),
            .I(N__36046));
    InMux I__3707 (
            .O(N__36046),
            .I(N__36041));
    InMux I__3706 (
            .O(N__36045),
            .I(N__36038));
    InMux I__3705 (
            .O(N__36044),
            .I(N__36035));
    LocalMux I__3704 (
            .O(N__36041),
            .I(\pid_alt.m35_e_3 ));
    LocalMux I__3703 (
            .O(N__36038),
            .I(\pid_alt.m35_e_3 ));
    LocalMux I__3702 (
            .O(N__36035),
            .I(\pid_alt.m35_e_3 ));
    CascadeMux I__3701 (
            .O(N__36028),
            .I(N__36022));
    InMux I__3700 (
            .O(N__36027),
            .I(N__36017));
    InMux I__3699 (
            .O(N__36026),
            .I(N__36014));
    InMux I__3698 (
            .O(N__36025),
            .I(N__36005));
    InMux I__3697 (
            .O(N__36022),
            .I(N__36005));
    InMux I__3696 (
            .O(N__36021),
            .I(N__36005));
    InMux I__3695 (
            .O(N__36020),
            .I(N__36005));
    LocalMux I__3694 (
            .O(N__36017),
            .I(\pid_alt.N_62_mux ));
    LocalMux I__3693 (
            .O(N__36014),
            .I(\pid_alt.N_62_mux ));
    LocalMux I__3692 (
            .O(N__36005),
            .I(\pid_alt.N_62_mux ));
    CascadeMux I__3691 (
            .O(N__35998),
            .I(\pid_alt.N_545_cascade_ ));
    InMux I__3690 (
            .O(N__35995),
            .I(N__35990));
    InMux I__3689 (
            .O(N__35994),
            .I(N__35987));
    InMux I__3688 (
            .O(N__35993),
            .I(N__35984));
    LocalMux I__3687 (
            .O(N__35990),
            .I(\pid_alt.error_i_acumm7lto12 ));
    LocalMux I__3686 (
            .O(N__35987),
            .I(\pid_alt.error_i_acumm7lto12 ));
    LocalMux I__3685 (
            .O(N__35984),
            .I(\pid_alt.error_i_acumm7lto12 ));
    CascadeMux I__3684 (
            .O(N__35977),
            .I(N__35970));
    CascadeMux I__3683 (
            .O(N__35976),
            .I(N__35966));
    CascadeMux I__3682 (
            .O(N__35975),
            .I(N__35962));
    InMux I__3681 (
            .O(N__35974),
            .I(N__35957));
    InMux I__3680 (
            .O(N__35973),
            .I(N__35944));
    InMux I__3679 (
            .O(N__35970),
            .I(N__35944));
    InMux I__3678 (
            .O(N__35969),
            .I(N__35944));
    InMux I__3677 (
            .O(N__35966),
            .I(N__35944));
    InMux I__3676 (
            .O(N__35965),
            .I(N__35944));
    InMux I__3675 (
            .O(N__35962),
            .I(N__35944));
    InMux I__3674 (
            .O(N__35961),
            .I(N__35941));
    InMux I__3673 (
            .O(N__35960),
            .I(N__35938));
    LocalMux I__3672 (
            .O(N__35957),
            .I(\pid_alt.N_158 ));
    LocalMux I__3671 (
            .O(N__35944),
            .I(\pid_alt.N_158 ));
    LocalMux I__3670 (
            .O(N__35941),
            .I(\pid_alt.N_158 ));
    LocalMux I__3669 (
            .O(N__35938),
            .I(\pid_alt.N_158 ));
    CascadeMux I__3668 (
            .O(N__35929),
            .I(\pid_alt.error_i_acumm_prereg_esr_RNIFJA3Z0Z_14_cascade_ ));
    CascadeMux I__3667 (
            .O(N__35926),
            .I(N__35923));
    InMux I__3666 (
            .O(N__35923),
            .I(N__35917));
    InMux I__3665 (
            .O(N__35922),
            .I(N__35914));
    InMux I__3664 (
            .O(N__35921),
            .I(N__35909));
    InMux I__3663 (
            .O(N__35920),
            .I(N__35909));
    LocalMux I__3662 (
            .O(N__35917),
            .I(\pid_alt.N_9_0 ));
    LocalMux I__3661 (
            .O(N__35914),
            .I(\pid_alt.N_9_0 ));
    LocalMux I__3660 (
            .O(N__35909),
            .I(\pid_alt.N_9_0 ));
    InMux I__3659 (
            .O(N__35902),
            .I(N__35898));
    InMux I__3658 (
            .O(N__35901),
            .I(N__35895));
    LocalMux I__3657 (
            .O(N__35898),
            .I(N__35892));
    LocalMux I__3656 (
            .O(N__35895),
            .I(N__35889));
    Span4Mux_h I__3655 (
            .O(N__35892),
            .I(N__35884));
    Span4Mux_v I__3654 (
            .O(N__35889),
            .I(N__35884));
    Span4Mux_v I__3653 (
            .O(N__35884),
            .I(N__35881));
    Span4Mux_s3_h I__3652 (
            .O(N__35881),
            .I(N__35878));
    Span4Mux_h I__3651 (
            .O(N__35878),
            .I(N__35875));
    Odrv4 I__3650 (
            .O(N__35875),
            .I(\pid_alt.error_p_regZ0Z_19 ));
    CascadeMux I__3649 (
            .O(N__35872),
            .I(\pid_alt.error_d_reg_prev_esr_RNI86IMZ0Z_19_cascade_ ));
    InMux I__3648 (
            .O(N__35869),
            .I(N__35866));
    LocalMux I__3647 (
            .O(N__35866),
            .I(\pid_alt.error_d_reg_prev_esr_RNI86IMZ0Z_19 ));
    CascadeMux I__3646 (
            .O(N__35863),
            .I(N__35860));
    InMux I__3645 (
            .O(N__35860),
            .I(N__35854));
    InMux I__3644 (
            .O(N__35859),
            .I(N__35854));
    LocalMux I__3643 (
            .O(N__35854),
            .I(\pid_alt.un1_pid_prereg_236_1 ));
    InMux I__3642 (
            .O(N__35851),
            .I(N__35844));
    InMux I__3641 (
            .O(N__35850),
            .I(N__35844));
    InMux I__3640 (
            .O(N__35849),
            .I(N__35841));
    LocalMux I__3639 (
            .O(N__35844),
            .I(N__35836));
    LocalMux I__3638 (
            .O(N__35841),
            .I(N__35836));
    Span12Mux_v I__3637 (
            .O(N__35836),
            .I(N__35833));
    Odrv12 I__3636 (
            .O(N__35833),
            .I(\pid_alt.error_d_regZ0Z_19 ));
    InMux I__3635 (
            .O(N__35830),
            .I(N__35826));
    InMux I__3634 (
            .O(N__35829),
            .I(N__35823));
    LocalMux I__3633 (
            .O(N__35826),
            .I(\pid_alt.error_d_reg_prevZ0Z_19 ));
    LocalMux I__3632 (
            .O(N__35823),
            .I(\pid_alt.error_d_reg_prevZ0Z_19 ));
    InMux I__3631 (
            .O(N__35818),
            .I(N__35809));
    InMux I__3630 (
            .O(N__35817),
            .I(N__35809));
    InMux I__3629 (
            .O(N__35816),
            .I(N__35809));
    LocalMux I__3628 (
            .O(N__35809),
            .I(N__35805));
    InMux I__3627 (
            .O(N__35808),
            .I(N__35801));
    Span4Mux_s2_h I__3626 (
            .O(N__35805),
            .I(N__35797));
    InMux I__3625 (
            .O(N__35804),
            .I(N__35794));
    LocalMux I__3624 (
            .O(N__35801),
            .I(N__35791));
    InMux I__3623 (
            .O(N__35800),
            .I(N__35788));
    Odrv4 I__3622 (
            .O(N__35797),
            .I(\pid_alt.error_d_reg_prevZ0Z_20 ));
    LocalMux I__3621 (
            .O(N__35794),
            .I(\pid_alt.error_d_reg_prevZ0Z_20 ));
    Odrv4 I__3620 (
            .O(N__35791),
            .I(\pid_alt.error_d_reg_prevZ0Z_20 ));
    LocalMux I__3619 (
            .O(N__35788),
            .I(\pid_alt.error_d_reg_prevZ0Z_20 ));
    InMux I__3618 (
            .O(N__35779),
            .I(N__35769));
    InMux I__3617 (
            .O(N__35778),
            .I(N__35769));
    InMux I__3616 (
            .O(N__35777),
            .I(N__35769));
    InMux I__3615 (
            .O(N__35776),
            .I(N__35766));
    LocalMux I__3614 (
            .O(N__35769),
            .I(N__35758));
    LocalMux I__3613 (
            .O(N__35766),
            .I(N__35758));
    InMux I__3612 (
            .O(N__35765),
            .I(N__35751));
    InMux I__3611 (
            .O(N__35764),
            .I(N__35751));
    InMux I__3610 (
            .O(N__35763),
            .I(N__35751));
    Sp12to4 I__3609 (
            .O(N__35758),
            .I(N__35746));
    LocalMux I__3608 (
            .O(N__35751),
            .I(N__35746));
    Span12Mux_s7_h I__3607 (
            .O(N__35746),
            .I(N__35743));
    Span12Mux_v I__3606 (
            .O(N__35743),
            .I(N__35740));
    Odrv12 I__3605 (
            .O(N__35740),
            .I(\pid_alt.error_d_regZ0Z_20 ));
    CascadeMux I__3604 (
            .O(N__35737),
            .I(N__35730));
    CascadeMux I__3603 (
            .O(N__35736),
            .I(N__35726));
    CascadeMux I__3602 (
            .O(N__35735),
            .I(N__35723));
    CascadeMux I__3601 (
            .O(N__35734),
            .I(N__35720));
    CascadeMux I__3600 (
            .O(N__35733),
            .I(N__35717));
    InMux I__3599 (
            .O(N__35730),
            .I(N__35712));
    InMux I__3598 (
            .O(N__35729),
            .I(N__35712));
    InMux I__3597 (
            .O(N__35726),
            .I(N__35705));
    InMux I__3596 (
            .O(N__35723),
            .I(N__35705));
    InMux I__3595 (
            .O(N__35720),
            .I(N__35705));
    InMux I__3594 (
            .O(N__35717),
            .I(N__35702));
    LocalMux I__3593 (
            .O(N__35712),
            .I(N__35699));
    LocalMux I__3592 (
            .O(N__35705),
            .I(\pid_alt.error_p_regZ0Z_20 ));
    LocalMux I__3591 (
            .O(N__35702),
            .I(\pid_alt.error_p_regZ0Z_20 ));
    Odrv12 I__3590 (
            .O(N__35699),
            .I(\pid_alt.error_p_regZ0Z_20 ));
    InMux I__3589 (
            .O(N__35692),
            .I(N__35689));
    LocalMux I__3588 (
            .O(N__35689),
            .I(N__35681));
    InMux I__3587 (
            .O(N__35688),
            .I(N__35674));
    InMux I__3586 (
            .O(N__35687),
            .I(N__35674));
    InMux I__3585 (
            .O(N__35686),
            .I(N__35674));
    InMux I__3584 (
            .O(N__35685),
            .I(N__35671));
    InMux I__3583 (
            .O(N__35684),
            .I(N__35668));
    Odrv4 I__3582 (
            .O(N__35681),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_20_c_RNISVKK ));
    LocalMux I__3581 (
            .O(N__35674),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_20_c_RNISVKK ));
    LocalMux I__3580 (
            .O(N__35671),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_20_c_RNISVKK ));
    LocalMux I__3579 (
            .O(N__35668),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_20_c_RNISVKK ));
    InMux I__3578 (
            .O(N__35659),
            .I(N__35656));
    LocalMux I__3577 (
            .O(N__35656),
            .I(N__35651));
    InMux I__3576 (
            .O(N__35655),
            .I(N__35646));
    InMux I__3575 (
            .O(N__35654),
            .I(N__35646));
    Odrv4 I__3574 (
            .O(N__35651),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_9_c_RNIQN3F ));
    LocalMux I__3573 (
            .O(N__35646),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_9_c_RNIQN3F ));
    InMux I__3572 (
            .O(N__35641),
            .I(N__35636));
    InMux I__3571 (
            .O(N__35640),
            .I(N__35631));
    InMux I__3570 (
            .O(N__35639),
            .I(N__35631));
    LocalMux I__3569 (
            .O(N__35636),
            .I(N__35628));
    LocalMux I__3568 (
            .O(N__35631),
            .I(N__35625));
    Odrv4 I__3567 (
            .O(N__35628),
            .I(\pid_alt.error_i_reg_esr_RNI7RNPZ0Z_12 ));
    Odrv4 I__3566 (
            .O(N__35625),
            .I(\pid_alt.error_i_reg_esr_RNI7RNPZ0Z_12 ));
    InMux I__3565 (
            .O(N__35620),
            .I(N__35614));
    InMux I__3564 (
            .O(N__35619),
            .I(N__35614));
    LocalMux I__3563 (
            .O(N__35614),
            .I(N__35611));
    Span4Mux_h I__3562 (
            .O(N__35611),
            .I(N__35608));
    Odrv4 I__3561 (
            .O(N__35608),
            .I(\pid_alt.error_d_reg_prev_esr_RNIMJHMZ0Z_13 ));
    InMux I__3560 (
            .O(N__35605),
            .I(N__35602));
    LocalMux I__3559 (
            .O(N__35602),
            .I(\pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14 ));
    CascadeMux I__3558 (
            .O(N__35599),
            .I(\pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18_cascade_ ));
    InMux I__3557 (
            .O(N__35596),
            .I(N__35593));
    LocalMux I__3556 (
            .O(N__35593),
            .I(\pid_alt.error_d_reg_prev_esr_RNI86IM_0Z0Z_19 ));
    CascadeMux I__3555 (
            .O(N__35590),
            .I(\pid_alt.error_d_reg_prev_esr_RNI86IM_0Z0Z_19_cascade_ ));
    InMux I__3554 (
            .O(N__35587),
            .I(N__35584));
    LocalMux I__3553 (
            .O(N__35584),
            .I(\pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18 ));
    InMux I__3552 (
            .O(N__35581),
            .I(N__35574));
    InMux I__3551 (
            .O(N__35580),
            .I(N__35574));
    InMux I__3550 (
            .O(N__35579),
            .I(N__35571));
    LocalMux I__3549 (
            .O(N__35574),
            .I(N__35568));
    LocalMux I__3548 (
            .O(N__35571),
            .I(N__35565));
    Span12Mux_s4_h I__3547 (
            .O(N__35568),
            .I(N__35562));
    Span4Mux_v I__3546 (
            .O(N__35565),
            .I(N__35559));
    Span12Mux_v I__3545 (
            .O(N__35562),
            .I(N__35556));
    Odrv4 I__3544 (
            .O(N__35559),
            .I(\pid_alt.error_d_regZ0Z_18 ));
    Odrv12 I__3543 (
            .O(N__35556),
            .I(\pid_alt.error_d_regZ0Z_18 ));
    CascadeMux I__3542 (
            .O(N__35551),
            .I(N__35548));
    InMux I__3541 (
            .O(N__35548),
            .I(N__35542));
    InMux I__3540 (
            .O(N__35547),
            .I(N__35542));
    LocalMux I__3539 (
            .O(N__35542),
            .I(N__35539));
    Span4Mux_v I__3538 (
            .O(N__35539),
            .I(N__35536));
    Span4Mux_h I__3537 (
            .O(N__35536),
            .I(N__35533));
    Span4Mux_v I__3536 (
            .O(N__35533),
            .I(N__35530));
    Odrv4 I__3535 (
            .O(N__35530),
            .I(\pid_alt.error_p_regZ0Z_18 ));
    InMux I__3534 (
            .O(N__35527),
            .I(N__35521));
    InMux I__3533 (
            .O(N__35526),
            .I(N__35521));
    LocalMux I__3532 (
            .O(N__35521),
            .I(N__35518));
    Span4Mux_v I__3531 (
            .O(N__35518),
            .I(N__35515));
    Odrv4 I__3530 (
            .O(N__35515),
            .I(\pid_alt.error_d_reg_prevZ0Z_18 ));
    CascadeMux I__3529 (
            .O(N__35512),
            .I(N__35509));
    InMux I__3528 (
            .O(N__35509),
            .I(N__35506));
    LocalMux I__3527 (
            .O(N__35506),
            .I(\pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18 ));
    InMux I__3526 (
            .O(N__35503),
            .I(N__35497));
    InMux I__3525 (
            .O(N__35502),
            .I(N__35497));
    LocalMux I__3524 (
            .O(N__35497),
            .I(N__35494));
    Span4Mux_h I__3523 (
            .O(N__35494),
            .I(N__35491));
    Span4Mux_v I__3522 (
            .O(N__35491),
            .I(N__35488));
    Odrv4 I__3521 (
            .O(N__35488),
            .I(\pid_alt.error_d_reg_prev_esr_RNI20IMZ0Z_17 ));
    CascadeMux I__3520 (
            .O(N__35485),
            .I(\pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18_cascade_ ));
    InMux I__3519 (
            .O(N__35482),
            .I(N__35479));
    LocalMux I__3518 (
            .O(N__35479),
            .I(N__35474));
    InMux I__3517 (
            .O(N__35478),
            .I(N__35469));
    InMux I__3516 (
            .O(N__35477),
            .I(N__35469));
    Odrv4 I__3515 (
            .O(N__35474),
            .I(\pid_alt.error_i_reg_esr_RNI9HOJZ0Z_18 ));
    LocalMux I__3514 (
            .O(N__35469),
            .I(\pid_alt.error_i_reg_esr_RNI9HOJZ0Z_18 ));
    InMux I__3513 (
            .O(N__35464),
            .I(N__35458));
    InMux I__3512 (
            .O(N__35463),
            .I(N__35458));
    LocalMux I__3511 (
            .O(N__35458),
            .I(\pid_alt.error_d_reg_prevZ0Z_12 ));
    InMux I__3510 (
            .O(N__35455),
            .I(N__35449));
    InMux I__3509 (
            .O(N__35454),
            .I(N__35449));
    LocalMux I__3508 (
            .O(N__35449),
            .I(N__35446));
    Span4Mux_h I__3507 (
            .O(N__35446),
            .I(N__35443));
    Span4Mux_v I__3506 (
            .O(N__35443),
            .I(N__35440));
    Odrv4 I__3505 (
            .O(N__35440),
            .I(\pid_alt.error_p_regZ0Z_12 ));
    InMux I__3504 (
            .O(N__35437),
            .I(N__35430));
    InMux I__3503 (
            .O(N__35436),
            .I(N__35430));
    InMux I__3502 (
            .O(N__35435),
            .I(N__35427));
    LocalMux I__3501 (
            .O(N__35430),
            .I(N__35422));
    LocalMux I__3500 (
            .O(N__35427),
            .I(N__35422));
    Span12Mux_v I__3499 (
            .O(N__35422),
            .I(N__35419));
    Odrv12 I__3498 (
            .O(N__35419),
            .I(\pid_alt.error_d_regZ0Z_12 ));
    InMux I__3497 (
            .O(N__35416),
            .I(N__35413));
    LocalMux I__3496 (
            .O(N__35413),
            .I(\pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12 ));
    InMux I__3495 (
            .O(N__35410),
            .I(N__35404));
    InMux I__3494 (
            .O(N__35409),
            .I(N__35404));
    LocalMux I__3493 (
            .O(N__35404),
            .I(N__35401));
    Span4Mux_h I__3492 (
            .O(N__35401),
            .I(N__35398));
    Odrv4 I__3491 (
            .O(N__35398),
            .I(\pid_alt.error_d_reg_prev_esr_RNIGDHMZ0Z_11 ));
    CascadeMux I__3490 (
            .O(N__35395),
            .I(\pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12_cascade_ ));
    InMux I__3489 (
            .O(N__35392),
            .I(N__35389));
    LocalMux I__3488 (
            .O(N__35389),
            .I(\pid_alt.error_d_reg_prev_esr_RNISPHM_0Z0Z_15 ));
    CascadeMux I__3487 (
            .O(N__35386),
            .I(\pid_alt.error_d_reg_prev_esr_RNISPHM_0Z0Z_15_cascade_ ));
    InMux I__3486 (
            .O(N__35383),
            .I(N__35377));
    InMux I__3485 (
            .O(N__35382),
            .I(N__35377));
    LocalMux I__3484 (
            .O(N__35377),
            .I(\pid_alt.error_d_reg_prev_esr_RNIPMHMZ0Z_14 ));
    InMux I__3483 (
            .O(N__35374),
            .I(N__35368));
    InMux I__3482 (
            .O(N__35373),
            .I(N__35368));
    LocalMux I__3481 (
            .O(N__35368),
            .I(N__35365));
    Span12Mux_h I__3480 (
            .O(N__35365),
            .I(N__35362));
    Odrv12 I__3479 (
            .O(N__35362),
            .I(\pid_alt.error_p_regZ0Z_14 ));
    CascadeMux I__3478 (
            .O(N__35359),
            .I(\pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14_cascade_ ));
    InMux I__3477 (
            .O(N__35356),
            .I(N__35347));
    InMux I__3476 (
            .O(N__35355),
            .I(N__35347));
    InMux I__3475 (
            .O(N__35354),
            .I(N__35347));
    LocalMux I__3474 (
            .O(N__35347),
            .I(N__35344));
    Span4Mux_h I__3473 (
            .O(N__35344),
            .I(N__35341));
    Span4Mux_v I__3472 (
            .O(N__35341),
            .I(N__35338));
    Span4Mux_v I__3471 (
            .O(N__35338),
            .I(N__35335));
    Odrv4 I__3470 (
            .O(N__35335),
            .I(\pid_alt.error_d_regZ0Z_14 ));
    CascadeMux I__3469 (
            .O(N__35332),
            .I(N__35329));
    InMux I__3468 (
            .O(N__35329),
            .I(N__35323));
    InMux I__3467 (
            .O(N__35328),
            .I(N__35323));
    LocalMux I__3466 (
            .O(N__35323),
            .I(\pid_alt.error_d_reg_prevZ0Z_14 ));
    InMux I__3465 (
            .O(N__35320),
            .I(N__35314));
    InMux I__3464 (
            .O(N__35319),
            .I(N__35314));
    LocalMux I__3463 (
            .O(N__35314),
            .I(\pid_alt.error_d_reg_prevZ0Z_5 ));
    CascadeMux I__3462 (
            .O(N__35311),
            .I(N__35308));
    InMux I__3461 (
            .O(N__35308),
            .I(N__35302));
    InMux I__3460 (
            .O(N__35307),
            .I(N__35302));
    LocalMux I__3459 (
            .O(N__35302),
            .I(N__35299));
    Span4Mux_h I__3458 (
            .O(N__35299),
            .I(N__35296));
    Span4Mux_v I__3457 (
            .O(N__35296),
            .I(N__35293));
    Span4Mux_s1_h I__3456 (
            .O(N__35293),
            .I(N__35290));
    Odrv4 I__3455 (
            .O(N__35290),
            .I(\pid_alt.error_p_regZ0Z_5 ));
    InMux I__3454 (
            .O(N__35287),
            .I(N__35278));
    InMux I__3453 (
            .O(N__35286),
            .I(N__35278));
    InMux I__3452 (
            .O(N__35285),
            .I(N__35278));
    LocalMux I__3451 (
            .O(N__35278),
            .I(N__35275));
    Span4Mux_v I__3450 (
            .O(N__35275),
            .I(N__35272));
    Span4Mux_v I__3449 (
            .O(N__35272),
            .I(N__35269));
    Odrv4 I__3448 (
            .O(N__35269),
            .I(\pid_alt.error_d_regZ0Z_5 ));
    InMux I__3447 (
            .O(N__35266),
            .I(N__35263));
    LocalMux I__3446 (
            .O(N__35263),
            .I(\pid_alt.error_d_reg_prev_esr_RNI9S511_0Z0Z_5 ));
    InMux I__3445 (
            .O(N__35260),
            .I(N__35254));
    InMux I__3444 (
            .O(N__35259),
            .I(N__35254));
    LocalMux I__3443 (
            .O(N__35254),
            .I(N__35251));
    Span4Mux_h I__3442 (
            .O(N__35251),
            .I(N__35248));
    Odrv4 I__3441 (
            .O(N__35248),
            .I(\pid_alt.error_d_reg_prev_esr_RNI6P511Z0Z_4 ));
    CascadeMux I__3440 (
            .O(N__35245),
            .I(\pid_alt.error_d_reg_prev_esr_RNI9S511_0Z0Z_5_cascade_ ));
    InMux I__3439 (
            .O(N__35242),
            .I(N__35237));
    InMux I__3438 (
            .O(N__35241),
            .I(N__35234));
    InMux I__3437 (
            .O(N__35240),
            .I(N__35231));
    LocalMux I__3436 (
            .O(N__35237),
            .I(N__35226));
    LocalMux I__3435 (
            .O(N__35234),
            .I(N__35226));
    LocalMux I__3434 (
            .O(N__35231),
            .I(N__35221));
    Span12Mux_h I__3433 (
            .O(N__35226),
            .I(N__35221));
    Odrv12 I__3432 (
            .O(N__35221),
            .I(\pid_alt.error_d_regZ0Z_13 ));
    InMux I__3431 (
            .O(N__35218),
            .I(N__35214));
    InMux I__3430 (
            .O(N__35217),
            .I(N__35211));
    LocalMux I__3429 (
            .O(N__35214),
            .I(\pid_alt.error_d_reg_prevZ0Z_13 ));
    LocalMux I__3428 (
            .O(N__35211),
            .I(\pid_alt.error_d_reg_prevZ0Z_13 ));
    InMux I__3427 (
            .O(N__35206),
            .I(N__35203));
    LocalMux I__3426 (
            .O(N__35203),
            .I(N__35199));
    InMux I__3425 (
            .O(N__35202),
            .I(N__35196));
    Span4Mux_h I__3424 (
            .O(N__35199),
            .I(N__35193));
    LocalMux I__3423 (
            .O(N__35196),
            .I(N__35190));
    Span4Mux_v I__3422 (
            .O(N__35193),
            .I(N__35187));
    Odrv12 I__3421 (
            .O(N__35190),
            .I(\pid_alt.error_p_regZ0Z_13 ));
    Odrv4 I__3420 (
            .O(N__35187),
            .I(\pid_alt.error_p_regZ0Z_13 ));
    InMux I__3419 (
            .O(N__35182),
            .I(N__35179));
    LocalMux I__3418 (
            .O(N__35179),
            .I(\pid_alt.error_d_reg_prev_esr_RNIMJHM_0Z0Z_13 ));
    CascadeMux I__3417 (
            .O(N__35176),
            .I(\pid_alt.error_d_reg_prev_esr_RNIMJHM_0Z0Z_13_cascade_ ));
    InMux I__3416 (
            .O(N__35173),
            .I(N__35167));
    InMux I__3415 (
            .O(N__35172),
            .I(N__35167));
    LocalMux I__3414 (
            .O(N__35167),
            .I(\pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12 ));
    InMux I__3413 (
            .O(N__35164),
            .I(N__35160));
    InMux I__3412 (
            .O(N__35163),
            .I(N__35157));
    LocalMux I__3411 (
            .O(N__35160),
            .I(N__35154));
    LocalMux I__3410 (
            .O(N__35157),
            .I(\pid_alt.error_p_regZ0Z_4 ));
    Odrv12 I__3409 (
            .O(N__35154),
            .I(\pid_alt.error_p_regZ0Z_4 ));
    InMux I__3408 (
            .O(N__35149),
            .I(N__35145));
    InMux I__3407 (
            .O(N__35148),
            .I(N__35142));
    LocalMux I__3406 (
            .O(N__35145),
            .I(N__35139));
    LocalMux I__3405 (
            .O(N__35142),
            .I(N__35136));
    Odrv4 I__3404 (
            .O(N__35139),
            .I(\pid_alt.error_d_reg_prevZ0Z_4 ));
    Odrv4 I__3403 (
            .O(N__35136),
            .I(\pid_alt.error_d_reg_prevZ0Z_4 ));
    InMux I__3402 (
            .O(N__35131),
            .I(N__35127));
    InMux I__3401 (
            .O(N__35130),
            .I(N__35123));
    LocalMux I__3400 (
            .O(N__35127),
            .I(N__35120));
    InMux I__3399 (
            .O(N__35126),
            .I(N__35117));
    LocalMux I__3398 (
            .O(N__35123),
            .I(N__35114));
    Span4Mux_v I__3397 (
            .O(N__35120),
            .I(N__35107));
    LocalMux I__3396 (
            .O(N__35117),
            .I(N__35107));
    Span4Mux_h I__3395 (
            .O(N__35114),
            .I(N__35107));
    Span4Mux_v I__3394 (
            .O(N__35107),
            .I(N__35104));
    Span4Mux_v I__3393 (
            .O(N__35104),
            .I(N__35101));
    Odrv4 I__3392 (
            .O(N__35101),
            .I(\pid_alt.error_d_regZ0Z_4 ));
    InMux I__3391 (
            .O(N__35098),
            .I(N__35092));
    InMux I__3390 (
            .O(N__35097),
            .I(N__35092));
    LocalMux I__3389 (
            .O(N__35092),
            .I(\pid_alt.error_d_reg_prev_esr_RNI6P511_0Z0Z_4 ));
    InMux I__3388 (
            .O(N__35089),
            .I(N__35082));
    InMux I__3387 (
            .O(N__35088),
            .I(N__35082));
    InMux I__3386 (
            .O(N__35087),
            .I(N__35079));
    LocalMux I__3385 (
            .O(N__35082),
            .I(N__35076));
    LocalMux I__3384 (
            .O(N__35079),
            .I(N__35073));
    Span4Mux_h I__3383 (
            .O(N__35076),
            .I(N__35070));
    Span4Mux_v I__3382 (
            .O(N__35073),
            .I(N__35067));
    Span4Mux_v I__3381 (
            .O(N__35070),
            .I(N__35064));
    Span4Mux_v I__3380 (
            .O(N__35067),
            .I(N__35061));
    Odrv4 I__3379 (
            .O(N__35064),
            .I(\pid_alt.error_d_regZ0Z_3 ));
    Odrv4 I__3378 (
            .O(N__35061),
            .I(\pid_alt.error_d_regZ0Z_3 ));
    InMux I__3377 (
            .O(N__35056),
            .I(N__35052));
    InMux I__3376 (
            .O(N__35055),
            .I(N__35049));
    LocalMux I__3375 (
            .O(N__35052),
            .I(\pid_alt.error_d_reg_prevZ0Z_3 ));
    LocalMux I__3374 (
            .O(N__35049),
            .I(\pid_alt.error_d_reg_prevZ0Z_3 ));
    InMux I__3373 (
            .O(N__35044),
            .I(N__35038));
    InMux I__3372 (
            .O(N__35043),
            .I(N__35038));
    LocalMux I__3371 (
            .O(N__35038),
            .I(\pid_alt.error_d_reg_prev_esr_RNI3M511_0Z0Z_3 ));
    CascadeMux I__3370 (
            .O(N__35035),
            .I(N__35032));
    InMux I__3369 (
            .O(N__35032),
            .I(N__35026));
    InMux I__3368 (
            .O(N__35031),
            .I(N__35026));
    LocalMux I__3367 (
            .O(N__35026),
            .I(N__35023));
    Odrv4 I__3366 (
            .O(N__35023),
            .I(\pid_alt.error_d_reg_prev_esr_RNI0J511Z0Z_2 ));
    InMux I__3365 (
            .O(N__35020),
            .I(N__35014));
    InMux I__3364 (
            .O(N__35019),
            .I(N__35014));
    LocalMux I__3363 (
            .O(N__35014),
            .I(\pid_alt.error_d_reg_prev_esr_RNII5LS3Z0Z_1 ));
    InMux I__3362 (
            .O(N__35011),
            .I(N__35008));
    LocalMux I__3361 (
            .O(N__35008),
            .I(\pid_alt.error_d_reg_prev_esr_RNI9S511Z0Z_5 ));
    CascadeMux I__3360 (
            .O(N__35005),
            .I(\pid_alt.error_d_reg_prev_esr_RNI9S511Z0Z_5_cascade_ ));
    InMux I__3359 (
            .O(N__35002),
            .I(N__34999));
    LocalMux I__3358 (
            .O(N__34999),
            .I(N__34995));
    InMux I__3357 (
            .O(N__34998),
            .I(N__34992));
    Span4Mux_v I__3356 (
            .O(N__34995),
            .I(N__34989));
    LocalMux I__3355 (
            .O(N__34992),
            .I(N__34986));
    Span4Mux_v I__3354 (
            .O(N__34989),
            .I(N__34983));
    Span4Mux_v I__3353 (
            .O(N__34986),
            .I(N__34980));
    Span4Mux_h I__3352 (
            .O(N__34983),
            .I(N__34977));
    Odrv4 I__3351 (
            .O(N__34980),
            .I(\pid_alt.error_p_regZ0Z_6 ));
    Odrv4 I__3350 (
            .O(N__34977),
            .I(\pid_alt.error_p_regZ0Z_6 ));
    InMux I__3349 (
            .O(N__34972),
            .I(N__34968));
    InMux I__3348 (
            .O(N__34971),
            .I(N__34965));
    LocalMux I__3347 (
            .O(N__34968),
            .I(N__34962));
    LocalMux I__3346 (
            .O(N__34965),
            .I(\pid_alt.error_d_reg_prevZ0Z_6 ));
    Odrv4 I__3345 (
            .O(N__34962),
            .I(\pid_alt.error_d_reg_prevZ0Z_6 ));
    InMux I__3344 (
            .O(N__34957),
            .I(N__34951));
    InMux I__3343 (
            .O(N__34956),
            .I(N__34951));
    LocalMux I__3342 (
            .O(N__34951),
            .I(N__34948));
    Span4Mux_s3_h I__3341 (
            .O(N__34948),
            .I(N__34944));
    InMux I__3340 (
            .O(N__34947),
            .I(N__34941));
    Sp12to4 I__3339 (
            .O(N__34944),
            .I(N__34936));
    LocalMux I__3338 (
            .O(N__34941),
            .I(N__34936));
    Span12Mux_v I__3337 (
            .O(N__34936),
            .I(N__34933));
    Odrv12 I__3336 (
            .O(N__34933),
            .I(\pid_alt.error_d_regZ0Z_6 ));
    InMux I__3335 (
            .O(N__34930),
            .I(N__34924));
    InMux I__3334 (
            .O(N__34929),
            .I(N__34924));
    LocalMux I__3333 (
            .O(N__34924),
            .I(\pid_alt.error_d_reg_prev_esr_RNICV511_0Z0Z_6 ));
    InMux I__3332 (
            .O(N__34921),
            .I(N__34918));
    LocalMux I__3331 (
            .O(N__34918),
            .I(N__34915));
    Span4Mux_s3_h I__3330 (
            .O(N__34915),
            .I(N__34912));
    Odrv4 I__3329 (
            .O(N__34912),
            .I(alt_ki_0));
    InMux I__3328 (
            .O(N__34909),
            .I(N__34906));
    LocalMux I__3327 (
            .O(N__34906),
            .I(N__34903));
    Span4Mux_s3_h I__3326 (
            .O(N__34903),
            .I(N__34900));
    Odrv4 I__3325 (
            .O(N__34900),
            .I(alt_ki_1));
    InMux I__3324 (
            .O(N__34897),
            .I(N__34894));
    LocalMux I__3323 (
            .O(N__34894),
            .I(N__34891));
    Span4Mux_s3_h I__3322 (
            .O(N__34891),
            .I(N__34888));
    Odrv4 I__3321 (
            .O(N__34888),
            .I(alt_ki_2));
    InMux I__3320 (
            .O(N__34885),
            .I(N__34882));
    LocalMux I__3319 (
            .O(N__34882),
            .I(N__34879));
    Span4Mux_s3_h I__3318 (
            .O(N__34879),
            .I(N__34876));
    Odrv4 I__3317 (
            .O(N__34876),
            .I(alt_ki_3));
    InMux I__3316 (
            .O(N__34873),
            .I(N__34870));
    LocalMux I__3315 (
            .O(N__34870),
            .I(N__34867));
    Span4Mux_v I__3314 (
            .O(N__34867),
            .I(N__34864));
    Span4Mux_h I__3313 (
            .O(N__34864),
            .I(N__34861));
    Odrv4 I__3312 (
            .O(N__34861),
            .I(alt_ki_4));
    InMux I__3311 (
            .O(N__34858),
            .I(N__34855));
    LocalMux I__3310 (
            .O(N__34855),
            .I(N__34852));
    Span4Mux_v I__3309 (
            .O(N__34852),
            .I(N__34849));
    Odrv4 I__3308 (
            .O(N__34849),
            .I(alt_ki_7));
    InMux I__3307 (
            .O(N__34846),
            .I(N__34843));
    LocalMux I__3306 (
            .O(N__34843),
            .I(N__34839));
    InMux I__3305 (
            .O(N__34842),
            .I(N__34836));
    Span4Mux_h I__3304 (
            .O(N__34839),
            .I(N__34831));
    LocalMux I__3303 (
            .O(N__34836),
            .I(N__34831));
    Span4Mux_v I__3302 (
            .O(N__34831),
            .I(N__34828));
    Span4Mux_v I__3301 (
            .O(N__34828),
            .I(N__34825));
    Odrv4 I__3300 (
            .O(N__34825),
            .I(\pid_alt.error_p_regZ0Z_3 ));
    InMux I__3299 (
            .O(N__34822),
            .I(N__34819));
    LocalMux I__3298 (
            .O(N__34819),
            .I(\pid_alt.error_d_reg_prev_esr_RNI3M511Z0Z_3 ));
    CascadeMux I__3297 (
            .O(N__34816),
            .I(\pid_alt.error_d_reg_prev_esr_RNI3M511Z0Z_3_cascade_ ));
    InMux I__3296 (
            .O(N__34813),
            .I(N__34810));
    LocalMux I__3295 (
            .O(N__34810),
            .I(N__34807));
    Odrv12 I__3294 (
            .O(N__34807),
            .I(\pid_alt.error_i_acummZ0Z_4 ));
    InMux I__3293 (
            .O(N__34804),
            .I(N__34801));
    LocalMux I__3292 (
            .O(N__34801),
            .I(N__34798));
    Span4Mux_s2_h I__3291 (
            .O(N__34798),
            .I(N__34795));
    Odrv4 I__3290 (
            .O(N__34795),
            .I(alt_kp_6));
    InMux I__3289 (
            .O(N__34792),
            .I(N__34789));
    LocalMux I__3288 (
            .O(N__34789),
            .I(N__34786));
    Span4Mux_s2_h I__3287 (
            .O(N__34786),
            .I(N__34783));
    Odrv4 I__3286 (
            .O(N__34783),
            .I(alt_kp_1));
    InMux I__3285 (
            .O(N__34780),
            .I(N__34777));
    LocalMux I__3284 (
            .O(N__34777),
            .I(N__34774));
    Span4Mux_s2_h I__3283 (
            .O(N__34774),
            .I(N__34771));
    Odrv4 I__3282 (
            .O(N__34771),
            .I(alt_kp_3));
    InMux I__3281 (
            .O(N__34768),
            .I(N__34765));
    LocalMux I__3280 (
            .O(N__34765),
            .I(N__34762));
    Span4Mux_h I__3279 (
            .O(N__34762),
            .I(N__34759));
    Span4Mux_v I__3278 (
            .O(N__34759),
            .I(N__34756));
    Span4Mux_v I__3277 (
            .O(N__34756),
            .I(N__34753));
    Odrv4 I__3276 (
            .O(N__34753),
            .I(\pid_front.O_0_9 ));
    InMux I__3275 (
            .O(N__34750),
            .I(N__34747));
    LocalMux I__3274 (
            .O(N__34747),
            .I(N__34744));
    Span4Mux_h I__3273 (
            .O(N__34744),
            .I(N__34741));
    Odrv4 I__3272 (
            .O(N__34741),
            .I(\pid_alt.O_3_23 ));
    CEMux I__3271 (
            .O(N__34738),
            .I(N__34690));
    CEMux I__3270 (
            .O(N__34737),
            .I(N__34690));
    CEMux I__3269 (
            .O(N__34736),
            .I(N__34690));
    CEMux I__3268 (
            .O(N__34735),
            .I(N__34690));
    CEMux I__3267 (
            .O(N__34734),
            .I(N__34690));
    CEMux I__3266 (
            .O(N__34733),
            .I(N__34690));
    CEMux I__3265 (
            .O(N__34732),
            .I(N__34690));
    CEMux I__3264 (
            .O(N__34731),
            .I(N__34690));
    CEMux I__3263 (
            .O(N__34730),
            .I(N__34690));
    CEMux I__3262 (
            .O(N__34729),
            .I(N__34690));
    CEMux I__3261 (
            .O(N__34728),
            .I(N__34690));
    CEMux I__3260 (
            .O(N__34727),
            .I(N__34690));
    CEMux I__3259 (
            .O(N__34726),
            .I(N__34690));
    CEMux I__3258 (
            .O(N__34725),
            .I(N__34690));
    CEMux I__3257 (
            .O(N__34724),
            .I(N__34690));
    CEMux I__3256 (
            .O(N__34723),
            .I(N__34690));
    GlobalMux I__3255 (
            .O(N__34690),
            .I(N__34687));
    gio2CtrlBuf I__3254 (
            .O(N__34687),
            .I(\pid_alt.N_933_0_g ));
    CascadeMux I__3253 (
            .O(N__34684),
            .I(N__34681));
    InMux I__3252 (
            .O(N__34681),
            .I(N__34677));
    InMux I__3251 (
            .O(N__34680),
            .I(N__34674));
    LocalMux I__3250 (
            .O(N__34677),
            .I(N__34671));
    LocalMux I__3249 (
            .O(N__34674),
            .I(\pid_alt.error_i_acummZ0Z_12 ));
    Odrv4 I__3248 (
            .O(N__34671),
            .I(\pid_alt.error_i_acummZ0Z_12 ));
    InMux I__3247 (
            .O(N__34666),
            .I(N__34663));
    LocalMux I__3246 (
            .O(N__34663),
            .I(N__34659));
    InMux I__3245 (
            .O(N__34662),
            .I(N__34656));
    Span4Mux_v I__3244 (
            .O(N__34659),
            .I(N__34653));
    LocalMux I__3243 (
            .O(N__34656),
            .I(\pid_alt.error_i_acummZ0Z_5 ));
    Odrv4 I__3242 (
            .O(N__34653),
            .I(\pid_alt.error_i_acummZ0Z_5 ));
    InMux I__3241 (
            .O(N__34648),
            .I(N__34645));
    LocalMux I__3240 (
            .O(N__34645),
            .I(N__34642));
    Odrv12 I__3239 (
            .O(N__34642),
            .I(\pid_alt.error_i_acummZ0Z_3 ));
    InMux I__3238 (
            .O(N__34639),
            .I(N__34636));
    LocalMux I__3237 (
            .O(N__34636),
            .I(N__34633));
    Odrv12 I__3236 (
            .O(N__34633),
            .I(\pid_alt.error_i_acummZ0Z_1 ));
    InMux I__3235 (
            .O(N__34630),
            .I(N__34627));
    LocalMux I__3234 (
            .O(N__34627),
            .I(N__34624));
    Odrv12 I__3233 (
            .O(N__34624),
            .I(\pid_alt.error_i_acummZ0Z_2 ));
    CascadeMux I__3232 (
            .O(N__34621),
            .I(\pid_alt.error_i_acumm_prereg_esr_RNICB6L2_0Z0Z_5_cascade_ ));
    InMux I__3231 (
            .O(N__34618),
            .I(N__34615));
    LocalMux I__3230 (
            .O(N__34615),
            .I(\pid_alt.error_i_acumm_prereg_esr_RNICB6L2Z0Z_5 ));
    InMux I__3229 (
            .O(N__34612),
            .I(N__34603));
    InMux I__3228 (
            .O(N__34611),
            .I(N__34603));
    InMux I__3227 (
            .O(N__34610),
            .I(N__34603));
    LocalMux I__3226 (
            .O(N__34603),
            .I(\pid_alt.N_159 ));
    CascadeMux I__3225 (
            .O(N__34600),
            .I(\pid_alt.N_159_cascade_ ));
    InMux I__3224 (
            .O(N__34597),
            .I(N__34591));
    InMux I__3223 (
            .O(N__34596),
            .I(N__34591));
    LocalMux I__3222 (
            .O(N__34591),
            .I(N__34588));
    Span4Mux_v I__3221 (
            .O(N__34588),
            .I(N__34585));
    Span4Mux_v I__3220 (
            .O(N__34585),
            .I(N__34582));
    Odrv4 I__3219 (
            .O(N__34582),
            .I(\pid_alt.error_i_regZ0Z_20 ));
    InMux I__3218 (
            .O(N__34579),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_20 ));
    InMux I__3217 (
            .O(N__34576),
            .I(N__34573));
    LocalMux I__3216 (
            .O(N__34573),
            .I(\pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16 ));
    InMux I__3215 (
            .O(N__34570),
            .I(N__34567));
    LocalMux I__3214 (
            .O(N__34567),
            .I(N__34562));
    InMux I__3213 (
            .O(N__34566),
            .I(N__34559));
    InMux I__3212 (
            .O(N__34565),
            .I(N__34556));
    Odrv4 I__3211 (
            .O(N__34562),
            .I(\pid_alt.error_i_reg_esr_RNI5BMJZ0Z_16 ));
    LocalMux I__3210 (
            .O(N__34559),
            .I(\pid_alt.error_i_reg_esr_RNI5BMJZ0Z_16 ));
    LocalMux I__3209 (
            .O(N__34556),
            .I(\pid_alt.error_i_reg_esr_RNI5BMJZ0Z_16 ));
    InMux I__3208 (
            .O(N__34549),
            .I(N__34545));
    InMux I__3207 (
            .O(N__34548),
            .I(N__34542));
    LocalMux I__3206 (
            .O(N__34545),
            .I(N__34539));
    LocalMux I__3205 (
            .O(N__34542),
            .I(\pid_alt.error_i_acummZ0Z_10 ));
    Odrv12 I__3204 (
            .O(N__34539),
            .I(\pid_alt.error_i_acummZ0Z_10 ));
    InMux I__3203 (
            .O(N__34534),
            .I(N__34530));
    InMux I__3202 (
            .O(N__34533),
            .I(N__34527));
    LocalMux I__3201 (
            .O(N__34530),
            .I(N__34524));
    LocalMux I__3200 (
            .O(N__34527),
            .I(\pid_alt.error_i_acummZ0Z_11 ));
    Odrv4 I__3199 (
            .O(N__34524),
            .I(\pid_alt.error_i_acummZ0Z_11 ));
    InMux I__3198 (
            .O(N__34519),
            .I(N__34515));
    InMux I__3197 (
            .O(N__34518),
            .I(N__34512));
    LocalMux I__3196 (
            .O(N__34515),
            .I(N__34509));
    LocalMux I__3195 (
            .O(N__34512),
            .I(\pid_alt.error_i_acummZ0Z_6 ));
    Odrv4 I__3194 (
            .O(N__34509),
            .I(\pid_alt.error_i_acummZ0Z_6 ));
    InMux I__3193 (
            .O(N__34504),
            .I(N__34500));
    InMux I__3192 (
            .O(N__34503),
            .I(N__34497));
    LocalMux I__3191 (
            .O(N__34500),
            .I(N__34494));
    LocalMux I__3190 (
            .O(N__34497),
            .I(\pid_alt.error_i_acummZ0Z_7 ));
    Odrv12 I__3189 (
            .O(N__34494),
            .I(\pid_alt.error_i_acummZ0Z_7 ));
    InMux I__3188 (
            .O(N__34489),
            .I(N__34485));
    InMux I__3187 (
            .O(N__34488),
            .I(N__34482));
    LocalMux I__3186 (
            .O(N__34485),
            .I(N__34479));
    LocalMux I__3185 (
            .O(N__34482),
            .I(\pid_alt.error_i_acummZ0Z_8 ));
    Odrv4 I__3184 (
            .O(N__34479),
            .I(\pid_alt.error_i_acummZ0Z_8 ));
    InMux I__3183 (
            .O(N__34474),
            .I(N__34470));
    InMux I__3182 (
            .O(N__34473),
            .I(N__34467));
    LocalMux I__3181 (
            .O(N__34470),
            .I(N__34462));
    LocalMux I__3180 (
            .O(N__34467),
            .I(N__34462));
    Odrv4 I__3179 (
            .O(N__34462),
            .I(\pid_alt.error_i_acummZ0Z_9 ));
    InMux I__3178 (
            .O(N__34459),
            .I(N__34456));
    LocalMux I__3177 (
            .O(N__34456),
            .I(N__34453));
    Span4Mux_h I__3176 (
            .O(N__34453),
            .I(N__34450));
    Span4Mux_v I__3175 (
            .O(N__34450),
            .I(N__34447));
    Odrv4 I__3174 (
            .O(N__34447),
            .I(\pid_alt.error_i_regZ0Z_12 ));
    InMux I__3173 (
            .O(N__34444),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_11 ));
    CascadeMux I__3172 (
            .O(N__34441),
            .I(N__34438));
    InMux I__3171 (
            .O(N__34438),
            .I(N__34435));
    LocalMux I__3170 (
            .O(N__34435),
            .I(N__34432));
    Span4Mux_v I__3169 (
            .O(N__34432),
            .I(N__34429));
    Odrv4 I__3168 (
            .O(N__34429),
            .I(\pid_alt.error_i_regZ0Z_13 ));
    InMux I__3167 (
            .O(N__34426),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_12 ));
    InMux I__3166 (
            .O(N__34423),
            .I(N__34420));
    LocalMux I__3165 (
            .O(N__34420),
            .I(N__34417));
    Span4Mux_v I__3164 (
            .O(N__34417),
            .I(N__34414));
    Span4Mux_v I__3163 (
            .O(N__34414),
            .I(N__34411));
    Odrv4 I__3162 (
            .O(N__34411),
            .I(\pid_alt.error_i_regZ0Z_14 ));
    InMux I__3161 (
            .O(N__34408),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_13 ));
    InMux I__3160 (
            .O(N__34405),
            .I(N__34402));
    LocalMux I__3159 (
            .O(N__34402),
            .I(N__34399));
    Span4Mux_v I__3158 (
            .O(N__34399),
            .I(N__34396));
    Span4Mux_v I__3157 (
            .O(N__34396),
            .I(N__34393));
    Odrv4 I__3156 (
            .O(N__34393),
            .I(\pid_alt.error_i_regZ0Z_15 ));
    InMux I__3155 (
            .O(N__34390),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_14 ));
    InMux I__3154 (
            .O(N__34387),
            .I(N__34384));
    LocalMux I__3153 (
            .O(N__34384),
            .I(N__34381));
    Span4Mux_v I__3152 (
            .O(N__34381),
            .I(N__34378));
    Span4Mux_v I__3151 (
            .O(N__34378),
            .I(N__34375));
    Odrv4 I__3150 (
            .O(N__34375),
            .I(\pid_alt.error_i_regZ0Z_16 ));
    InMux I__3149 (
            .O(N__34372),
            .I(bfn_2_18_0_));
    InMux I__3148 (
            .O(N__34369),
            .I(N__34366));
    LocalMux I__3147 (
            .O(N__34366),
            .I(N__34363));
    Span4Mux_h I__3146 (
            .O(N__34363),
            .I(N__34360));
    Span4Mux_v I__3145 (
            .O(N__34360),
            .I(N__34357));
    Odrv4 I__3144 (
            .O(N__34357),
            .I(\pid_alt.error_i_regZ0Z_17 ));
    InMux I__3143 (
            .O(N__34354),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_16 ));
    InMux I__3142 (
            .O(N__34351),
            .I(N__34348));
    LocalMux I__3141 (
            .O(N__34348),
            .I(N__34345));
    Span4Mux_v I__3140 (
            .O(N__34345),
            .I(N__34342));
    Span4Mux_v I__3139 (
            .O(N__34342),
            .I(N__34339));
    Odrv4 I__3138 (
            .O(N__34339),
            .I(\pid_alt.error_i_regZ0Z_18 ));
    InMux I__3137 (
            .O(N__34336),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_17 ));
    InMux I__3136 (
            .O(N__34333),
            .I(N__34330));
    LocalMux I__3135 (
            .O(N__34330),
            .I(N__34327));
    Span4Mux_v I__3134 (
            .O(N__34327),
            .I(N__34324));
    Span4Mux_v I__3133 (
            .O(N__34324),
            .I(N__34321));
    Odrv4 I__3132 (
            .O(N__34321),
            .I(\pid_alt.error_i_regZ0Z_19 ));
    InMux I__3131 (
            .O(N__34318),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_18 ));
    InMux I__3130 (
            .O(N__34315),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_19 ));
    CascadeMux I__3129 (
            .O(N__34312),
            .I(N__34309));
    InMux I__3128 (
            .O(N__34309),
            .I(N__34306));
    LocalMux I__3127 (
            .O(N__34306),
            .I(\pid_alt.error_i_regZ0Z_4 ));
    InMux I__3126 (
            .O(N__34303),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_3 ));
    CascadeMux I__3125 (
            .O(N__34300),
            .I(N__34297));
    InMux I__3124 (
            .O(N__34297),
            .I(N__34294));
    LocalMux I__3123 (
            .O(N__34294),
            .I(\pid_alt.error_i_regZ0Z_5 ));
    InMux I__3122 (
            .O(N__34291),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_4 ));
    CascadeMux I__3121 (
            .O(N__34288),
            .I(N__34285));
    InMux I__3120 (
            .O(N__34285),
            .I(N__34282));
    LocalMux I__3119 (
            .O(N__34282),
            .I(N__34279));
    Span4Mux_v I__3118 (
            .O(N__34279),
            .I(N__34276));
    Odrv4 I__3117 (
            .O(N__34276),
            .I(\pid_alt.error_i_regZ0Z_6 ));
    InMux I__3116 (
            .O(N__34273),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_5 ));
    CascadeMux I__3115 (
            .O(N__34270),
            .I(N__34267));
    InMux I__3114 (
            .O(N__34267),
            .I(N__34264));
    LocalMux I__3113 (
            .O(N__34264),
            .I(N__34261));
    Span4Mux_v I__3112 (
            .O(N__34261),
            .I(N__34258));
    Odrv4 I__3111 (
            .O(N__34258),
            .I(\pid_alt.error_i_regZ0Z_7 ));
    InMux I__3110 (
            .O(N__34255),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_6 ));
    CascadeMux I__3109 (
            .O(N__34252),
            .I(N__34249));
    InMux I__3108 (
            .O(N__34249),
            .I(N__34246));
    LocalMux I__3107 (
            .O(N__34246),
            .I(N__34243));
    Span4Mux_v I__3106 (
            .O(N__34243),
            .I(N__34240));
    Odrv4 I__3105 (
            .O(N__34240),
            .I(\pid_alt.error_i_regZ0Z_8 ));
    InMux I__3104 (
            .O(N__34237),
            .I(bfn_2_17_0_));
    CascadeMux I__3103 (
            .O(N__34234),
            .I(N__34231));
    InMux I__3102 (
            .O(N__34231),
            .I(N__34228));
    LocalMux I__3101 (
            .O(N__34228),
            .I(N__34225));
    Span4Mux_v I__3100 (
            .O(N__34225),
            .I(N__34222));
    Span4Mux_v I__3099 (
            .O(N__34222),
            .I(N__34219));
    Odrv4 I__3098 (
            .O(N__34219),
            .I(\pid_alt.error_i_regZ0Z_9 ));
    InMux I__3097 (
            .O(N__34216),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_8 ));
    CascadeMux I__3096 (
            .O(N__34213),
            .I(N__34210));
    InMux I__3095 (
            .O(N__34210),
            .I(N__34207));
    LocalMux I__3094 (
            .O(N__34207),
            .I(N__34204));
    Odrv12 I__3093 (
            .O(N__34204),
            .I(\pid_alt.error_i_regZ0Z_10 ));
    InMux I__3092 (
            .O(N__34201),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_9 ));
    CascadeMux I__3091 (
            .O(N__34198),
            .I(N__34195));
    InMux I__3090 (
            .O(N__34195),
            .I(N__34192));
    LocalMux I__3089 (
            .O(N__34192),
            .I(N__34189));
    Span4Mux_v I__3088 (
            .O(N__34189),
            .I(N__34186));
    Odrv4 I__3087 (
            .O(N__34186),
            .I(\pid_alt.error_i_regZ0Z_11 ));
    InMux I__3086 (
            .O(N__34183),
            .I(N__34180));
    LocalMux I__3085 (
            .O(N__34180),
            .I(N__34175));
    InMux I__3084 (
            .O(N__34179),
            .I(N__34170));
    InMux I__3083 (
            .O(N__34178),
            .I(N__34170));
    Odrv4 I__3082 (
            .O(N__34175),
            .I(\pid_alt.error_i_reg_esr_RNI4NMPZ0Z_11 ));
    LocalMux I__3081 (
            .O(N__34170),
            .I(\pid_alt.error_i_reg_esr_RNI4NMPZ0Z_11 ));
    InMux I__3080 (
            .O(N__34165),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_10 ));
    CascadeMux I__3079 (
            .O(N__34162),
            .I(N__34159));
    InMux I__3078 (
            .O(N__34159),
            .I(N__34156));
    LocalMux I__3077 (
            .O(N__34156),
            .I(\pid_alt.error_i_regZ0Z_1 ));
    InMux I__3076 (
            .O(N__34153),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_0 ));
    CascadeMux I__3075 (
            .O(N__34150),
            .I(N__34147));
    InMux I__3074 (
            .O(N__34147),
            .I(N__34144));
    LocalMux I__3073 (
            .O(N__34144),
            .I(N__34141));
    Span4Mux_v I__3072 (
            .O(N__34141),
            .I(N__34138));
    Odrv4 I__3071 (
            .O(N__34138),
            .I(\pid_alt.error_i_regZ0Z_2 ));
    InMux I__3070 (
            .O(N__34135),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_1 ));
    CascadeMux I__3069 (
            .O(N__34132),
            .I(N__34129));
    InMux I__3068 (
            .O(N__34129),
            .I(N__34126));
    LocalMux I__3067 (
            .O(N__34126),
            .I(N__34123));
    Span4Mux_v I__3066 (
            .O(N__34123),
            .I(N__34120));
    Odrv4 I__3065 (
            .O(N__34120),
            .I(\pid_alt.error_i_regZ0Z_3 ));
    InMux I__3064 (
            .O(N__34117),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_2 ));
    InMux I__3063 (
            .O(N__34114),
            .I(N__34105));
    InMux I__3062 (
            .O(N__34113),
            .I(N__34105));
    InMux I__3061 (
            .O(N__34112),
            .I(N__34105));
    LocalMux I__3060 (
            .O(N__34105),
            .I(\pid_alt.error_p_regZ0Z_1 ));
    CascadeMux I__3059 (
            .O(N__34102),
            .I(N__34098));
    InMux I__3058 (
            .O(N__34101),
            .I(N__34090));
    InMux I__3057 (
            .O(N__34098),
            .I(N__34090));
    InMux I__3056 (
            .O(N__34097),
            .I(N__34090));
    LocalMux I__3055 (
            .O(N__34090),
            .I(\pid_alt.error_d_reg_prevZ0Z_1 ));
    InMux I__3054 (
            .O(N__34087),
            .I(N__34081));
    InMux I__3053 (
            .O(N__34086),
            .I(N__34074));
    InMux I__3052 (
            .O(N__34085),
            .I(N__34074));
    InMux I__3051 (
            .O(N__34084),
            .I(N__34074));
    LocalMux I__3050 (
            .O(N__34081),
            .I(N__34069));
    LocalMux I__3049 (
            .O(N__34074),
            .I(N__34069));
    Sp12to4 I__3048 (
            .O(N__34069),
            .I(N__34066));
    Odrv12 I__3047 (
            .O(N__34066),
            .I(\pid_alt.error_d_regZ0Z_1 ));
    InMux I__3046 (
            .O(N__34063),
            .I(N__34060));
    LocalMux I__3045 (
            .O(N__34060),
            .I(\pid_alt.un1_pid_prereg_16_0 ));
    CascadeMux I__3044 (
            .O(N__34057),
            .I(\pid_alt.error_d_reg_prev_esr_RNITF511_0Z0Z_1_cascade_ ));
    InMux I__3043 (
            .O(N__34054),
            .I(N__34049));
    InMux I__3042 (
            .O(N__34053),
            .I(N__34044));
    InMux I__3041 (
            .O(N__34052),
            .I(N__34044));
    LocalMux I__3040 (
            .O(N__34049),
            .I(\pid_alt.error_d_regZ0Z_2 ));
    LocalMux I__3039 (
            .O(N__34044),
            .I(\pid_alt.error_d_regZ0Z_2 ));
    InMux I__3038 (
            .O(N__34039),
            .I(N__34035));
    InMux I__3037 (
            .O(N__34038),
            .I(N__34032));
    LocalMux I__3036 (
            .O(N__34035),
            .I(\pid_alt.error_d_reg_prevZ0Z_2 ));
    LocalMux I__3035 (
            .O(N__34032),
            .I(\pid_alt.error_d_reg_prevZ0Z_2 ));
    InMux I__3034 (
            .O(N__34027),
            .I(N__34024));
    LocalMux I__3033 (
            .O(N__34024),
            .I(\pid_alt.error_d_reg_prevZ0Z_0 ));
    InMux I__3032 (
            .O(N__34021),
            .I(N__34018));
    LocalMux I__3031 (
            .O(N__34018),
            .I(\pid_alt.error_d_reg_prev_esr_RNITF511Z0Z_1 ));
    InMux I__3030 (
            .O(N__34015),
            .I(N__34011));
    InMux I__3029 (
            .O(N__34014),
            .I(N__34008));
    LocalMux I__3028 (
            .O(N__34011),
            .I(\pid_alt.error_p_reg_esr_RNIOI4PZ0Z_0 ));
    LocalMux I__3027 (
            .O(N__34008),
            .I(\pid_alt.error_p_reg_esr_RNIOI4PZ0Z_0 ));
    CascadeMux I__3026 (
            .O(N__34003),
            .I(N__34000));
    InMux I__3025 (
            .O(N__34000),
            .I(N__33997));
    LocalMux I__3024 (
            .O(N__33997),
            .I(\pid_alt.error_d_reg_prev_esr_RNI0J511_0Z0Z_2 ));
    InMux I__3023 (
            .O(N__33994),
            .I(N__33990));
    InMux I__3022 (
            .O(N__33993),
            .I(N__33987));
    LocalMux I__3021 (
            .O(N__33990),
            .I(\pid_alt.error_d_reg_prev_esr_RNITF511_0Z0Z_1 ));
    LocalMux I__3020 (
            .O(N__33987),
            .I(\pid_alt.error_d_reg_prev_esr_RNITF511_0Z0Z_1 ));
    InMux I__3019 (
            .O(N__33982),
            .I(N__33979));
    LocalMux I__3018 (
            .O(N__33979),
            .I(N__33975));
    InMux I__3017 (
            .O(N__33978),
            .I(N__33971));
    Span4Mux_v I__3016 (
            .O(N__33975),
            .I(N__33968));
    InMux I__3015 (
            .O(N__33974),
            .I(N__33965));
    LocalMux I__3014 (
            .O(N__33971),
            .I(N__33962));
    Span4Mux_v I__3013 (
            .O(N__33968),
            .I(N__33959));
    LocalMux I__3012 (
            .O(N__33965),
            .I(N__33954));
    Span12Mux_v I__3011 (
            .O(N__33962),
            .I(N__33954));
    Odrv4 I__3010 (
            .O(N__33959),
            .I(\pid_alt.error_d_regZ0Z_17 ));
    Odrv12 I__3009 (
            .O(N__33954),
            .I(\pid_alt.error_d_regZ0Z_17 ));
    InMux I__3008 (
            .O(N__33949),
            .I(N__33945));
    CascadeMux I__3007 (
            .O(N__33948),
            .I(N__33942));
    LocalMux I__3006 (
            .O(N__33945),
            .I(N__33939));
    InMux I__3005 (
            .O(N__33942),
            .I(N__33936));
    Span4Mux_v I__3004 (
            .O(N__33939),
            .I(N__33931));
    LocalMux I__3003 (
            .O(N__33936),
            .I(N__33931));
    Span4Mux_v I__3002 (
            .O(N__33931),
            .I(N__33928));
    Odrv4 I__3001 (
            .O(N__33928),
            .I(\pid_alt.error_d_reg_prevZ0Z_17 ));
    InMux I__3000 (
            .O(N__33925),
            .I(N__33922));
    LocalMux I__2999 (
            .O(N__33922),
            .I(N__33919));
    Span4Mux_h I__2998 (
            .O(N__33919),
            .I(N__33916));
    Odrv4 I__2997 (
            .O(N__33916),
            .I(\pid_alt.O_4_12 ));
    InMux I__2996 (
            .O(N__33913),
            .I(N__33910));
    LocalMux I__2995 (
            .O(N__33910),
            .I(N__33907));
    Span4Mux_h I__2994 (
            .O(N__33907),
            .I(N__33904));
    Odrv4 I__2993 (
            .O(N__33904),
            .I(\pid_alt.O_4_14 ));
    InMux I__2992 (
            .O(N__33901),
            .I(N__33898));
    LocalMux I__2991 (
            .O(N__33898),
            .I(N__33895));
    Odrv4 I__2990 (
            .O(N__33895),
            .I(\pid_alt.O_4_4 ));
    InMux I__2989 (
            .O(N__33892),
            .I(N__33889));
    LocalMux I__2988 (
            .O(N__33889),
            .I(N__33886));
    Odrv12 I__2987 (
            .O(N__33886),
            .I(alt_ki_5));
    InMux I__2986 (
            .O(N__33883),
            .I(N__33880));
    LocalMux I__2985 (
            .O(N__33880),
            .I(N__33877));
    Span4Mux_s2_h I__2984 (
            .O(N__33877),
            .I(N__33874));
    Odrv4 I__2983 (
            .O(N__33874),
            .I(alt_ki_6));
    InMux I__2982 (
            .O(N__33871),
            .I(N__33867));
    InMux I__2981 (
            .O(N__33870),
            .I(N__33864));
    LocalMux I__2980 (
            .O(N__33867),
            .I(N__33859));
    LocalMux I__2979 (
            .O(N__33864),
            .I(N__33859));
    Odrv4 I__2978 (
            .O(N__33859),
            .I(\pid_alt.error_p_regZ0Z_2 ));
    CascadeMux I__2977 (
            .O(N__33856),
            .I(\pid_alt.error_d_reg_prev_esr_RNI0J511_0Z0Z_2_cascade_ ));
    InMux I__2976 (
            .O(N__33853),
            .I(N__33850));
    LocalMux I__2975 (
            .O(N__33850),
            .I(N__33847));
    Odrv4 I__2974 (
            .O(N__33847),
            .I(\pid_alt.O_5_20 ));
    InMux I__2973 (
            .O(N__33844),
            .I(N__33838));
    InMux I__2972 (
            .O(N__33843),
            .I(N__33838));
    LocalMux I__2971 (
            .O(N__33838),
            .I(N__33835));
    Odrv12 I__2970 (
            .O(N__33835),
            .I(\pid_alt.error_p_regZ0Z_16 ));
    InMux I__2969 (
            .O(N__33832),
            .I(N__33829));
    LocalMux I__2968 (
            .O(N__33829),
            .I(N__33826));
    Odrv4 I__2967 (
            .O(N__33826),
            .I(\pid_alt.O_3_5 ));
    InMux I__2966 (
            .O(N__33823),
            .I(N__33820));
    LocalMux I__2965 (
            .O(N__33820),
            .I(N__33817));
    Span4Mux_s2_h I__2964 (
            .O(N__33817),
            .I(N__33814));
    Odrv4 I__2963 (
            .O(N__33814),
            .I(alt_kd_0));
    InMux I__2962 (
            .O(N__33811),
            .I(N__33808));
    LocalMux I__2961 (
            .O(N__33808),
            .I(N__33805));
    Span4Mux_s2_h I__2960 (
            .O(N__33805),
            .I(N__33802));
    Odrv4 I__2959 (
            .O(N__33802),
            .I(alt_kd_1));
    InMux I__2958 (
            .O(N__33799),
            .I(N__33796));
    LocalMux I__2957 (
            .O(N__33796),
            .I(N__33793));
    Span4Mux_s2_h I__2956 (
            .O(N__33793),
            .I(N__33790));
    Odrv4 I__2955 (
            .O(N__33790),
            .I(alt_kd_2));
    InMux I__2954 (
            .O(N__33787),
            .I(N__33784));
    LocalMux I__2953 (
            .O(N__33784),
            .I(N__33781));
    Span4Mux_s2_h I__2952 (
            .O(N__33781),
            .I(N__33778));
    Odrv4 I__2951 (
            .O(N__33778),
            .I(alt_kd_3));
    InMux I__2950 (
            .O(N__33775),
            .I(N__33772));
    LocalMux I__2949 (
            .O(N__33772),
            .I(N__33769));
    Span4Mux_v I__2948 (
            .O(N__33769),
            .I(N__33766));
    Odrv4 I__2947 (
            .O(N__33766),
            .I(alt_kd_4));
    InMux I__2946 (
            .O(N__33763),
            .I(N__33760));
    LocalMux I__2945 (
            .O(N__33760),
            .I(N__33757));
    Span4Mux_v I__2944 (
            .O(N__33757),
            .I(N__33754));
    Odrv4 I__2943 (
            .O(N__33754),
            .I(alt_kd_5));
    InMux I__2942 (
            .O(N__33751),
            .I(N__33748));
    LocalMux I__2941 (
            .O(N__33748),
            .I(N__33745));
    Span4Mux_s3_h I__2940 (
            .O(N__33745),
            .I(N__33742));
    Odrv4 I__2939 (
            .O(N__33742),
            .I(alt_kd_6));
    InMux I__2938 (
            .O(N__33739),
            .I(N__33736));
    LocalMux I__2937 (
            .O(N__33736),
            .I(N__33733));
    Span4Mux_s3_h I__2936 (
            .O(N__33733),
            .I(N__33730));
    Odrv4 I__2935 (
            .O(N__33730),
            .I(alt_kd_7));
    InMux I__2934 (
            .O(N__33727),
            .I(N__33724));
    LocalMux I__2933 (
            .O(N__33724),
            .I(N__33721));
    Odrv4 I__2932 (
            .O(N__33721),
            .I(\pid_alt.O_5_11 ));
    InMux I__2931 (
            .O(N__33718),
            .I(N__33715));
    LocalMux I__2930 (
            .O(N__33715),
            .I(N__33712));
    Odrv4 I__2929 (
            .O(N__33712),
            .I(\pid_alt.O_5_12 ));
    InMux I__2928 (
            .O(N__33709),
            .I(N__33706));
    LocalMux I__2927 (
            .O(N__33706),
            .I(N__33703));
    Odrv4 I__2926 (
            .O(N__33703),
            .I(\pid_alt.O_5_13 ));
    InMux I__2925 (
            .O(N__33700),
            .I(N__33697));
    LocalMux I__2924 (
            .O(N__33697),
            .I(\pid_alt.O_5_7 ));
    InMux I__2923 (
            .O(N__33694),
            .I(N__33691));
    LocalMux I__2922 (
            .O(N__33691),
            .I(\pid_alt.O_5_15 ));
    InMux I__2921 (
            .O(N__33688),
            .I(N__33682));
    InMux I__2920 (
            .O(N__33687),
            .I(N__33682));
    LocalMux I__2919 (
            .O(N__33682),
            .I(N__33679));
    Odrv12 I__2918 (
            .O(N__33679),
            .I(\pid_alt.error_p_regZ0Z_11 ));
    InMux I__2917 (
            .O(N__33676),
            .I(N__33673));
    LocalMux I__2916 (
            .O(N__33673),
            .I(N__33670));
    Odrv4 I__2915 (
            .O(N__33670),
            .I(\pid_alt.O_5_16 ));
    InMux I__2914 (
            .O(N__33667),
            .I(N__33664));
    LocalMux I__2913 (
            .O(N__33664),
            .I(\pid_alt.O_5_14 ));
    InMux I__2912 (
            .O(N__33661),
            .I(N__33655));
    InMux I__2911 (
            .O(N__33660),
            .I(N__33655));
    LocalMux I__2910 (
            .O(N__33655),
            .I(N__33652));
    Span4Mux_v I__2909 (
            .O(N__33652),
            .I(N__33649));
    Odrv4 I__2908 (
            .O(N__33649),
            .I(\pid_alt.error_p_regZ0Z_10 ));
    InMux I__2907 (
            .O(N__33646),
            .I(N__33643));
    LocalMux I__2906 (
            .O(N__33643),
            .I(N__33640));
    Odrv4 I__2905 (
            .O(N__33640),
            .I(\pid_alt.O_5_18 ));
    InMux I__2904 (
            .O(N__33637),
            .I(N__33634));
    LocalMux I__2903 (
            .O(N__33634),
            .I(N__33631));
    Odrv4 I__2902 (
            .O(N__33631),
            .I(\pid_alt.O_5_19 ));
    InMux I__2901 (
            .O(N__33628),
            .I(N__33623));
    InMux I__2900 (
            .O(N__33627),
            .I(N__33618));
    InMux I__2899 (
            .O(N__33626),
            .I(N__33618));
    LocalMux I__2898 (
            .O(N__33623),
            .I(N__33613));
    LocalMux I__2897 (
            .O(N__33618),
            .I(N__33613));
    Span12Mux_v I__2896 (
            .O(N__33613),
            .I(N__33610));
    Odrv12 I__2895 (
            .O(N__33610),
            .I(\pid_alt.error_d_regZ0Z_16 ));
    InMux I__2894 (
            .O(N__33607),
            .I(N__33601));
    InMux I__2893 (
            .O(N__33606),
            .I(N__33601));
    LocalMux I__2892 (
            .O(N__33601),
            .I(\pid_alt.error_d_reg_prevZ0Z_16 ));
    InMux I__2891 (
            .O(N__33598),
            .I(N__33595));
    LocalMux I__2890 (
            .O(N__33595),
            .I(N__33592));
    Odrv4 I__2889 (
            .O(N__33592),
            .I(\pid_alt.O_5_4 ));
    CascadeMux I__2888 (
            .O(N__33589),
            .I(N__33586));
    InMux I__2887 (
            .O(N__33586),
            .I(N__33580));
    InMux I__2886 (
            .O(N__33585),
            .I(N__33580));
    LocalMux I__2885 (
            .O(N__33580),
            .I(N__33577));
    Odrv12 I__2884 (
            .O(N__33577),
            .I(\pid_alt.error_p_regZ0Z_0 ));
    InMux I__2883 (
            .O(N__33574),
            .I(N__33571));
    LocalMux I__2882 (
            .O(N__33571),
            .I(N__33568));
    Odrv4 I__2881 (
            .O(N__33568),
            .I(\pid_alt.O_5_10 ));
    InMux I__2880 (
            .O(N__33565),
            .I(N__33562));
    LocalMux I__2879 (
            .O(N__33562),
            .I(N__33559));
    Span4Mux_h I__2878 (
            .O(N__33559),
            .I(N__33556));
    Odrv4 I__2877 (
            .O(N__33556),
            .I(\pid_alt.O_5_22 ));
    InMux I__2876 (
            .O(N__33553),
            .I(N__33550));
    LocalMux I__2875 (
            .O(N__33550),
            .I(N__33547));
    Span4Mux_h I__2874 (
            .O(N__33547),
            .I(N__33544));
    Odrv4 I__2873 (
            .O(N__33544),
            .I(\pid_alt.O_5_23 ));
    InMux I__2872 (
            .O(N__33541),
            .I(N__33538));
    LocalMux I__2871 (
            .O(N__33538),
            .I(N__33535));
    Odrv4 I__2870 (
            .O(N__33535),
            .I(\pid_alt.O_5_17 ));
    InMux I__2869 (
            .O(N__33532),
            .I(N__33529));
    LocalMux I__2868 (
            .O(N__33529),
            .I(N__33526));
    Odrv4 I__2867 (
            .O(N__33526),
            .I(\pid_alt.O_5_9 ));
    InMux I__2866 (
            .O(N__33523),
            .I(N__33520));
    LocalMux I__2865 (
            .O(N__33520),
            .I(N__33517));
    Odrv4 I__2864 (
            .O(N__33517),
            .I(\pid_alt.O_5_21 ));
    InMux I__2863 (
            .O(N__33514),
            .I(N__33511));
    LocalMux I__2862 (
            .O(N__33511),
            .I(N__33508));
    Span4Mux_v I__2861 (
            .O(N__33508),
            .I(N__33504));
    InMux I__2860 (
            .O(N__33507),
            .I(N__33501));
    Span4Mux_v I__2859 (
            .O(N__33504),
            .I(N__33496));
    LocalMux I__2858 (
            .O(N__33501),
            .I(N__33496));
    Odrv4 I__2857 (
            .O(N__33496),
            .I(\pid_alt.error_p_regZ0Z_17 ));
    CascadeMux I__2856 (
            .O(N__33493),
            .I(\pid_alt.error_d_reg_prev_esr_RNIL8611Z0Z_9_cascade_ ));
    InMux I__2855 (
            .O(N__33490),
            .I(N__33487));
    LocalMux I__2854 (
            .O(N__33487),
            .I(\pid_alt.error_d_reg_prev_esr_RNIL8611Z0Z_9 ));
    InMux I__2853 (
            .O(N__33484),
            .I(N__33478));
    InMux I__2852 (
            .O(N__33483),
            .I(N__33478));
    LocalMux I__2851 (
            .O(N__33478),
            .I(\pid_alt.error_d_reg_prev_esr_RNIDAHM_0Z0Z_10 ));
    InMux I__2850 (
            .O(N__33475),
            .I(N__33472));
    LocalMux I__2849 (
            .O(N__33472),
            .I(\pid_alt.error_d_reg_prev_esr_RNI20IM_0Z0Z_17 ));
    CascadeMux I__2848 (
            .O(N__33469),
            .I(\pid_alt.error_d_reg_prev_esr_RNI20IM_0Z0Z_17_cascade_ ));
    InMux I__2847 (
            .O(N__33466),
            .I(N__33460));
    InMux I__2846 (
            .O(N__33465),
            .I(N__33460));
    LocalMux I__2845 (
            .O(N__33460),
            .I(\pid_alt.error_d_reg_prev_esr_RNIVSHMZ0Z_16 ));
    CascadeMux I__2844 (
            .O(N__33457),
            .I(\pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16_cascade_ ));
    CascadeMux I__2843 (
            .O(N__33454),
            .I(\pid_alt.error_d_reg_prev_esr_RNIGDHM_0Z0Z_11_cascade_ ));
    InMux I__2842 (
            .O(N__33451),
            .I(N__33448));
    LocalMux I__2841 (
            .O(N__33448),
            .I(\pid_alt.error_d_reg_prev_esr_RNIDAHMZ0Z_10 ));
    InMux I__2840 (
            .O(N__33445),
            .I(N__33442));
    LocalMux I__2839 (
            .O(N__33442),
            .I(\pid_alt.error_d_reg_prev_esr_RNIGDHM_0Z0Z_11 ));
    CascadeMux I__2838 (
            .O(N__33439),
            .I(\pid_alt.error_d_reg_prev_esr_RNIDAHMZ0Z_10_cascade_ ));
    InMux I__2837 (
            .O(N__33436),
            .I(N__33430));
    InMux I__2836 (
            .O(N__33435),
            .I(N__33430));
    LocalMux I__2835 (
            .O(N__33430),
            .I(N__33427));
    Span12Mux_v I__2834 (
            .O(N__33427),
            .I(N__33424));
    Odrv12 I__2833 (
            .O(N__33424),
            .I(\pid_alt.error_d_reg_prevZ0Z_10 ));
    InMux I__2832 (
            .O(N__33421),
            .I(N__33414));
    InMux I__2831 (
            .O(N__33420),
            .I(N__33414));
    InMux I__2830 (
            .O(N__33419),
            .I(N__33411));
    LocalMux I__2829 (
            .O(N__33414),
            .I(N__33408));
    LocalMux I__2828 (
            .O(N__33411),
            .I(N__33403));
    Span12Mux_v I__2827 (
            .O(N__33408),
            .I(N__33403));
    Odrv12 I__2826 (
            .O(N__33403),
            .I(\pid_alt.error_d_regZ0Z_10 ));
    InMux I__2825 (
            .O(N__33400),
            .I(N__33394));
    InMux I__2824 (
            .O(N__33399),
            .I(N__33394));
    LocalMux I__2823 (
            .O(N__33394),
            .I(\pid_alt.error_d_reg_prevZ0Z_11 ));
    InMux I__2822 (
            .O(N__33391),
            .I(N__33382));
    InMux I__2821 (
            .O(N__33390),
            .I(N__33382));
    InMux I__2820 (
            .O(N__33389),
            .I(N__33382));
    LocalMux I__2819 (
            .O(N__33382),
            .I(N__33379));
    Span12Mux_v I__2818 (
            .O(N__33379),
            .I(N__33376));
    Odrv12 I__2817 (
            .O(N__33376),
            .I(\pid_alt.error_d_regZ0Z_11 ));
    InMux I__2816 (
            .O(N__33373),
            .I(N__33370));
    LocalMux I__2815 (
            .O(N__33370),
            .I(N__33367));
    Span4Mux_h I__2814 (
            .O(N__33367),
            .I(N__33364));
    Span4Mux_v I__2813 (
            .O(N__33364),
            .I(N__33361));
    Odrv4 I__2812 (
            .O(N__33361),
            .I(\pid_alt.O_5_24 ));
    CascadeMux I__2811 (
            .O(N__33358),
            .I(\pid_alt.error_p_reg_esr_RNIOI4PZ0Z_0_cascade_ ));
    InMux I__2810 (
            .O(N__33355),
            .I(N__33346));
    InMux I__2809 (
            .O(N__33354),
            .I(N__33346));
    InMux I__2808 (
            .O(N__33353),
            .I(N__33346));
    LocalMux I__2807 (
            .O(N__33346),
            .I(N__33343));
    Odrv4 I__2806 (
            .O(N__33343),
            .I(\pid_alt.error_d_regZ0Z_0 ));
    InMux I__2805 (
            .O(N__33340),
            .I(N__33337));
    LocalMux I__2804 (
            .O(N__33337),
            .I(N__33334));
    Odrv4 I__2803 (
            .O(N__33334),
            .I(\pid_front.O_0_23 ));
    InMux I__2802 (
            .O(N__33331),
            .I(N__33328));
    LocalMux I__2801 (
            .O(N__33328),
            .I(N__33325));
    Span4Mux_v I__2800 (
            .O(N__33325),
            .I(N__33322));
    Odrv4 I__2799 (
            .O(N__33322),
            .I(\pid_alt.O_4_5 ));
    InMux I__2798 (
            .O(N__33319),
            .I(N__33316));
    LocalMux I__2797 (
            .O(N__33316),
            .I(N__33313));
    Span4Mux_v I__2796 (
            .O(N__33313),
            .I(N__33310));
    Odrv4 I__2795 (
            .O(N__33310),
            .I(\pid_alt.O_4_8 ));
    InMux I__2794 (
            .O(N__33307),
            .I(N__33304));
    LocalMux I__2793 (
            .O(N__33304),
            .I(N__33301));
    Span4Mux_v I__2792 (
            .O(N__33301),
            .I(N__33298));
    Odrv4 I__2791 (
            .O(N__33298),
            .I(\pid_alt.O_4_9 ));
    InMux I__2790 (
            .O(N__33295),
            .I(N__33292));
    LocalMux I__2789 (
            .O(N__33292),
            .I(N__33289));
    Odrv4 I__2788 (
            .O(N__33289),
            .I(\pid_alt.O_4_6 ));
    InMux I__2787 (
            .O(N__33286),
            .I(N__33283));
    LocalMux I__2786 (
            .O(N__33283),
            .I(N__33280));
    Span4Mux_v I__2785 (
            .O(N__33280),
            .I(N__33277));
    Span4Mux_v I__2784 (
            .O(N__33277),
            .I(N__33274));
    Odrv4 I__2783 (
            .O(N__33274),
            .I(\pid_alt.O_5_6 ));
    InMux I__2782 (
            .O(N__33271),
            .I(N__33268));
    LocalMux I__2781 (
            .O(N__33268),
            .I(N__33265));
    Span4Mux_v I__2780 (
            .O(N__33265),
            .I(N__33262));
    Span4Mux_v I__2779 (
            .O(N__33262),
            .I(N__33259));
    Odrv4 I__2778 (
            .O(N__33259),
            .I(\pid_alt.O_3_6 ));
    InMux I__2777 (
            .O(N__33256),
            .I(N__33253));
    LocalMux I__2776 (
            .O(N__33253),
            .I(N__33250));
    Span4Mux_v I__2775 (
            .O(N__33250),
            .I(N__33247));
    Span4Mux_v I__2774 (
            .O(N__33247),
            .I(N__33244));
    Odrv4 I__2773 (
            .O(N__33244),
            .I(\pid_alt.O_5_8 ));
    InMux I__2772 (
            .O(N__33241),
            .I(N__33238));
    LocalMux I__2771 (
            .O(N__33238),
            .I(N__33235));
    Odrv4 I__2770 (
            .O(N__33235),
            .I(\pid_alt.O_4_22 ));
    InMux I__2769 (
            .O(N__33232),
            .I(N__33229));
    LocalMux I__2768 (
            .O(N__33229),
            .I(N__33226));
    Odrv4 I__2767 (
            .O(N__33226),
            .I(\pid_alt.O_4_24 ));
    InMux I__2766 (
            .O(N__33223),
            .I(N__33220));
    LocalMux I__2765 (
            .O(N__33220),
            .I(\pid_alt.O_4_7 ));
    InMux I__2764 (
            .O(N__33217),
            .I(N__33214));
    LocalMux I__2763 (
            .O(N__33214),
            .I(\pid_alt.O_4_15 ));
    InMux I__2762 (
            .O(N__33211),
            .I(N__33208));
    LocalMux I__2761 (
            .O(N__33208),
            .I(\pid_alt.O_4_10 ));
    InMux I__2760 (
            .O(N__33205),
            .I(N__33202));
    LocalMux I__2759 (
            .O(N__33202),
            .I(\pid_alt.O_4_11 ));
    InMux I__2758 (
            .O(N__33199),
            .I(N__33196));
    LocalMux I__2757 (
            .O(N__33196),
            .I(\pid_alt.O_4_21 ));
    InMux I__2756 (
            .O(N__33193),
            .I(N__33190));
    LocalMux I__2755 (
            .O(N__33190),
            .I(N__33187));
    Span4Mux_v I__2754 (
            .O(N__33187),
            .I(N__33184));
    Odrv4 I__2753 (
            .O(N__33184),
            .I(\pid_alt.O_3_4 ));
    InMux I__2752 (
            .O(N__33181),
            .I(N__33178));
    LocalMux I__2751 (
            .O(N__33178),
            .I(N__33175));
    Span4Mux_v I__2750 (
            .O(N__33175),
            .I(N__33172));
    Span4Mux_v I__2749 (
            .O(N__33172),
            .I(N__33169));
    Odrv4 I__2748 (
            .O(N__33169),
            .I(\pid_alt.O_5_5 ));
    InMux I__2747 (
            .O(N__33166),
            .I(N__33163));
    LocalMux I__2746 (
            .O(N__33163),
            .I(\pid_alt.O_3_13 ));
    InMux I__2745 (
            .O(N__33160),
            .I(N__33157));
    LocalMux I__2744 (
            .O(N__33157),
            .I(\pid_alt.O_3_16 ));
    InMux I__2743 (
            .O(N__33154),
            .I(N__33151));
    LocalMux I__2742 (
            .O(N__33151),
            .I(N__33148));
    Span4Mux_h I__2741 (
            .O(N__33148),
            .I(N__33145));
    Odrv4 I__2740 (
            .O(N__33145),
            .I(\pid_alt.O_4_13 ));
    InMux I__2739 (
            .O(N__33142),
            .I(N__33139));
    LocalMux I__2738 (
            .O(N__33139),
            .I(N__33136));
    Odrv4 I__2737 (
            .O(N__33136),
            .I(\pid_alt.O_4_18 ));
    InMux I__2736 (
            .O(N__33133),
            .I(N__33130));
    LocalMux I__2735 (
            .O(N__33130),
            .I(N__33127));
    Odrv4 I__2734 (
            .O(N__33127),
            .I(\pid_alt.O_4_19 ));
    InMux I__2733 (
            .O(N__33124),
            .I(N__33121));
    LocalMux I__2732 (
            .O(N__33121),
            .I(N__33118));
    Odrv4 I__2731 (
            .O(N__33118),
            .I(\pid_alt.O_4_20 ));
    InMux I__2730 (
            .O(N__33115),
            .I(N__33112));
    LocalMux I__2729 (
            .O(N__33112),
            .I(N__33109));
    Odrv4 I__2728 (
            .O(N__33109),
            .I(\pid_alt.O_4_16 ));
    InMux I__2727 (
            .O(N__33106),
            .I(N__33103));
    LocalMux I__2726 (
            .O(N__33103),
            .I(N__33100));
    Odrv4 I__2725 (
            .O(N__33100),
            .I(\pid_alt.O_4_17 ));
    InMux I__2724 (
            .O(N__33097),
            .I(N__33094));
    LocalMux I__2723 (
            .O(N__33094),
            .I(N__33091));
    Odrv4 I__2722 (
            .O(N__33091),
            .I(\pid_alt.O_4_23 ));
    InMux I__2721 (
            .O(N__33088),
            .I(N__33085));
    LocalMux I__2720 (
            .O(N__33085),
            .I(N__33082));
    Odrv4 I__2719 (
            .O(N__33082),
            .I(\pid_alt.O_3_19 ));
    InMux I__2718 (
            .O(N__33079),
            .I(N__33076));
    LocalMux I__2717 (
            .O(N__33076),
            .I(\pid_alt.O_3_21 ));
    InMux I__2716 (
            .O(N__33073),
            .I(N__33070));
    LocalMux I__2715 (
            .O(N__33070),
            .I(\pid_alt.O_3_17 ));
    InMux I__2714 (
            .O(N__33067),
            .I(N__33064));
    LocalMux I__2713 (
            .O(N__33064),
            .I(N__33061));
    Odrv4 I__2712 (
            .O(N__33061),
            .I(\pid_alt.O_3_24 ));
    InMux I__2711 (
            .O(N__33058),
            .I(N__33055));
    LocalMux I__2710 (
            .O(N__33055),
            .I(\pid_alt.O_3_7 ));
    InMux I__2709 (
            .O(N__33052),
            .I(N__33049));
    LocalMux I__2708 (
            .O(N__33049),
            .I(\pid_alt.O_3_15 ));
    InMux I__2707 (
            .O(N__33046),
            .I(N__33043));
    LocalMux I__2706 (
            .O(N__33043),
            .I(\pid_alt.O_3_9 ));
    InMux I__2705 (
            .O(N__33040),
            .I(N__33037));
    LocalMux I__2704 (
            .O(N__33037),
            .I(\pid_alt.O_3_10 ));
    InMux I__2703 (
            .O(N__33034),
            .I(N__33031));
    LocalMux I__2702 (
            .O(N__33031),
            .I(\pid_alt.O_3_11 ));
    InMux I__2701 (
            .O(N__33028),
            .I(N__33025));
    LocalMux I__2700 (
            .O(N__33025),
            .I(\pid_alt.O_3_12 ));
    InMux I__2699 (
            .O(N__33022),
            .I(N__33019));
    LocalMux I__2698 (
            .O(N__33019),
            .I(\pid_alt.O_3_14 ));
    InMux I__2697 (
            .O(N__33016),
            .I(N__33013));
    LocalMux I__2696 (
            .O(N__33013),
            .I(\pid_alt.O_3_8 ));
    InMux I__2695 (
            .O(N__33010),
            .I(N__33007));
    LocalMux I__2694 (
            .O(N__33007),
            .I(N__33004));
    Odrv4 I__2693 (
            .O(N__33004),
            .I(\pid_alt.O_3_18 ));
    InMux I__2692 (
            .O(N__33001),
            .I(N__32998));
    LocalMux I__2691 (
            .O(N__32998),
            .I(N__32995));
    Odrv4 I__2690 (
            .O(N__32995),
            .I(\pid_alt.O_3_22 ));
    InMux I__2689 (
            .O(N__32992),
            .I(N__32989));
    LocalMux I__2688 (
            .O(N__32989),
            .I(N__32986));
    Odrv4 I__2687 (
            .O(N__32986),
            .I(\pid_alt.O_3_20 ));
    IoInMux I__2686 (
            .O(N__32983),
            .I(N__32980));
    LocalMux I__2685 (
            .O(N__32980),
            .I(N__32977));
    IoSpan4Mux I__2684 (
            .O(N__32977),
            .I(N__32974));
    Span4Mux_s2_v I__2683 (
            .O(N__32974),
            .I(N__32971));
    Span4Mux_h I__2682 (
            .O(N__32971),
            .I(N__32968));
    Sp12to4 I__2681 (
            .O(N__32968),
            .I(N__32965));
    Span12Mux_s8_v I__2680 (
            .O(N__32965),
            .I(N__32962));
    Span12Mux_v I__2679 (
            .O(N__32962),
            .I(N__32959));
    Odrv12 I__2678 (
            .O(N__32959),
            .I(\Pc2drone_pll_inst.clk_system_pll ));
    defparam IN_MUX_bfv_16_4_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_4_0_));
    defparam IN_MUX_bfv_16_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_5_0_ (
            .carryinitin(\pid_side.un1_pid_prereg_0_cry_6 ),
            .carryinitout(bfn_16_5_0_));
    defparam IN_MUX_bfv_16_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_6_0_ (
            .carryinitin(\pid_side.un1_pid_prereg_0_cry_14 ),
            .carryinitout(bfn_16_6_0_));
    defparam IN_MUX_bfv_16_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_7_0_ (
            .carryinitin(\pid_side.un1_pid_prereg_0_cry_22 ),
            .carryinitout(bfn_16_7_0_));
    defparam IN_MUX_bfv_13_23_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_23_0_));
    defparam IN_MUX_bfv_13_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_24_0_ (
            .carryinitin(\pid_front.un1_pid_prereg_0_cry_6 ),
            .carryinitout(bfn_13_24_0_));
    defparam IN_MUX_bfv_13_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_25_0_ (
            .carryinitin(\pid_front.un1_pid_prereg_0_cry_14 ),
            .carryinitout(bfn_13_25_0_));
    defparam IN_MUX_bfv_13_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_26_0_ (
            .carryinitin(\pid_front.un1_pid_prereg_0_cry_22 ),
            .carryinitout(bfn_13_26_0_));
    defparam IN_MUX_bfv_4_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_13_0_));
    defparam IN_MUX_bfv_4_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_14_0_ (
            .carryinitin(\pid_alt.un1_pid_prereg_0_cry_6 ),
            .carryinitout(bfn_4_14_0_));
    defparam IN_MUX_bfv_4_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_15_0_ (
            .carryinitin(\pid_alt.un1_pid_prereg_0_cry_14 ),
            .carryinitout(bfn_4_15_0_));
    defparam IN_MUX_bfv_4_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_16_0_ (
            .carryinitin(\pid_alt.un1_pid_prereg_0_cry_22 ),
            .carryinitout(bfn_4_16_0_));
    defparam IN_MUX_bfv_8_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_11_0_));
    defparam IN_MUX_bfv_8_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_12_0_ (
            .carryinitin(\scaler_4.un3_source_data_0_cry_7 ),
            .carryinitout(bfn_8_12_0_));
    defparam IN_MUX_bfv_7_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_11_0_));
    defparam IN_MUX_bfv_7_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_12_0_ (
            .carryinitin(\scaler_4.un2_source_data_0_cry_8 ),
            .carryinitout(bfn_7_12_0_));
    defparam IN_MUX_bfv_11_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_13_0_));
    defparam IN_MUX_bfv_11_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_14_0_ (
            .carryinitin(\reset_module_System.count_1_cry_8 ),
            .carryinitout(bfn_11_14_0_));
    defparam IN_MUX_bfv_11_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_15_0_ (
            .carryinitin(\reset_module_System.count_1_cry_16 ),
            .carryinitout(bfn_11_15_0_));
    defparam IN_MUX_bfv_4_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_9_0_));
    defparam IN_MUX_bfv_4_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_10_0_ (
            .carryinitin(\ppm_encoder_1.un1_throttle_cry_7 ),
            .carryinitout(bfn_4_10_0_));
    defparam IN_MUX_bfv_7_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_9_0_));
    defparam IN_MUX_bfv_7_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_10_0_ (
            .carryinitin(\ppm_encoder_1.un1_rudder_cry_13 ),
            .carryinitout(bfn_7_10_0_));
    defparam IN_MUX_bfv_10_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_7_0_));
    defparam IN_MUX_bfv_10_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_8_0_ (
            .carryinitin(\ppm_encoder_1.un1_elevator_cry_7 ),
            .carryinitout(bfn_10_8_0_));
    defparam IN_MUX_bfv_10_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_10_0_));
    defparam IN_MUX_bfv_10_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_11_0_ (
            .carryinitin(\ppm_encoder_1.un1_aileron_cry_7 ),
            .carryinitout(bfn_10_11_0_));
    defparam IN_MUX_bfv_8_1_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_1_0_));
    defparam IN_MUX_bfv_8_2_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_2_0_ (
            .carryinitin(\ppm_encoder_1.un1_init_pulses_3_cry_7 ),
            .carryinitout(bfn_8_2_0_));
    defparam IN_MUX_bfv_8_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_3_0_ (
            .carryinitin(\ppm_encoder_1.un1_init_pulses_3_cry_15 ),
            .carryinitout(bfn_8_3_0_));
    defparam IN_MUX_bfv_9_2_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_2_0_));
    defparam IN_MUX_bfv_9_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_3_0_ (
            .carryinitin(\ppm_encoder_1.un1_init_pulses_0_cry_7 ),
            .carryinitout(bfn_9_3_0_));
    defparam IN_MUX_bfv_9_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_4_0_ (
            .carryinitin(\ppm_encoder_1.un1_init_pulses_0_cry_15 ),
            .carryinitout(bfn_9_4_0_));
    defparam IN_MUX_bfv_10_1_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_1_0_));
    defparam IN_MUX_bfv_10_2_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_2_0_ (
            .carryinitin(\ppm_encoder_1.counter24_0_data_tmp_7 ),
            .carryinitout(bfn_10_2_0_));
    defparam IN_MUX_bfv_14_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_3_0_));
    defparam IN_MUX_bfv_14_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_4_0_ (
            .carryinitin(\pid_side.un11lto30_i_a2_6 ),
            .carryinitout(bfn_14_4_0_));
    defparam IN_MUX_bfv_11_22_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_22_0_));
    defparam IN_MUX_bfv_11_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_23_0_ (
            .carryinitin(\pid_front.un11lto30_i_a2_6 ),
            .carryinitout(bfn_11_23_0_));
    defparam IN_MUX_bfv_4_18_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_18_0_));
    defparam IN_MUX_bfv_4_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_19_0_ (
            .carryinitin(\pid_alt.error_cry_7 ),
            .carryinitout(bfn_4_19_0_));
    defparam IN_MUX_bfv_7_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_19_0_));
    defparam IN_MUX_bfv_10_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_12_0_));
    defparam IN_MUX_bfv_12_2_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_2_0_));
    defparam IN_MUX_bfv_12_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_3_0_ (
            .carryinitin(\ppm_encoder_1.un1_counter_13_cry_7 ),
            .carryinitout(bfn_12_3_0_));
    defparam IN_MUX_bfv_12_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_4_0_ (
            .carryinitin(\ppm_encoder_1.un1_counter_13_cry_15 ),
            .carryinitout(bfn_12_4_0_));
    defparam IN_MUX_bfv_15_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_8_0_));
    defparam IN_MUX_bfv_15_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_9_0_ (
            .carryinitin(\pid_side.un1_error_i_acumm_prereg_cry_7 ),
            .carryinitout(bfn_15_9_0_));
    defparam IN_MUX_bfv_15_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_10_0_ (
            .carryinitin(\pid_side.un1_error_i_acumm_prereg_cry_15 ),
            .carryinitout(bfn_15_10_0_));
    defparam IN_MUX_bfv_15_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_11_0_ (
            .carryinitin(\pid_side.un1_error_i_acumm_prereg_cry_23 ),
            .carryinitout(bfn_15_11_0_));
    defparam IN_MUX_bfv_20_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_20_15_0_));
    defparam IN_MUX_bfv_20_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_16_0_ (
            .carryinitin(\pid_side.error_cry_3_0 ),
            .carryinitout(bfn_20_16_0_));
    defparam IN_MUX_bfv_15_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_19_0_));
    defparam IN_MUX_bfv_15_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_20_0_ (
            .carryinitin(\pid_front.un1_error_i_acumm_prereg_cry_7 ),
            .carryinitout(bfn_15_20_0_));
    defparam IN_MUX_bfv_15_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_21_0_ (
            .carryinitin(\pid_front.un1_error_i_acumm_prereg_cry_15 ),
            .carryinitout(bfn_15_21_0_));
    defparam IN_MUX_bfv_15_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_22_0_ (
            .carryinitin(\pid_front.un1_error_i_acumm_prereg_cry_23 ),
            .carryinitout(bfn_15_22_0_));
    defparam IN_MUX_bfv_12_18_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_18_0_));
    defparam IN_MUX_bfv_12_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_19_0_ (
            .carryinitin(\pid_front.error_cry_3_0 ),
            .carryinitout(bfn_12_19_0_));
    defparam IN_MUX_bfv_2_16_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_16_0_));
    defparam IN_MUX_bfv_2_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_17_0_ (
            .carryinitin(\pid_alt.un1_error_i_acumm_prereg_cry_7 ),
            .carryinitout(bfn_2_17_0_));
    defparam IN_MUX_bfv_2_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_18_0_ (
            .carryinitin(\pid_alt.un1_error_i_acumm_prereg_cry_15 ),
            .carryinitout(bfn_2_18_0_));
    defparam IN_MUX_bfv_8_18_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_18_0_));
    defparam IN_MUX_bfv_8_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_19_0_ (
            .carryinitin(\dron_frame_decoder_1.un1_WDT_cry_7 ),
            .carryinitout(bfn_8_19_0_));
    defparam IN_MUX_bfv_8_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_13_0_));
    defparam IN_MUX_bfv_8_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_14_0_ (
            .carryinitin(\Commands_frame_decoder.un1_WDT_cry_7 ),
            .carryinitout(bfn_8_14_0_));
    ICE_GB \reset_module_System.reset_RNITC69  (
            .USERSIGNALTOGLOBALBUFFER(N__71045),
            .GLOBALBUFFEROUTPUT(N_934_g));
    ICE_GB \reset_module_System.reset_iso_RNI7G1  (
            .USERSIGNALTOGLOBALBUFFER(N__51655),
            .GLOBALBUFFEROUTPUT(reset_module_System_reset_iso_g));
    ICE_GB \pid_alt.state_RNICP2N1_0_0  (
            .USERSIGNALTOGLOBALBUFFER(N__45202),
            .GLOBALBUFFEROUTPUT(\pid_alt.N_933_0_g ));
    ICE_GB \pid_side.state_RNIV8D6_0_0  (
            .USERSIGNALTOGLOBALBUFFER(N__56344),
            .GLOBALBUFFEROUTPUT(\pid_side.state_0_g_0 ));
    ICE_GB \pid_alt.state_RNIR49E_0_0  (
            .USERSIGNALTOGLOBALBUFFER(N__61279),
            .GLOBALBUFFEROUTPUT(\pid_alt.state_0_g_0 ));
    ICE_GB \Pc2drone_pll_inst.PLLOUTCORE_derived_clock_RNI5FOA  (
            .USERSIGNALTOGLOBALBUFFER(N__32983),
            .GLOBALBUFFEROUTPUT(clk_system_pll_g));
    ICE_GB \pid_front.state_RNI3OO4_0_0  (
            .USERSIGNALTOGLOBALBUFFER(N__41518),
            .GLOBALBUFFEROUTPUT(\pid_front.state_0_g_0 ));
    ICE_GB \pid_side.state_RNIIIOO_0_0  (
            .USERSIGNALTOGLOBALBUFFER(N__60832),
            .GLOBALBUFFEROUTPUT(\pid_side.N_2054_g ));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \pid_alt.error_d_reg_esr_8_LC_1_5_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_8_LC_1_5_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_8_LC_1_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_8_LC_1_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33028),
            .lcout(\pid_alt.error_d_regZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94198),
            .ce(N__34725),
            .sr(N__92967));
    defparam \pid_alt.error_d_reg_esr_10_LC_1_5_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_10_LC_1_5_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_10_LC_1_5_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_10_LC_1_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33022),
            .lcout(\pid_alt.error_d_regZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94198),
            .ce(N__34725),
            .sr(N__92967));
    defparam \pid_alt.error_d_reg_esr_4_LC_1_5_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_4_LC_1_5_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_4_LC_1_5_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_4_LC_1_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33016),
            .lcout(\pid_alt.error_d_regZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94198),
            .ce(N__34725),
            .sr(N__92967));
    defparam \pid_alt.error_d_reg_esr_14_LC_1_5_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_14_LC_1_5_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_14_LC_1_5_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_14_LC_1_5_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33010),
            .lcout(\pid_alt.error_d_regZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94198),
            .ce(N__34725),
            .sr(N__92967));
    defparam \pid_alt.error_d_reg_esr_18_LC_1_5_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_18_LC_1_5_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_18_LC_1_5_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_18_LC_1_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33001),
            .lcout(\pid_alt.error_d_regZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94198),
            .ce(N__34725),
            .sr(N__92967));
    defparam \pid_alt.error_d_reg_esr_16_LC_1_5_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_16_LC_1_5_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_16_LC_1_5_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_16_LC_1_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32992),
            .lcout(\pid_alt.error_d_regZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94198),
            .ce(N__34725),
            .sr(N__92967));
    defparam \pid_alt.error_d_reg_esr_15_LC_1_5_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_15_LC_1_5_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_15_LC_1_5_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_15_LC_1_5_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33088),
            .lcout(\pid_alt.error_d_regZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94198),
            .ce(N__34725),
            .sr(N__92967));
    defparam \pid_alt.error_d_reg_esr_17_LC_1_6_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_17_LC_1_6_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_17_LC_1_6_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_17_LC_1_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33079),
            .lcout(\pid_alt.error_d_regZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94216),
            .ce(N__34726),
            .sr(N__92968));
    defparam \pid_alt.error_d_reg_esr_13_LC_1_6_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_13_LC_1_6_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_13_LC_1_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_13_LC_1_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33073),
            .lcout(\pid_alt.error_d_regZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94216),
            .ce(N__34726),
            .sr(N__92968));
    defparam \pid_alt.error_d_reg_esr_20_LC_1_6_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_20_LC_1_6_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_20_LC_1_6_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_20_LC_1_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33067),
            .lcout(\pid_alt.error_d_regZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94216),
            .ce(N__34726),
            .sr(N__92968));
    defparam \pid_alt.error_d_reg_esr_3_LC_1_6_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_3_LC_1_6_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_3_LC_1_6_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_3_LC_1_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33058),
            .lcout(\pid_alt.error_d_regZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94216),
            .ce(N__34726),
            .sr(N__92968));
    defparam \pid_alt.error_d_reg_esr_11_LC_1_6_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_11_LC_1_6_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_11_LC_1_6_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_11_LC_1_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33052),
            .lcout(\pid_alt.error_d_regZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94216),
            .ce(N__34726),
            .sr(N__92968));
    defparam \pid_alt.error_d_reg_esr_5_LC_1_6_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_5_LC_1_6_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_5_LC_1_6_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_5_LC_1_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33046),
            .lcout(\pid_alt.error_d_regZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94216),
            .ce(N__34726),
            .sr(N__92968));
    defparam \pid_alt.error_d_reg_esr_6_LC_1_6_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_6_LC_1_6_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_6_LC_1_6_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_6_LC_1_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33040),
            .lcout(\pid_alt.error_d_regZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94216),
            .ce(N__34726),
            .sr(N__92968));
    defparam \pid_alt.error_d_reg_esr_7_LC_1_6_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_7_LC_1_6_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_7_LC_1_6_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_7_LC_1_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33034),
            .lcout(\pid_alt.error_d_regZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94216),
            .ce(N__34726),
            .sr(N__92968));
    defparam \pid_alt.error_d_reg_esr_9_LC_1_7_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_9_LC_1_7_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_9_LC_1_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_9_LC_1_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33166),
            .lcout(\pid_alt.error_d_regZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94232),
            .ce(N__34727),
            .sr(N__92969));
    defparam \pid_alt.error_d_reg_esr_12_LC_1_7_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_12_LC_1_7_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_12_LC_1_7_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_12_LC_1_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33160),
            .lcout(\pid_alt.error_d_regZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94232),
            .ce(N__34727),
            .sr(N__92969));
    defparam \pid_alt.error_d_reg_prev_esr_10_LC_1_8_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_10_LC_1_8_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_10_LC_1_8_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_10_LC_1_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33419),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94248),
            .ce(N__40516),
            .sr(N__86514));
    defparam \pid_alt.error_i_reg_esr_9_LC_1_9_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_9_LC_1_9_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_9_LC_1_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_9_LC_1_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33154),
            .lcout(\pid_alt.error_i_regZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94265),
            .ce(N__34728),
            .sr(N__92970));
    defparam \pid_alt.error_i_reg_esr_14_LC_1_10_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_14_LC_1_10_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_14_LC_1_10_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_i_reg_esr_14_LC_1_10_0  (
            .in0(N__33142),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_i_regZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94284),
            .ce(N__34730),
            .sr(N__92972));
    defparam \pid_alt.error_i_reg_esr_15_LC_1_10_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_15_LC_1_10_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_15_LC_1_10_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_i_reg_esr_15_LC_1_10_1  (
            .in0(N__33133),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_i_regZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94284),
            .ce(N__34730),
            .sr(N__92972));
    defparam \pid_alt.error_i_reg_esr_16_LC_1_10_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_16_LC_1_10_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_16_LC_1_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_16_LC_1_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33124),
            .lcout(\pid_alt.error_i_regZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94284),
            .ce(N__34730),
            .sr(N__92972));
    defparam \pid_alt.error_i_reg_esr_12_LC_1_10_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_12_LC_1_10_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_12_LC_1_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_12_LC_1_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33115),
            .lcout(\pid_alt.error_i_regZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94284),
            .ce(N__34730),
            .sr(N__92972));
    defparam \pid_alt.error_i_reg_esr_13_LC_1_10_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_13_LC_1_10_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_13_LC_1_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_13_LC_1_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33106),
            .lcout(\pid_alt.error_i_regZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94284),
            .ce(N__34730),
            .sr(N__92972));
    defparam \pid_alt.error_i_reg_esr_19_LC_1_10_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_19_LC_1_10_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_19_LC_1_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_19_LC_1_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33097),
            .lcout(\pid_alt.error_i_regZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94284),
            .ce(N__34730),
            .sr(N__92972));
    defparam \pid_alt.error_i_reg_esr_18_LC_1_10_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_18_LC_1_10_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_18_LC_1_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_18_LC_1_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33241),
            .lcout(\pid_alt.error_i_regZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94284),
            .ce(N__34730),
            .sr(N__92972));
    defparam \pid_alt.error_i_reg_esr_20_LC_1_10_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_20_LC_1_10_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_20_LC_1_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_20_LC_1_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33232),
            .lcout(\pid_alt.error_i_regZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94284),
            .ce(N__34730),
            .sr(N__92972));
    defparam \pid_alt.error_i_reg_esr_3_LC_1_11_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_3_LC_1_11_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_3_LC_1_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_3_LC_1_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33223),
            .lcout(\pid_alt.error_i_regZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94299),
            .ce(N__34731),
            .sr(N__92973));
    defparam \pid_alt.error_i_reg_esr_11_LC_1_11_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_11_LC_1_11_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_11_LC_1_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_11_LC_1_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33217),
            .lcout(\pid_alt.error_i_regZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94299),
            .ce(N__34731),
            .sr(N__92973));
    defparam \pid_alt.error_i_reg_esr_6_LC_1_11_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_6_LC_1_11_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_6_LC_1_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_6_LC_1_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33211),
            .lcout(\pid_alt.error_i_regZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94299),
            .ce(N__34731),
            .sr(N__92973));
    defparam \pid_alt.error_i_reg_esr_7_LC_1_11_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_7_LC_1_11_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_7_LC_1_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_7_LC_1_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33205),
            .lcout(\pid_alt.error_i_regZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94299),
            .ce(N__34731),
            .sr(N__92973));
    defparam \pid_alt.error_i_reg_esr_17_LC_1_11_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_17_LC_1_11_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_17_LC_1_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_17_LC_1_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33199),
            .lcout(\pid_alt.error_i_regZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94299),
            .ce(N__34731),
            .sr(N__92973));
    defparam \pid_alt.error_d_reg_esr_0_LC_1_11_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_0_LC_1_11_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_0_LC_1_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_0_LC_1_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33193),
            .lcout(\pid_alt.error_d_regZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94299),
            .ce(N__34731),
            .sr(N__92973));
    defparam \pid_alt.error_p_reg_esr_1_LC_1_12_5 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_1_LC_1_12_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_1_LC_1_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_1_LC_1_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33181),
            .lcout(\pid_alt.error_p_regZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94314),
            .ce(N__34732),
            .sr(N__92976));
    defparam \pid_alt.error_i_reg_esr_2_LC_1_12_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_2_LC_1_12_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_2_LC_1_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_2_LC_1_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33295),
            .lcout(\pid_alt.error_i_regZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94314),
            .ce(N__34732),
            .sr(N__92976));
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_2_LC_1_13_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_2_LC_1_13_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_2_LC_1_13_0 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI0J511_2_LC_1_13_0  (
            .in0(N__33871),
            .in1(N__34039),
            .in2(_gnd_net_),
            .in3(N__34054),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI0J511Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_2_LC_1_13_1 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_2_LC_1_13_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_2_LC_1_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_2_LC_1_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33286),
            .lcout(\pid_alt.error_p_regZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94331),
            .ce(N__34733),
            .sr(N__92977));
    defparam \pid_alt.error_d_reg_esr_2_LC_1_13_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_2_LC_1_13_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_2_LC_1_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_2_LC_1_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33271),
            .lcout(\pid_alt.error_d_regZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94331),
            .ce(N__34733),
            .sr(N__92977));
    defparam \pid_alt.error_d_reg_prev_esr_RNI20IM_17_LC_1_13_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI20IM_17_LC_1_13_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI20IM_17_LC_1_13_3 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI20IM_17_LC_1_13_3  (
            .in0(N__33514),
            .in1(N__33949),
            .in2(_gnd_net_),
            .in3(N__33974),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI20IMZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI6P511_4_LC_1_13_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI6P511_4_LC_1_13_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI6P511_4_LC_1_13_6 .LUT_INIT=16'b1000100011101110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI6P511_4_LC_1_13_6  (
            .in0(N__35126),
            .in1(N__35163),
            .in2(_gnd_net_),
            .in3(N__35149),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI6P511Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_4_LC_1_13_7 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_4_LC_1_13_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_4_LC_1_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_4_LC_1_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33256),
            .lcout(\pid_alt.error_p_regZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94331),
            .ce(N__34733),
            .sr(N__92977));
    defparam \pid_alt.error_d_reg_prev_esr_RNICV511_6_LC_1_14_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNICV511_6_LC_1_14_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNICV511_6_LC_1_14_0 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNICV511_6_LC_1_14_0  (
            .in0(N__34998),
            .in1(N__34971),
            .in2(_gnd_net_),
            .in3(N__34956),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNICV511Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_RNIOI4P_0_LC_1_14_1 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNIOI4P_0_LC_1_14_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNIOI4P_0_LC_1_14_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pid_alt.error_p_reg_esr_RNIOI4P_0_LC_1_14_1  (
            .in0(_gnd_net_),
            .in1(N__33585),
            .in2(_gnd_net_),
            .in3(N__33353),
            .lcout(\pid_alt.error_p_reg_esr_RNIOI4PZ0Z_0 ),
            .ltout(\pid_alt.error_p_reg_esr_RNIOI4PZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIFPN33_1_LC_1_14_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIFPN33_1_LC_1_14_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIFPN33_1_LC_1_14_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIFPN33_1_LC_1_14_2  (
            .in0(N__38861),
            .in1(_gnd_net_),
            .in2(N__33358),
            .in3(N__33994),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIFPN33Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_6_LC_1_14_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_6_LC_1_14_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_6_LC_1_14_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_6_LC_1_14_3  (
            .in0(N__34957),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94346),
            .ce(N__40513),
            .sr(N__86494));
    defparam \pid_alt.error_d_reg_prev_esr_0_LC_1_14_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_0_LC_1_14_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_0_LC_1_14_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_0_LC_1_14_4  (
            .in0(N__33355),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94346),
            .ce(N__40513),
            .sr(N__86494));
    defparam \pid_alt.error_p_reg_esr_RNI3SMI1_0_LC_1_14_6 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNI3SMI1_0_LC_1_14_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNI3SMI1_0_LC_1_14_6 .LUT_INIT=16'b1010010110100101;
    LogicCell40 \pid_alt.error_p_reg_esr_RNI3SMI1_0_LC_1_14_6  (
            .in0(N__33354),
            .in1(_gnd_net_),
            .in2(N__33589),
            .in3(N__36762),
            .lcout(\pid_alt.error_p_reg_esr_RNI3SMI1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIMJHM_13_LC_1_14_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIMJHM_13_LC_1_14_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIMJHM_13_LC_1_14_7 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIMJHM_13_LC_1_14_7  (
            .in0(N__35202),
            .in1(N__35218),
            .in2(_gnd_net_),
            .in3(N__35240),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIMJHMZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_19_LC_1_15_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_19_LC_1_15_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_19_LC_1_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_19_LC_1_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33340),
            .lcout(\pid_front.error_p_regZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94361),
            .ce(N__93355),
            .sr(N__92978));
    defparam \pid_alt.error_i_reg_esr_1_LC_1_16_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_1_LC_1_16_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_1_LC_1_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_1_LC_1_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33331),
            .lcout(\pid_alt.error_i_regZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94369),
            .ce(N__34734),
            .sr(N__92979));
    defparam \pid_alt.error_i_reg_esr_4_LC_1_16_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_4_LC_1_16_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_4_LC_1_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_4_LC_1_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33319),
            .lcout(\pid_alt.error_i_regZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94369),
            .ce(N__34734),
            .sr(N__92979));
    defparam \pid_alt.error_i_reg_esr_5_LC_1_16_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_5_LC_1_16_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_5_LC_1_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_5_LC_1_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33307),
            .lcout(\pid_alt.error_i_regZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94369),
            .ce(N__34734),
            .sr(N__92979));
    defparam \pid_alt.error_d_reg_prev_esr_RNIGDHM_0_11_LC_1_17_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGDHM_0_11_LC_1_17_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGDHM_0_11_LC_1_17_1 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIGDHM_0_11_LC_1_17_1  (
            .in0(N__33687),
            .in1(N__33399),
            .in2(_gnd_net_),
            .in3(N__33389),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIGDHM_0Z0Z_11 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIGDHM_0Z0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI1FP62_10_LC_1_17_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI1FP62_10_LC_1_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI1FP62_10_LC_1_17_2 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI1FP62_10_LC_1_17_2  (
            .in0(_gnd_net_),
            .in1(N__33451),
            .in2(N__33454),
            .in3(N__34179),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI1FP62Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIDAHM_10_LC_1_17_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIDAHM_10_LC_1_17_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIDAHM_10_LC_1_17_3 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIDAHM_10_LC_1_17_3  (
            .in0(N__33661),
            .in1(N__33436),
            .in2(_gnd_net_),
            .in3(N__33421),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIDAHMZ0Z_10 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIDAHMZ0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNITPKD4_10_LC_1_17_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNITPKD4_10_LC_1_17_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNITPKD4_10_LC_1_17_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNITPKD4_10_LC_1_17_4  (
            .in0(N__33445),
            .in1(N__37299),
            .in2(N__33439),
            .in3(N__34178),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNITPKD4Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIDAHM_0_10_LC_1_17_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIDAHM_0_10_LC_1_17_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIDAHM_0_10_LC_1_17_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIDAHM_0_10_LC_1_17_5  (
            .in0(N__33660),
            .in1(N__33435),
            .in2(_gnd_net_),
            .in3(N__33420),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIDAHM_0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_11_LC_1_17_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_11_LC_1_17_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_11_LC_1_17_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_11_LC_1_17_6  (
            .in0(N__33391),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94377),
            .ce(N__40506),
            .sr(N__86476));
    defparam \pid_alt.error_d_reg_prev_esr_RNIGDHM_11_LC_1_17_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGDHM_11_LC_1_17_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGDHM_11_LC_1_17_7 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIGDHM_11_LC_1_17_7  (
            .in0(N__33688),
            .in1(N__33400),
            .in2(_gnd_net_),
            .in3(N__33390),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIGDHMZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNICG9B1_20_LC_1_18_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNICG9B1_20_LC_1_18_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNICG9B1_20_LC_1_18_0 .LUT_INIT=16'b1111110101000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNICG9B1_20_LC_1_18_0  (
            .in0(N__35816),
            .in1(N__35777),
            .in2(N__35734),
            .in3(N__35686),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNICG9B1Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNICG9B1_2_20_LC_1_18_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNICG9B1_2_20_LC_1_18_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNICG9B1_2_20_LC_1_18_2 .LUT_INIT=16'b0100001010111101;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNICG9B1_2_20_LC_1_18_2  (
            .in0(N__35817),
            .in1(N__35778),
            .in2(N__35735),
            .in3(N__35687),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNICG9B1_2Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_20_LC_1_18_3 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_20_LC_1_18_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_20_LC_1_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_20_LC_1_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33373),
            .lcout(\pid_alt.error_p_regZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94385),
            .ce(N__34735),
            .sr(N__92983));
    defparam \pid_alt.error_d_reg_prev_esr_RNIL8611_9_LC_1_18_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIL8611_9_LC_1_18_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIL8611_9_LC_1_18_4 .LUT_INIT=16'b1101110101000100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIL8611_9_LC_1_18_4  (
            .in0(N__37612),
            .in1(N__37698),
            .in2(_gnd_net_),
            .in3(N__37636),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIL8611Z0Z_9 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIL8611Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNICI045_9_LC_1_18_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNICI045_9_LC_1_18_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNICI045_9_LC_1_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNICI045_9_LC_1_18_5  (
            .in0(N__37669),
            .in1(N__33483),
            .in2(N__33493),
            .in3(N__35654),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNICI045Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNO_0_24_LC_1_18_6 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNO_0_24_LC_1_18_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNO_0_24_LC_1_18_6 .LUT_INIT=16'b1011111111111101;
    LogicCell40 \pid_alt.pid_prereg_esr_RNO_0_24_LC_1_18_6  (
            .in0(N__35818),
            .in1(N__35779),
            .in2(N__35736),
            .in3(N__35688),
            .lcout(\pid_alt.un1_pid_prereg_0_axb_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNISAR62_9_LC_1_18_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNISAR62_9_LC_1_18_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNISAR62_9_LC_1_18_7 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNISAR62_9_LC_1_18_7  (
            .in0(N__33490),
            .in1(N__33484),
            .in2(_gnd_net_),
            .in3(N__35655),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNISAR62Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI8DL14_16_LC_1_19_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI8DL14_16_LC_1_19_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI8DL14_16_LC_1_19_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI8DL14_16_LC_1_19_0  (
            .in0(N__33475),
            .in1(N__36197),
            .in2(N__37122),
            .in3(N__33465),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI8DL14Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI20IM_0_17_LC_1_19_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI20IM_0_17_LC_1_19_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI20IM_0_17_LC_1_19_1 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI20IM_0_17_LC_1_19_1  (
            .in0(N__33978),
            .in1(_gnd_net_),
            .in2(N__33948),
            .in3(N__33507),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI20IM_0Z0Z_17 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNI20IM_0Z0Z_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI8BR02_16_LC_1_19_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI8BR02_16_LC_1_19_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI8BR02_16_LC_1_19_2 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI8BR02_16_LC_1_19_2  (
            .in0(_gnd_net_),
            .in1(N__36198),
            .in2(N__33469),
            .in3(N__33466),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI8BR02Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIVSHM_16_LC_1_19_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIVSHM_16_LC_1_19_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIVSHM_16_LC_1_19_3 .LUT_INIT=16'b1101110101000100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIVSHM_16_LC_1_19_3  (
            .in0(N__33607),
            .in1(N__33844),
            .in2(_gnd_net_),
            .in3(N__33628),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIVSHMZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIVSHM_0_16_LC_1_19_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIVSHM_0_16_LC_1_19_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIVSHM_0_16_LC_1_19_4 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIVSHM_0_16_LC_1_19_4  (
            .in0(N__33843),
            .in1(N__33606),
            .in2(_gnd_net_),
            .in3(N__33626),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI02Q02_15_LC_1_19_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI02Q02_15_LC_1_19_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI02Q02_15_LC_1_19_5 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI02Q02_15_LC_1_19_5  (
            .in0(_gnd_net_),
            .in1(N__34566),
            .in2(N__33457),
            .in3(N__40267),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI02Q02Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_16_LC_1_19_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_16_LC_1_19_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_16_LC_1_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_16_LC_1_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33627),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94390),
            .ce(N__40501),
            .sr(N__86463));
    defparam \pid_alt.error_p_reg_esr_0_LC_1_21_0 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_0_LC_1_21_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_0_LC_1_21_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_0_LC_1_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33598),
            .lcout(\pid_alt.error_p_regZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94400),
            .ce(N__34736),
            .sr(N__92988));
    defparam \pid_alt.error_p_reg_esr_6_LC_1_21_4 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_6_LC_1_21_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_6_LC_1_21_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_6_LC_1_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33574),
            .lcout(\pid_alt.error_p_regZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94400),
            .ce(N__34736),
            .sr(N__92988));
    defparam \pid_alt.error_p_reg_esr_18_LC_1_22_0 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_18_LC_1_22_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_18_LC_1_22_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_18_LC_1_22_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33565),
            .lcout(\pid_alt.error_p_regZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94405),
            .ce(N__34737),
            .sr(N__92991));
    defparam \pid_alt.error_p_reg_esr_19_LC_1_22_1 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_19_LC_1_22_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_19_LC_1_22_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_19_LC_1_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33553),
            .lcout(\pid_alt.error_p_regZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94405),
            .ce(N__34737),
            .sr(N__92991));
    defparam \pid_alt.error_p_reg_esr_13_LC_1_22_2 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_13_LC_1_22_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_13_LC_1_22_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_p_reg_esr_13_LC_1_22_2  (
            .in0(N__33541),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_p_regZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94405),
            .ce(N__34737),
            .sr(N__92991));
    defparam \pid_alt.error_p_reg_esr_5_LC_1_22_3 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_5_LC_1_22_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_5_LC_1_22_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_p_reg_esr_5_LC_1_22_3  (
            .in0(N__33532),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_p_regZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94405),
            .ce(N__34737),
            .sr(N__92991));
    defparam \pid_alt.error_p_reg_esr_17_LC_1_22_4 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_17_LC_1_22_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_17_LC_1_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_17_LC_1_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33523),
            .lcout(\pid_alt.error_p_regZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94405),
            .ce(N__34737),
            .sr(N__92991));
    defparam \pid_alt.error_p_reg_esr_7_LC_1_22_5 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_7_LC_1_22_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_7_LC_1_22_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_7_LC_1_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33727),
            .lcout(\pid_alt.error_p_regZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94405),
            .ce(N__34737),
            .sr(N__92991));
    defparam \pid_alt.error_p_reg_esr_8_LC_1_22_6 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_8_LC_1_22_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_8_LC_1_22_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_8_LC_1_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33718),
            .lcout(\pid_alt.error_p_regZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94405),
            .ce(N__34737),
            .sr(N__92991));
    defparam \pid_alt.error_p_reg_esr_9_LC_1_22_7 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_9_LC_1_22_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_9_LC_1_22_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_9_LC_1_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33709),
            .lcout(\pid_alt.error_p_regZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94405),
            .ce(N__34737),
            .sr(N__92991));
    defparam \pid_alt.error_p_reg_esr_3_LC_1_23_1 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_3_LC_1_23_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_3_LC_1_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_3_LC_1_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33700),
            .lcout(\pid_alt.error_p_regZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94409),
            .ce(N__34738),
            .sr(N__92995));
    defparam \pid_alt.error_p_reg_esr_11_LC_1_23_2 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_11_LC_1_23_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_11_LC_1_23_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_p_reg_esr_11_LC_1_23_2  (
            .in0(N__33694),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_p_regZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94409),
            .ce(N__34738),
            .sr(N__92995));
    defparam \pid_alt.error_p_reg_esr_12_LC_1_23_3 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_12_LC_1_23_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_12_LC_1_23_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_p_reg_esr_12_LC_1_23_3  (
            .in0(N__33676),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_p_regZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94409),
            .ce(N__34738),
            .sr(N__92995));
    defparam \pid_alt.error_p_reg_esr_10_LC_1_23_4 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_10_LC_1_23_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_10_LC_1_23_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_10_LC_1_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33667),
            .lcout(\pid_alt.error_p_regZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94409),
            .ce(N__34738),
            .sr(N__92995));
    defparam \pid_alt.error_p_reg_esr_14_LC_1_23_5 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_14_LC_1_23_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_14_LC_1_23_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_14_LC_1_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33646),
            .lcout(\pid_alt.error_p_regZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94409),
            .ce(N__34738),
            .sr(N__92995));
    defparam \pid_alt.error_p_reg_esr_15_LC_1_23_6 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_15_LC_1_23_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_15_LC_1_23_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_15_LC_1_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33637),
            .lcout(\pid_alt.error_p_regZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94409),
            .ce(N__34738),
            .sr(N__92995));
    defparam \pid_alt.error_p_reg_esr_16_LC_1_23_7 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_16_LC_1_23_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_16_LC_1_23_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_16_LC_1_23_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33853),
            .lcout(\pid_alt.error_p_regZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94409),
            .ce(N__34738),
            .sr(N__92995));
    defparam \pid_alt.error_d_reg_esr_1_LC_2_5_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_1_LC_2_5_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_1_LC_2_5_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_1_LC_2_5_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33832),
            .lcout(\pid_alt.error_d_regZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94188),
            .ce(N__34724),
            .sr(N__92966));
    defparam \Commands_frame_decoder.source_alt_kd_0_LC_2_9_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kd_0_LC_2_9_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kd_0_LC_2_9_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kd_0_LC_2_9_0  (
            .in0(_gnd_net_),
            .in1(N__88280),
            .in2(_gnd_net_),
            .in3(N__93126),
            .lcout(alt_kd_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94253),
            .ce(N__51607),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kd_1_LC_2_9_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kd_1_LC_2_9_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kd_1_LC_2_9_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_kd_1_LC_2_9_1  (
            .in0(N__93127),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85526),
            .lcout(alt_kd_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94253),
            .ce(N__51607),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kd_2_LC_2_9_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kd_2_LC_2_9_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kd_2_LC_2_9_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kd_2_LC_2_9_2  (
            .in0(_gnd_net_),
            .in1(N__92521),
            .in2(_gnd_net_),
            .in3(N__93128),
            .lcout(alt_kd_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94253),
            .ce(N__51607),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kd_3_LC_2_9_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kd_3_LC_2_9_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kd_3_LC_2_9_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_kd_3_LC_2_9_3  (
            .in0(N__93129),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__92326),
            .lcout(alt_kd_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94253),
            .ce(N__51607),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kd_4_LC_2_9_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kd_4_LC_2_9_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kd_4_LC_2_9_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kd_4_LC_2_9_4  (
            .in0(_gnd_net_),
            .in1(N__88861),
            .in2(_gnd_net_),
            .in3(N__93130),
            .lcout(alt_kd_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94253),
            .ce(N__51607),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kd_5_LC_2_9_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kd_5_LC_2_9_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kd_5_LC_2_9_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_kd_5_LC_2_9_5  (
            .in0(N__93131),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88695),
            .lcout(alt_kd_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94253),
            .ce(N__51607),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kd_6_LC_2_9_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kd_6_LC_2_9_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kd_6_LC_2_9_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kd_6_LC_2_9_6  (
            .in0(_gnd_net_),
            .in1(N__88506),
            .in2(_gnd_net_),
            .in3(N__93132),
            .lcout(alt_kd_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94253),
            .ce(N__51607),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kd_7_LC_2_9_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kd_7_LC_2_9_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kd_7_LC_2_9_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_kd_7_LC_2_9_7  (
            .in0(N__93133),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__92127),
            .lcout(alt_kd_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94253),
            .ce(N__51607),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_8_LC_2_10_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_8_LC_2_10_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_8_LC_2_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_8_LC_2_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33925),
            .lcout(\pid_alt.error_i_regZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94271),
            .ce(N__34729),
            .sr(N__92971));
    defparam \pid_alt.error_i_reg_esr_10_LC_2_10_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_10_LC_2_10_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_10_LC_2_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_10_LC_2_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33913),
            .lcout(\pid_alt.error_i_regZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94271),
            .ce(N__34729),
            .sr(N__92971));
    defparam \pid_alt.error_i_reg_esr_0_LC_2_10_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_0_LC_2_10_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_0_LC_2_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_0_LC_2_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33901),
            .lcout(\pid_alt.error_i_regZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94271),
            .ce(N__34729),
            .sr(N__92971));
    defparam \Commands_frame_decoder.source_alt_ki_5_LC_2_11_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_5_LC_2_11_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_5_LC_2_11_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_5_LC_2_11_3  (
            .in0(_gnd_net_),
            .in1(N__88702),
            .in2(_gnd_net_),
            .in3(N__93140),
            .lcout(alt_ki_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94287),
            .ce(N__42735),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_ki_6_LC_2_11_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_6_LC_2_11_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_6_LC_2_11_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_6_LC_2_11_4  (
            .in0(N__93141),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88509),
            .lcout(alt_ki_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94287),
            .ce(N__42735),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_1_LC_2_12_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_1_LC_2_12_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_1_LC_2_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_1_LC_2_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34087),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94301),
            .ce(N__40515),
            .sr(N__86501));
    defparam \pid_alt.error_d_reg_prev_esr_18_LC_2_12_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_18_LC_2_12_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_18_LC_2_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_18_LC_2_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35579),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94301),
            .ce(N__40515),
            .sr(N__86501));
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_0_2_LC_2_13_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_0_2_LC_2_13_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_0_2_LC_2_13_0 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI0J511_0_2_LC_2_13_0  (
            .in0(N__33870),
            .in1(N__34038),
            .in2(_gnd_net_),
            .in3(N__34052),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI0J511_0Z0Z_2 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNI0J511_0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIT2B22_1_LC_2_13_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIT2B22_1_LC_2_13_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIT2B22_1_LC_2_13_1 .LUT_INIT=16'b0100101111010010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIT2B22_1_LC_2_13_1  (
            .in0(N__34114),
            .in1(N__34101),
            .in2(N__33856),
            .in3(N__34086),
            .lcout(\pid_alt.un1_pid_prereg_16_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNITF511_1_LC_2_13_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNITF511_1_LC_2_13_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNITF511_1_LC_2_13_2 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNITF511_1_LC_2_13_2  (
            .in0(N__34085),
            .in1(_gnd_net_),
            .in2(N__34102),
            .in3(N__34113),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNITF511Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNITF511_0_1_LC_2_13_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNITF511_0_1_LC_2_13_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNITF511_0_1_LC_2_13_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNITF511_0_1_LC_2_13_5  (
            .in0(N__34112),
            .in1(N__34097),
            .in2(_gnd_net_),
            .in3(N__34084),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNITF511_0Z0Z_1 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNITF511_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIF0465_1_LC_2_13_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIF0465_1_LC_2_13_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIF0465_1_LC_2_13_6 .LUT_INIT=16'b0011110011001100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIF0465_1_LC_2_13_6  (
            .in0(N__37071),
            .in1(N__34063),
            .in2(N__34057),
            .in3(N__34015),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIF0465Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_2_LC_2_13_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_2_LC_2_13_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_2_LC_2_13_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_2_LC_2_13_7  (
            .in0(N__34053),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94319),
            .ce(N__40514),
            .sr(N__86495));
    defparam \pid_alt.error_d_reg_prev_esr_RNI2Q08_0_LC_2_14_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI2Q08_0_LC_2_14_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI2Q08_0_LC_2_14_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI2Q08_0_LC_2_14_3  (
            .in0(N__34027),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prev_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNII5LS3_1_LC_2_14_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNII5LS3_1_LC_2_14_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNII5LS3_1_LC_2_14_6 .LUT_INIT=16'b1110100010100000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNII5LS3_1_LC_2_14_6  (
            .in0(N__34021),
            .in1(N__34014),
            .in2(N__34003),
            .in3(N__33993),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNII5LS3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI3M511_0_3_LC_2_14_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI3M511_0_3_LC_2_14_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI3M511_0_3_LC_2_14_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI3M511_0_3_LC_2_14_7  (
            .in0(N__34842),
            .in1(N__35055),
            .in2(_gnd_net_),
            .in3(N__35087),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI3M511_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_13_LC_2_15_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_13_LC_2_15_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_13_LC_2_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_13_LC_2_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35242),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94349),
            .ce(N__40509),
            .sr(N__86483));
    defparam \pid_alt.error_d_reg_prev_esr_17_LC_2_15_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_17_LC_2_15_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_17_LC_2_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_17_LC_2_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33982),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94349),
            .ce(N__40509),
            .sr(N__86483));
    defparam \pid_alt.error_d_reg_prev_esr_4_LC_2_15_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_4_LC_2_15_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_4_LC_2_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_4_LC_2_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35131),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94349),
            .ce(N__40509),
            .sr(N__86483));
    defparam \pid_alt.error_i_acumm_prereg_esr_16_LC_2_15_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_16_LC_2_15_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_16_LC_2_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_16_LC_2_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34570),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94349),
            .ce(N__40509),
            .sr(N__86483));
    defparam \pid_alt.error_i_acumm_prereg_esr_21_LC_2_15_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_21_LC_2_15_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_21_LC_2_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_21_LC_2_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35692),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94349),
            .ce(N__40509),
            .sr(N__86483));
    defparam \pid_alt.error_i_acumm_prereg_esr_18_LC_2_15_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_18_LC_2_15_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_18_LC_2_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_18_LC_2_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35482),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94349),
            .ce(N__40509),
            .sr(N__86483));
    defparam \pid_alt.error_i_acumm_prereg_esr_11_LC_2_15_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_11_LC_2_15_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_11_LC_2_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_11_LC_2_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34183),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94349),
            .ce(N__40509),
            .sr(N__86483));
    defparam \pid_alt.error_i_acumm_esr_RNIB9IP_0_LC_2_16_0 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_esr_RNIB9IP_0_LC_2_16_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_esr_RNIB9IP_0_LC_2_16_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pid_alt.error_i_acumm_esr_RNIB9IP_0_LC_2_16_0  (
            .in0(_gnd_net_),
            .in1(N__38742),
            .in2(N__38772),
            .in3(_gnd_net_),
            .lcout(\pid_alt.un1_pid_prereg_0 ),
            .ltout(),
            .carryin(bfn_2_16_0_),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_RNIQMD91_1_LC_2_16_1 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_esr_RNIQMD91_1_LC_2_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_esr_RNIQMD91_1_LC_2_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_acumm_esr_RNIQMD91_1_LC_2_16_1  (
            .in0(_gnd_net_),
            .in1(N__34639),
            .in2(N__34162),
            .in3(N__34153),
            .lcout(\pid_alt.error_i_acumm_esr_RNIQMD91Z0Z_1 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_0 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_RNITQE91_2_LC_2_16_2 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_esr_RNITQE91_2_LC_2_16_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_esr_RNITQE91_2_LC_2_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_acumm_esr_RNITQE91_2_LC_2_16_2  (
            .in0(_gnd_net_),
            .in1(N__34630),
            .in2(N__34150),
            .in3(N__34135),
            .lcout(\pid_alt.error_i_acumm_esr_RNITQE91Z0Z_2 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_1 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_RNI0VF91_3_LC_2_16_3 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_esr_RNI0VF91_3_LC_2_16_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_esr_RNI0VF91_3_LC_2_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_acumm_esr_RNI0VF91_3_LC_2_16_3  (
            .in0(_gnd_net_),
            .in1(N__34648),
            .in2(N__34132),
            .in3(N__34117),
            .lcout(\pid_alt.error_i_acumm_esr_RNI0VF91Z0Z_3 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_2 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_RNI33H91_4_LC_2_16_4 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_esr_RNI33H91_4_LC_2_16_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_esr_RNI33H91_4_LC_2_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_acumm_esr_RNI33H91_4_LC_2_16_4  (
            .in0(_gnd_net_),
            .in1(N__34813),
            .in2(N__34312),
            .in3(N__34303),
            .lcout(\pid_alt.error_i_acumm_esr_RNI33H91Z0Z_4 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_3 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_RNIT8KA1_5_LC_2_16_5 .C_ON=1'b1;
    defparam \pid_alt.error_i_reg_esr_RNIT8KA1_5_LC_2_16_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_reg_esr_RNIT8KA1_5_LC_2_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_reg_esr_RNIT8KA1_5_LC_2_16_5  (
            .in0(_gnd_net_),
            .in1(N__34666),
            .in2(N__34300),
            .in3(N__34291),
            .lcout(\pid_alt.error_i_reg_esr_RNIT8KA1Z0Z_5 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_4 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ_LC_2_16_6 .C_ON=1'b1;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ_LC_2_16_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ_LC_2_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ_LC_2_16_6  (
            .in0(_gnd_net_),
            .in1(N__34519),
            .in2(N__34288),
            .in3(N__34273),
            .lcout(\pid_alt.un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_5 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ_LC_2_16_7 .C_ON=1'b1;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ_LC_2_16_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ_LC_2_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ_LC_2_16_7  (
            .in0(_gnd_net_),
            .in1(N__34504),
            .in2(N__34270),
            .in3(N__34255),
            .lcout(\pid_alt.un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_6 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ_LC_2_17_0 .C_ON=1'b1;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ_LC_2_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ_LC_2_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ_LC_2_17_0  (
            .in0(_gnd_net_),
            .in1(N__34489),
            .in2(N__34252),
            .in3(N__34237),
            .lcout(\pid_alt.un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ ),
            .ltout(),
            .carryin(bfn_2_17_0_),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_8_c_RNI9POQ_LC_2_17_1 .C_ON=1'b1;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_8_c_RNI9POQ_LC_2_17_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_8_c_RNI9POQ_LC_2_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_8_c_RNI9POQ_LC_2_17_1  (
            .in0(_gnd_net_),
            .in1(N__34473),
            .in2(N__34234),
            .in3(N__34216),
            .lcout(\pid_alt.un1_error_i_acumm_prereg_cry_8_c_RNI9POQ ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_8 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_9_c_RNIQN3F_LC_2_17_2 .C_ON=1'b1;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_9_c_RNIQN3F_LC_2_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_9_c_RNIQN3F_LC_2_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_9_c_RNIQN3F_LC_2_17_2  (
            .in0(_gnd_net_),
            .in1(N__34549),
            .in2(N__34213),
            .in3(N__34201),
            .lcout(\pid_alt.un1_error_i_acumm_prereg_cry_9_c_RNIQN3F ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_9 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_RNI4NMP_11_LC_2_17_3 .C_ON=1'b1;
    defparam \pid_alt.error_i_reg_esr_RNI4NMP_11_LC_2_17_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_reg_esr_RNI4NMP_11_LC_2_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_reg_esr_RNI4NMP_11_LC_2_17_3  (
            .in0(_gnd_net_),
            .in1(N__34534),
            .in2(N__34198),
            .in3(N__34165),
            .lcout(\pid_alt.error_i_reg_esr_RNI4NMPZ0Z_11 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_10 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_RNI7RNP_12_LC_2_17_4 .C_ON=1'b1;
    defparam \pid_alt.error_i_reg_esr_RNI7RNP_12_LC_2_17_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_reg_esr_RNI7RNP_12_LC_2_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_reg_esr_RNI7RNP_12_LC_2_17_4  (
            .in0(_gnd_net_),
            .in1(N__34459),
            .in2(N__34684),
            .in3(N__34444),
            .lcout(\pid_alt.error_i_reg_esr_RNI7RNPZ0Z_12 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_11 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_RNIJ6LM_13_LC_2_17_5 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_esr_RNIJ6LM_13_LC_2_17_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_esr_RNIJ6LM_13_LC_2_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_acumm_esr_RNIJ6LM_13_LC_2_17_5  (
            .in0(_gnd_net_),
            .in1(N__57544),
            .in2(N__34441),
            .in3(N__34426),
            .lcout(\pid_alt.error_i_acumm_esr_RNIJ6LMZ0Z_13 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_12 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_RNI15KJ_14_LC_2_17_6 .C_ON=1'b1;
    defparam \pid_alt.error_i_reg_esr_RNI15KJ_14_LC_2_17_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_reg_esr_RNI15KJ_14_LC_2_17_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_i_reg_esr_RNI15KJ_14_LC_2_17_6  (
            .in0(_gnd_net_),
            .in1(N__34423),
            .in2(_gnd_net_),
            .in3(N__34408),
            .lcout(\pid_alt.error_i_reg_esr_RNI15KJZ0Z_14 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_13 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_RNI38LJ_15_LC_2_17_7 .C_ON=1'b1;
    defparam \pid_alt.error_i_reg_esr_RNI38LJ_15_LC_2_17_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_reg_esr_RNI38LJ_15_LC_2_17_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_i_reg_esr_RNI38LJ_15_LC_2_17_7  (
            .in0(_gnd_net_),
            .in1(N__34405),
            .in2(_gnd_net_),
            .in3(N__34390),
            .lcout(\pid_alt.error_i_reg_esr_RNI38LJZ0Z_15 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_14 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_RNI5BMJ_16_LC_2_18_0 .C_ON=1'b1;
    defparam \pid_alt.error_i_reg_esr_RNI5BMJ_16_LC_2_18_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_reg_esr_RNI5BMJ_16_LC_2_18_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_i_reg_esr_RNI5BMJ_16_LC_2_18_0  (
            .in0(_gnd_net_),
            .in1(N__34387),
            .in2(_gnd_net_),
            .in3(N__34372),
            .lcout(\pid_alt.error_i_reg_esr_RNI5BMJZ0Z_16 ),
            .ltout(),
            .carryin(bfn_2_18_0_),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_RNI7ENJ_17_LC_2_18_1 .C_ON=1'b1;
    defparam \pid_alt.error_i_reg_esr_RNI7ENJ_17_LC_2_18_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_reg_esr_RNI7ENJ_17_LC_2_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_i_reg_esr_RNI7ENJ_17_LC_2_18_1  (
            .in0(_gnd_net_),
            .in1(N__34369),
            .in2(_gnd_net_),
            .in3(N__34354),
            .lcout(\pid_alt.error_i_reg_esr_RNI7ENJZ0Z_17 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_16 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_RNI9HOJ_18_LC_2_18_2 .C_ON=1'b1;
    defparam \pid_alt.error_i_reg_esr_RNI9HOJ_18_LC_2_18_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_reg_esr_RNI9HOJ_18_LC_2_18_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_i_reg_esr_RNI9HOJ_18_LC_2_18_2  (
            .in0(_gnd_net_),
            .in1(N__34351),
            .in2(_gnd_net_),
            .in3(N__34336),
            .lcout(\pid_alt.error_i_reg_esr_RNI9HOJZ0Z_18 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_17 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_RNIBKPJ_19_LC_2_18_3 .C_ON=1'b1;
    defparam \pid_alt.error_i_reg_esr_RNIBKPJ_19_LC_2_18_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_reg_esr_RNIBKPJ_19_LC_2_18_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_i_reg_esr_RNIBKPJ_19_LC_2_18_3  (
            .in0(_gnd_net_),
            .in1(N__34333),
            .in2(_gnd_net_),
            .in3(N__34318),
            .lcout(\pid_alt.error_i_reg_esr_RNIBKPJZ0Z_19 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_18 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ_LC_2_18_4 .C_ON=1'b1;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ_LC_2_18_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ_LC_2_18_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ_LC_2_18_4  (
            .in0(_gnd_net_),
            .in1(N__34596),
            .in2(_gnd_net_),
            .in3(N__34315),
            .lcout(\pid_alt.un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_19 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_20_c_RNISVKK_LC_2_18_5 .C_ON=1'b0;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_20_c_RNISVKK_LC_2_18_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_20_c_RNISVKK_LC_2_18_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_20_c_RNISVKK_LC_2_18_5  (
            .in0(N__34597),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34579),
            .lcout(\pid_alt.un1_error_i_acumm_prereg_cry_20_c_RNISVKK ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIOQI14_15_LC_2_18_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOQI14_15_LC_2_18_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOQI14_15_LC_2_18_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIOQI14_15_LC_2_18_6  (
            .in0(N__34576),
            .in1(N__40263),
            .in2(N__37150),
            .in3(N__34565),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIOQI14Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNICG9B1_0_20_LC_2_18_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNICG9B1_0_20_LC_2_18_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNICG9B1_0_20_LC_2_18_7 .LUT_INIT=16'b0100001010111101;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNICG9B1_0_20_LC_2_18_7  (
            .in0(N__35808),
            .in1(N__35776),
            .in2(N__35733),
            .in3(N__35684),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNICG9B1_0Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_10_LC_2_19_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_10_LC_2_19_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_10_LC_2_19_0 .LUT_INIT=16'b1110111000101110;
    LogicCell40 \pid_alt.error_i_acumm_10_LC_2_19_0  (
            .in0(N__34548),
            .in1(N__69014),
            .in2(N__35975),
            .in3(N__36097),
            .lcout(\pid_alt.error_i_acummZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94388),
            .ce(),
            .sr(N__57489));
    defparam \pid_alt.error_i_acumm_11_LC_2_19_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_11_LC_2_19_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_11_LC_2_19_1 .LUT_INIT=16'b1011111110110000;
    LogicCell40 \pid_alt.error_i_acumm_11_LC_2_19_1  (
            .in0(N__38081),
            .in1(N__35965),
            .in2(N__69025),
            .in3(N__34533),
            .lcout(\pid_alt.error_i_acummZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94388),
            .ce(),
            .sr(N__57489));
    defparam \pid_alt.error_i_acumm_6_LC_2_19_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_6_LC_2_19_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_6_LC_2_19_2 .LUT_INIT=16'b1110111000101110;
    LogicCell40 \pid_alt.error_i_acumm_6_LC_2_19_2  (
            .in0(N__34518),
            .in1(N__69020),
            .in2(N__35976),
            .in3(N__38686),
            .lcout(\pid_alt.error_i_acummZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94388),
            .ce(),
            .sr(N__57489));
    defparam \pid_alt.error_i_acumm_7_LC_2_19_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_7_LC_2_19_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_7_LC_2_19_3 .LUT_INIT=16'b1111011110100010;
    LogicCell40 \pid_alt.error_i_acumm_7_LC_2_19_3  (
            .in0(N__69021),
            .in1(N__35969),
            .in2(N__38710),
            .in3(N__34503),
            .lcout(\pid_alt.error_i_acummZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94388),
            .ce(),
            .sr(N__57489));
    defparam \pid_alt.error_i_acumm_8_LC_2_19_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_8_LC_2_19_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_8_LC_2_19_4 .LUT_INIT=16'b1110111000101110;
    LogicCell40 \pid_alt.error_i_acumm_8_LC_2_19_4  (
            .in0(N__34488),
            .in1(N__69022),
            .in2(N__35977),
            .in3(N__38106),
            .lcout(\pid_alt.error_i_acummZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94388),
            .ce(),
            .sr(N__57489));
    defparam \pid_alt.error_i_acumm_9_LC_2_19_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_9_LC_2_19_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_9_LC_2_19_5 .LUT_INIT=16'b1110010011101110;
    LogicCell40 \pid_alt.error_i_acumm_9_LC_2_19_5  (
            .in0(N__69023),
            .in1(N__34474),
            .in2(N__38137),
            .in3(N__35973),
            .lcout(\pid_alt.error_i_acummZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94388),
            .ce(),
            .sr(N__57489));
    defparam \pid_alt.error_i_acumm_12_LC_2_19_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_12_LC_2_19_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_12_LC_2_19_6 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \pid_alt.error_i_acumm_12_LC_2_19_6  (
            .in0(N__34680),
            .in1(N__69018),
            .in2(N__35926),
            .in3(N__35995),
            .lcout(\pid_alt.error_i_acummZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94388),
            .ce(),
            .sr(N__57489));
    defparam \pid_alt.error_i_acumm_5_LC_2_19_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_5_LC_2_19_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_5_LC_2_19_7 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \pid_alt.error_i_acumm_5_LC_2_19_7  (
            .in0(N__69019),
            .in1(N__36026),
            .in2(N__38616),
            .in3(N__34662),
            .lcout(\pid_alt.error_i_acummZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94388),
            .ce(),
            .sr(N__57489));
    defparam \pid_alt.error_i_acumm_esr_3_LC_2_20_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_esr_3_LC_2_20_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_esr_3_LC_2_20_0 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \pid_alt.error_i_acumm_esr_3_LC_2_20_0  (
            .in0(N__38809),
            .in1(N__36025),
            .in2(N__36064),
            .in3(N__34612),
            .lcout(\pid_alt.error_i_acummZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94394),
            .ce(N__57509),
            .sr(N__57478));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNICB6L2_5_LC_2_20_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNICB6L2_5_LC_2_20_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNICB6L2_5_LC_2_20_1 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNICB6L2_5_LC_2_20_1  (
            .in0(N__38658),
            .in1(N__36044),
            .in2(N__38615),
            .in3(N__35920),
            .lcout(\pid_alt.error_i_acumm_prereg_esr_RNICB6L2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_1_LC_2_20_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_esr_1_LC_2_20_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_esr_1_LC_2_20_2 .LUT_INIT=16'b1110000001000000;
    LogicCell40 \pid_alt.error_i_acumm_esr_1_LC_2_20_2  (
            .in0(N__38807),
            .in1(N__34610),
            .in2(N__38830),
            .in3(N__36021),
            .lcout(\pid_alt.error_i_acummZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94394),
            .ce(N__57509),
            .sr(N__57478));
    defparam \pid_alt.error_i_acumm_esr_2_LC_2_20_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_esr_2_LC_2_20_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_esr_2_LC_2_20_3 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \pid_alt.error_i_acumm_esr_2_LC_2_20_3  (
            .in0(N__34611),
            .in1(N__36079),
            .in2(N__36028),
            .in3(N__38808),
            .lcout(\pid_alt.error_i_acummZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94394),
            .ce(N__57509),
            .sr(N__57478));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNICB6L2_0_5_LC_2_20_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNICB6L2_0_5_LC_2_20_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNICB6L2_0_5_LC_2_20_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNICB6L2_0_5_LC_2_20_4  (
            .in0(N__35921),
            .in1(N__36045),
            .in2(N__38608),
            .in3(N__38659),
            .lcout(),
            .ltout(\pid_alt.error_i_acumm_prereg_esr_RNICB6L2_0Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIPTHL5_5_LC_2_20_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIPTHL5_5_LC_2_20_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIPTHL5_5_LC_2_20_5 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNIPTHL5_5_LC_2_20_5  (
            .in0(_gnd_net_),
            .in1(N__35961),
            .in2(N__34621),
            .in3(N__34618),
            .lcout(\pid_alt.N_159 ),
            .ltout(\pid_alt.N_159_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_0_LC_2_20_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_esr_0_LC_2_20_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_esr_0_LC_2_20_6 .LUT_INIT=16'b1101100000000000;
    LogicCell40 \pid_alt.error_i_acumm_esr_0_LC_2_20_6  (
            .in0(N__38806),
            .in1(N__36020),
            .in2(N__34600),
            .in3(N__38725),
            .lcout(\pid_alt.error_i_acummZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94394),
            .ce(N__57509),
            .sr(N__57478));
    defparam \pid_alt.error_i_acumm_esr_4_LC_2_21_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_esr_4_LC_2_21_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_esr_4_LC_2_21_5 .LUT_INIT=16'b1111111100110101;
    LogicCell40 \pid_alt.error_i_acumm_esr_4_LC_2_21_5  (
            .in0(N__35974),
            .in1(N__36027),
            .in2(N__38617),
            .in3(N__38805),
            .lcout(\pid_alt.error_i_acummZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94397),
            .ce(N__57516),
            .sr(N__57485));
    defparam \Commands_frame_decoder.source_alt_kp_e_0_5_LC_2_22_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_5_LC_2_22_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_5_LC_2_22_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_e_0_5_LC_2_22_0  (
            .in0(N__88480),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__93154),
            .lcout(alt_kp_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94403),
            .ce(N__48701),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kp_e_0_1_LC_2_23_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_1_LC_2_23_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_1_LC_2_23_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_e_0_1_LC_2_23_2  (
            .in0(_gnd_net_),
            .in1(N__85489),
            .in2(_gnd_net_),
            .in3(N__93155),
            .lcout(alt_kp_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94408),
            .ce(N__48709),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kp_e_0_3_LC_2_23_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_3_LC_2_23_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_3_LC_2_23_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_e_0_3_LC_2_23_3  (
            .in0(N__93156),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__92331),
            .lcout(alt_kp_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94408),
            .ce(N__48709),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_5_LC_2_26_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_5_LC_2_26_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_5_LC_2_26_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_5_LC_2_26_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34768),
            .lcout(\pid_front.error_p_regZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94411),
            .ce(N__93409),
            .sr(N__92999));
    defparam \pid_alt.error_d_reg_esr_19_LC_3_5_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_19_LC_3_5_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_19_LC_3_5_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_19_LC_3_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34750),
            .lcout(\pid_alt.error_d_regZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94174),
            .ce(N__34723),
            .sr(N__92965));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_4_LC_3_6_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_4_LC_3_6_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_4_LC_3_6_4 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_4_LC_3_6_4  (
            .in0(N__54259),
            .in1(N__54115),
            .in2(_gnd_net_),
            .in3(N__39041),
            .lcout(\ppm_encoder_1.N_406 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_13_LC_3_6_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_13_LC_3_6_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_13_LC_3_6_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_13_LC_3_6_6  (
            .in0(_gnd_net_),
            .in1(N__50921),
            .in2(_gnd_net_),
            .in3(N__41881),
            .lcout(\ppm_encoder_1.N_440 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_esr_5_LC_3_7_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_5_LC_3_7_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_esr_5_LC_3_7_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.rudder_esr_5_LC_3_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42955),
            .lcout(\ppm_encoder_1.rudderZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94203),
            .ce(N__47984),
            .sr(N__86511));
    defparam \Commands_frame_decoder.source_alt_ki_0_LC_3_10_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_0_LC_3_10_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_0_LC_3_10_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_0_LC_3_10_0  (
            .in0(_gnd_net_),
            .in1(N__88306),
            .in2(_gnd_net_),
            .in3(N__93134),
            .lcout(alt_ki_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94254),
            .ce(N__42739),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_ki_1_LC_3_10_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_1_LC_3_10_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_1_LC_3_10_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_1_LC_3_10_1  (
            .in0(N__93135),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85527),
            .lcout(alt_ki_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94254),
            .ce(N__42739),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_ki_2_LC_3_10_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_2_LC_3_10_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_2_LC_3_10_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_2_LC_3_10_2  (
            .in0(_gnd_net_),
            .in1(N__92520),
            .in2(_gnd_net_),
            .in3(N__93136),
            .lcout(alt_ki_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94254),
            .ce(N__42739),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_ki_3_LC_3_10_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_3_LC_3_10_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_3_LC_3_10_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_3_LC_3_10_3  (
            .in0(N__93137),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__92330),
            .lcout(alt_ki_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94254),
            .ce(N__42739),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_ki_4_LC_3_10_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_4_LC_3_10_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_4_LC_3_10_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_4_LC_3_10_4  (
            .in0(_gnd_net_),
            .in1(N__88858),
            .in2(_gnd_net_),
            .in3(N__93138),
            .lcout(alt_ki_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94254),
            .ce(N__42739),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_ki_7_LC_3_10_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_7_LC_3_10_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_7_LC_3_10_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_7_LC_3_10_7  (
            .in0(N__93139),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__92131),
            .lcout(alt_ki_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94254),
            .ce(N__42739),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI11TA9_3_LC_3_13_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI11TA9_3_LC_3_13_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI11TA9_3_LC_3_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI11TA9_3_LC_3_13_0  (
            .in0(N__34822),
            .in1(N__36224),
            .in2(N__36964),
            .in3(N__35097),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI11TA9Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI3M511_3_LC_3_13_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI3M511_3_LC_3_13_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI3M511_3_LC_3_13_1 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI3M511_3_LC_3_13_1  (
            .in0(N__34846),
            .in1(N__35056),
            .in2(_gnd_net_),
            .in3(N__35088),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI3M511Z0Z_3 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNI3M511Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNICISB3_3_LC_3_13_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNICISB3_3_LC_3_13_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNICISB3_3_LC_3_13_2 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNICISB3_3_LC_3_13_2  (
            .in0(_gnd_net_),
            .in1(N__35098),
            .in2(N__34816),
            .in3(N__36225),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNICISB3Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI6P511_0_4_LC_3_13_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI6P511_0_4_LC_3_13_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI6P511_0_4_LC_3_13_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI6P511_0_4_LC_3_13_3  (
            .in0(N__35164),
            .in1(N__35148),
            .in2(_gnd_net_),
            .in3(N__35130),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI6P511_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_3_LC_3_13_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_3_LC_3_13_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_3_LC_3_13_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_3_LC_3_13_4  (
            .in0(N__35089),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94302),
            .ce(N__40512),
            .sr(N__86491));
    defparam \pid_alt.error_d_reg_prev_esr_RNILE0V5_2_LC_3_13_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNILE0V5_2_LC_3_13_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNILE0V5_2_LC_3_13_6 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNILE0V5_2_LC_3_13_6  (
            .in0(N__35020),
            .in1(_gnd_net_),
            .in2(N__35035),
            .in3(N__35044),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNILE0V5Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNILDG87_2_LC_3_13_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNILDG87_2_LC_3_13_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNILDG87_2_LC_3_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNILDG87_2_LC_3_13_7  (
            .in0(N__35043),
            .in1(N__35031),
            .in2(N__37020),
            .in3(N__35019),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNILDG87Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI171A6_5_LC_3_14_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI171A6_5_LC_3_14_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI171A6_5_LC_3_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI171A6_5_LC_3_14_0  (
            .in0(N__34929),
            .in1(N__35011),
            .in2(N__36904),
            .in3(N__37763),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI171A6Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI9S511_5_LC_3_14_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI9S511_5_LC_3_14_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI9S511_5_LC_3_14_1 .LUT_INIT=16'b1000100011101110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI9S511_5_LC_3_14_1  (
            .in0(N__35285),
            .in1(N__35307),
            .in2(_gnd_net_),
            .in3(N__35319),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI9S511Z0Z_5 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNI9S511Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIL81T2_5_LC_3_14_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIL81T2_5_LC_3_14_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIL81T2_5_LC_3_14_2 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIL81T2_5_LC_3_14_2  (
            .in0(N__34930),
            .in1(_gnd_net_),
            .in2(N__35005),
            .in3(N__37764),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIL81T2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNICV511_0_6_LC_3_14_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNICV511_0_6_LC_3_14_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNICV511_0_6_LC_3_14_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNICV511_0_6_LC_3_14_3  (
            .in0(N__35002),
            .in1(N__34972),
            .in2(_gnd_net_),
            .in3(N__34947),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNICV511_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_5_LC_3_14_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_5_LC_3_14_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_5_LC_3_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_5_LC_3_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35287),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94320),
            .ce(N__40510),
            .sr(N__86484));
    defparam \pid_alt.error_d_reg_prev_esr_RNICUVC3_4_LC_3_14_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNICUVC3_4_LC_3_14_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNICUVC3_4_LC_3_14_5 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNICUVC3_4_LC_3_14_5  (
            .in0(N__35260),
            .in1(N__35266),
            .in2(_gnd_net_),
            .in3(N__38634),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNICUVC3Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI9S511_0_5_LC_3_14_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI9S511_0_5_LC_3_14_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI9S511_0_5_LC_3_14_6 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI9S511_0_5_LC_3_14_6  (
            .in0(N__35320),
            .in1(_gnd_net_),
            .in2(N__35311),
            .in3(N__35286),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI9S511_0Z0Z_5 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNI9S511_0Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIOGSO6_4_LC_3_14_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOGSO6_4_LC_3_14_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOGSO6_4_LC_3_14_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIOGSO6_4_LC_3_14_7  (
            .in0(N__35259),
            .in1(N__36927),
            .in2(N__35245),
            .in3(N__38633),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIOGSO6Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI64JA4_12_LC_3_15_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI64JA4_12_LC_3_15_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI64JA4_12_LC_3_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI64JA4_12_LC_3_15_0  (
            .in0(N__35182),
            .in1(N__35172),
            .in2(N__37240),
            .in3(N__36113),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI64JA4Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIMJHM_0_13_LC_3_15_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIMJHM_0_13_LC_3_15_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIMJHM_0_13_LC_3_15_1 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIMJHM_0_13_LC_3_15_1  (
            .in0(N__35241),
            .in1(N__35217),
            .in2(_gnd_net_),
            .in3(N__35206),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIMJHM_0Z0Z_13 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIMJHM_0Z0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNISAO32_12_LC_3_15_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNISAO32_12_LC_3_15_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNISAO32_12_LC_3_15_2 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNISAO32_12_LC_3_15_2  (
            .in0(_gnd_net_),
            .in1(N__35173),
            .in2(N__35176),
            .in3(N__36114),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNISAO32Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIJGHM_12_LC_3_15_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIJGHM_12_LC_3_15_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIJGHM_12_LC_3_15_3 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIJGHM_12_LC_3_15_3  (
            .in0(N__35454),
            .in1(N__35463),
            .in2(_gnd_net_),
            .in3(N__35435),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_12_LC_3_15_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_12_LC_3_15_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_12_LC_3_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_12_LC_3_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35437),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94335),
            .ce(N__40507),
            .sr(N__86477));
    defparam \pid_alt.error_d_reg_prev_esr_RNIAPQ62_11_LC_3_15_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIAPQ62_11_LC_3_15_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIAPQ62_11_LC_3_15_5 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIAPQ62_11_LC_3_15_5  (
            .in0(N__35410),
            .in1(N__35416),
            .in2(_gnd_net_),
            .in3(N__35640),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIAPQ62Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIJGHM_0_12_LC_3_15_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIJGHM_0_12_LC_3_15_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIJGHM_0_12_LC_3_15_6 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIJGHM_0_12_LC_3_15_6  (
            .in0(N__35464),
            .in1(N__35455),
            .in2(_gnd_net_),
            .in3(N__35436),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIB8KD4_11_LC_3_15_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIB8KD4_11_LC_3_15_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIB8KD4_11_LC_3_15_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIB8KD4_11_LC_3_15_7  (
            .in0(N__35409),
            .in1(N__37275),
            .in2(N__35395),
            .in3(N__35639),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIB8KD4Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI88G14_14_LC_3_16_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI88G14_14_LC_3_16_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI88G14_14_LC_3_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI88G14_14_LC_3_16_0  (
            .in0(N__35392),
            .in1(N__35382),
            .in2(N__37183),
            .in3(N__36164),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI88G14Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNISPHM_0_15_LC_3_16_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNISPHM_0_15_LC_3_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNISPHM_0_15_LC_3_16_1 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNISPHM_0_15_LC_3_16_1  (
            .in0(N__40297),
            .in1(N__40534),
            .in2(_gnd_net_),
            .in3(N__40557),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNISPHM_0Z0Z_15 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNISPHM_0Z0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIOOO02_14_LC_3_16_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOOO02_14_LC_3_16_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOOO02_14_LC_3_16_2 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIOOO02_14_LC_3_16_2  (
            .in0(_gnd_net_),
            .in1(N__35383),
            .in2(N__35386),
            .in3(N__36165),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIOOO02Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIPMHM_14_LC_3_16_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIPMHM_14_LC_3_16_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIPMHM_14_LC_3_16_3 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIPMHM_14_LC_3_16_3  (
            .in0(N__35355),
            .in1(_gnd_net_),
            .in2(N__35332),
            .in3(N__35374),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIPMHMZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIPMHM_0_14_LC_3_16_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIPMHM_0_14_LC_3_16_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIPMHM_0_14_LC_3_16_4 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIPMHM_0_14_LC_3_16_4  (
            .in0(N__35373),
            .in1(N__35328),
            .in2(_gnd_net_),
            .in3(N__35354),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNICQF44_13_LC_3_16_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNICQF44_13_LC_3_16_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNICQF44_13_LC_3_16_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNICQF44_13_LC_3_16_5  (
            .in0(N__35619),
            .in1(N__37209),
            .in2(N__35359),
            .in3(N__37364),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNICQF44Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_14_LC_3_16_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_14_LC_3_16_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_14_LC_3_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_14_LC_3_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35356),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94350),
            .ce(N__40503),
            .sr(N__86467));
    defparam \pid_alt.error_d_reg_prev_esr_RNIGFN02_13_LC_3_16_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGFN02_13_LC_3_16_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGFN02_13_LC_3_16_7 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIGFN02_13_LC_3_16_7  (
            .in0(N__35620),
            .in1(N__35605),
            .in2(_gnd_net_),
            .in3(N__37365),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIGFN02Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIGKS02_17_LC_3_17_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGKS02_17_LC_3_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGKS02_17_LC_3_17_0 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIGKS02_17_LC_3_17_0  (
            .in0(N__35478),
            .in1(_gnd_net_),
            .in2(N__35512),
            .in3(N__35503),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIGKS02Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI53IM_18_LC_3_17_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI53IM_18_LC_3_17_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI53IM_18_LC_3_17_1 .LUT_INIT=16'b1111010101010000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI53IM_18_LC_3_17_1  (
            .in0(N__35527),
            .in1(_gnd_net_),
            .in2(N__35551),
            .in3(N__35581),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI8IQ14_18_LC_3_17_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI8IQ14_18_LC_3_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI8IQ14_18_LC_3_17_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI8IQ14_18_LC_3_17_2  (
            .in0(N__35596),
            .in1(N__37521),
            .in2(N__35599),
            .in3(N__37736),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI8IQ14Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI86IM_0_19_LC_3_17_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI86IM_0_19_LC_3_17_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI86IM_0_19_LC_3_17_4 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI86IM_0_19_LC_3_17_4  (
            .in0(N__35901),
            .in1(N__35829),
            .in2(_gnd_net_),
            .in3(N__35849),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI86IM_0Z0Z_19 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNI86IM_0Z0Z_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIOTT02_18_LC_3_17_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOTT02_18_LC_3_17_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOTT02_18_LC_3_17_5 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIOTT02_18_LC_3_17_5  (
            .in0(N__37737),
            .in1(_gnd_net_),
            .in2(N__35590),
            .in3(N__35587),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIOTT02Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI53IM_0_18_LC_3_17_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI53IM_0_18_LC_3_17_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI53IM_0_18_LC_3_17_6 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI53IM_0_18_LC_3_17_6  (
            .in0(N__35580),
            .in1(N__35547),
            .in2(_gnd_net_),
            .in3(N__35526),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIOVN14_17_LC_3_17_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOVN14_17_LC_3_17_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOVN14_17_LC_3_17_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIOVN14_17_LC_3_17_7  (
            .in0(N__35502),
            .in1(N__37566),
            .in2(N__35485),
            .in3(N__35477),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIOVN14Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_20_LC_3_18_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_20_LC_3_18_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_20_LC_3_18_1 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_20_LC_3_18_1  (
            .in0(_gnd_net_),
            .in1(N__35765),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94371),
            .ce(N__40499),
            .sr(N__86458));
    defparam \pid_alt.error_d_reg_prev_esr_RNI86IM_19_LC_3_18_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI86IM_19_LC_3_18_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI86IM_19_LC_3_18_2 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI86IM_19_LC_3_18_2  (
            .in0(N__35902),
            .in1(N__35830),
            .in2(_gnd_net_),
            .in3(N__35850),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI86IMZ0Z_19 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNI86IMZ0Z_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIK3024_19_LC_3_18_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIK3024_19_LC_3_18_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIK3024_19_LC_3_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIK3024_19_LC_3_18_3  (
            .in0(N__37491),
            .in1(N__35859),
            .in2(N__35872),
            .in3(N__36137),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIK3024Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIS5212_19_LC_3_18_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIS5212_19_LC_3_18_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIS5212_19_LC_3_18_4 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIS5212_19_LC_3_18_4  (
            .in0(N__36138),
            .in1(_gnd_net_),
            .in2(N__35863),
            .in3(N__35869),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIS5212Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIGGKM_20_LC_3_18_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGGKM_20_LC_3_18_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGGKM_20_LC_3_18_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIGGKM_20_LC_3_18_5  (
            .in0(N__35729),
            .in1(N__35763),
            .in2(_gnd_net_),
            .in3(N__35800),
            .lcout(\pid_alt.un1_pid_prereg_236_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_19_LC_3_18_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_19_LC_3_18_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_19_LC_3_18_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_19_LC_3_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35851),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94371),
            .ce(N__40499),
            .sr(N__86458));
    defparam \pid_alt.error_d_reg_prev_esr_RNICG9B1_1_20_LC_3_18_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNICG9B1_1_20_LC_3_18_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNICG9B1_1_20_LC_3_18_7 .LUT_INIT=16'b0100001010111101;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNICG9B1_1_20_LC_3_18_7  (
            .in0(N__35804),
            .in1(N__35764),
            .in2(N__35737),
            .in3(N__35685),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNICG9B1_1Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI4CCV_10_LC_3_19_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI4CCV_10_LC_3_19_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI4CCV_10_LC_3_19_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNI4CCV_10_LC_3_19_0  (
            .in0(N__38105),
            .in1(N__38130),
            .in2(N__38083),
            .in3(N__36096),
            .lcout(\pid_alt.m35_e_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_10_LC_3_19_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_10_LC_3_19_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_10_LC_3_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_10_LC_3_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35659),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94379),
            .ce(N__40498),
            .sr(N__86453));
    defparam \pid_alt.error_i_acumm_prereg_esr_12_LC_3_19_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_12_LC_3_19_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_12_LC_3_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_12_LC_3_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35641),
            .lcout(\pid_alt.error_i_acumm7lto12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94379),
            .ce(N__40498),
            .sr(N__86453));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNICP62_10_LC_3_19_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNICP62_10_LC_3_19_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNICP62_10_LC_3_19_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNICP62_10_LC_3_19_4  (
            .in0(_gnd_net_),
            .in1(N__36095),
            .in2(_gnd_net_),
            .in3(N__35993),
            .lcout(),
            .ltout(\pid_alt.m21_e_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIIO7C2_2_LC_3_19_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIIO7C2_2_LC_3_19_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIIO7C2_2_LC_3_19_5 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNIIO7C2_2_LC_3_19_5  (
            .in0(N__38047),
            .in1(N__36060),
            .in2(N__36082),
            .in3(N__36075),
            .lcout(\pid_alt.m21_e_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_2_LC_3_19_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_2_LC_3_19_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_2_LC_3_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_2_LC_3_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37070),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94379),
            .ce(N__40498),
            .sr(N__86453));
    defparam \pid_alt.error_i_acumm_prereg_esr_3_LC_3_19_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_3_LC_3_19_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_3_LC_3_19_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_3_LC_3_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37013),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94379),
            .ce(N__40498),
            .sr(N__86453));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI4SOH2_10_LC_3_20_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI4SOH2_10_LC_3_20_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI4SOH2_10_LC_3_20_0 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNI4SOH2_10_LC_3_20_0  (
            .in0(N__38657),
            .in1(N__35960),
            .in2(N__36049),
            .in3(N__35922),
            .lcout(\pid_alt.N_62_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIRRP7_14_LC_3_20_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIRRP7_14_LC_3_20_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIRRP7_14_LC_3_20_2 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNIRRP7_14_LC_3_20_2  (
            .in0(N__36238),
            .in1(N__36151),
            .in2(N__36184),
            .in3(N__37351),
            .lcout(\pid_alt.N_545 ),
            .ltout(\pid_alt.N_545_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI175B_12_LC_3_20_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI175B_12_LC_3_20_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI175B_12_LC_3_20_3 .LUT_INIT=16'b1011101011111010;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNI175B_12_LC_3_20_3  (
            .in0(N__57611),
            .in1(N__57558),
            .in2(N__35998),
            .in3(N__35994),
            .lcout(\pid_alt.N_158 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIFJA3_14_LC_3_20_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIFJA3_14_LC_3_20_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIFJA3_14_LC_3_20_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNIFJA3_14_LC_3_20_4  (
            .in0(N__36180),
            .in1(N__36150),
            .in2(_gnd_net_),
            .in3(N__37350),
            .lcout(),
            .ltout(\pid_alt.error_i_acumm_prereg_esr_RNIFJA3Z0Z_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIAP1A_13_LC_3_20_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIAP1A_13_LC_3_20_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIAP1A_13_LC_3_20_5 .LUT_INIT=16'b1011101010101010;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNIAP1A_13_LC_3_20_5  (
            .in0(N__57610),
            .in1(N__57557),
            .in2(N__35929),
            .in3(N__36237),
            .lcout(\pid_alt.N_9_0 ),
            .ltout(\pid_alt.N_9_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIO7B05_21_LC_3_20_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIO7B05_21_LC_3_20_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIO7B05_21_LC_3_20_6 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNIO7B05_21_LC_3_20_6  (
            .in0(N__57612),
            .in1(N__38782),
            .in2(N__36274),
            .in3(N__36271),
            .lcout(\pid_alt.N_111 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIC8F4_16_LC_3_20_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIC8F4_16_LC_3_20_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIC8F4_16_LC_3_20_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNIC8F4_16_LC_3_20_7  (
            .in0(N__37723),
            .in1(N__36265),
            .in2(N__36253),
            .in3(N__36124),
            .lcout(\pid_alt.m7_e_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_4_LC_3_21_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_4_LC_3_21_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_4_LC_3_21_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_4_LC_3_21_0  (
            .in0(N__36229),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_i_acumm7lto4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94395),
            .ce(N__40496),
            .sr(N__86445));
    defparam \pid_alt.error_i_acumm_prereg_esr_17_LC_3_21_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_17_LC_3_21_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_17_LC_3_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_17_LC_3_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36205),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94395),
            .ce(N__40496),
            .sr(N__86445));
    defparam \pid_alt.error_i_acumm_prereg_esr_15_LC_3_21_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_15_LC_3_21_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_15_LC_3_21_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_15_LC_3_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36172),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94395),
            .ce(N__40496),
            .sr(N__86445));
    defparam \pid_alt.error_i_acumm_prereg_esr_8_LC_3_21_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_8_LC_3_21_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_8_LC_3_21_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_8_LC_3_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39433),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94395),
            .ce(N__40496),
            .sr(N__86445));
    defparam \pid_alt.error_i_acumm_prereg_esr_20_LC_3_21_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_20_LC_3_21_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_20_LC_3_21_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_20_LC_3_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36142),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94395),
            .ce(N__40496),
            .sr(N__86445));
    defparam \pid_alt.error_i_acumm_prereg_esr_13_LC_3_21_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_13_LC_3_21_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_13_LC_3_21_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_13_LC_3_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36118),
            .lcout(\pid_alt.error_i_acumm7lto13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94395),
            .ce(N__40496),
            .sr(N__86445));
    defparam \Commands_frame_decoder.source_alt_kp_0_e_0_4_LC_3_22_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_0_e_0_4_LC_3_22_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kp_0_e_0_4_LC_3_22_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_0_e_0_4_LC_3_22_4  (
            .in0(_gnd_net_),
            .in1(N__88685),
            .in2(_gnd_net_),
            .in3(N__93151),
            .lcout(alt_kp_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94398),
            .ce(N__48692),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kp_e_0_6_LC_3_22_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_6_LC_3_22_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_6_LC_3_22_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_e_0_6_LC_3_22_5  (
            .in0(N__93152),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__92123),
            .lcout(alt_kp_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94398),
            .ce(N__48692),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kp_e_0_0_LC_3_23_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_0_LC_3_23_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_0_LC_3_23_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_e_0_0_LC_3_23_1  (
            .in0(_gnd_net_),
            .in1(N__88307),
            .in2(_gnd_net_),
            .in3(N__93153),
            .lcout(alt_kp_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94404),
            .ce(N__48708),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIBHIH2_2_LC_4_2_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIBHIH2_2_LC_4_2_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIBHIH2_2_LC_4_2_0 .LUT_INIT=16'b1110000100011110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIBHIH2_2_LC_4_2_0  (
            .in0(N__44328),
            .in1(N__47480),
            .in2(N__46645),
            .in3(N__41786),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI3K6R5_5_LC_4_2_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI3K6R5_5_LC_4_2_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI3K6R5_5_LC_4_2_1 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI3K6R5_5_LC_4_2_1  (
            .in0(N__43944),
            .in1(N__36352),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\ppm_encoder_1.init_pulses_RNI3K6R5Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIT9FE2_13_LC_4_2_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIT9FE2_13_LC_4_2_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIT9FE2_13_LC_4_2_2 .LUT_INIT=16'b1110000100011110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIT9FE2_13_LC_4_2_2  (
            .in0(N__44329),
            .in1(N__47481),
            .in2(N__41880),
            .in3(N__41787),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_2_LC_4_2_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_2_LC_4_2_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_2_LC_4_2_4 .LUT_INIT=16'b0011000001110101;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_2_LC_4_2_4  (
            .in0(N__47434),
            .in1(N__36454),
            .in2(N__50594),
            .in3(N__40813),
            .lcout(),
            .ltout(\ppm_encoder_1.pulses2count_9_i_3_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_2_LC_4_2_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_2_LC_4_2_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_2_LC_4_2_5 .LUT_INIT=16'b1111101011111110;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_2_LC_4_2_5  (
            .in0(N__47483),
            .in1(N__50960),
            .in2(N__36283),
            .in3(N__46642),
            .lcout(\ppm_encoder_1.pulses2count_9_i_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_1_LC_4_2_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_1_LC_4_2_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_1_LC_4_2_6 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_1_LC_4_2_6  (
            .in0(N__50959),
            .in1(N__36280),
            .in2(_gnd_net_),
            .in3(N__40415),
            .lcout(\ppm_encoder_1.pulses2count_9_0_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_1_LC_4_2_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_1_LC_4_2_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_1_LC_4_2_7 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_1_LC_4_2_7  (
            .in0(N__47482),
            .in1(N__40696),
            .in2(_gnd_net_),
            .in3(N__47433),
            .lcout(\ppm_encoder_1.pulses2count_9_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIPH6J4_5_LC_4_3_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIPH6J4_5_LC_4_3_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIPH6J4_5_LC_4_3_0 .LUT_INIT=16'b1010010110010110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIPH6J4_5_LC_4_3_0  (
            .in0(N__41772),
            .in1(N__44456),
            .in2(N__49968),
            .in3(N__36334),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIDN3K_2_LC_4_3_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIDN3K_2_LC_4_3_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIDN3K_2_LC_4_3_1 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIDN3K_2_LC_4_3_1  (
            .in0(N__44906),
            .in1(_gnd_net_),
            .in2(N__42080),
            .in3(N__38952),
            .lcout(\ppm_encoder_1.N_513 ),
            .ltout(\ppm_encoder_1.N_513_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIFLIH2_6_LC_4_3_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIFLIH2_6_LC_4_3_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIFLIH2_6_LC_4_3_2 .LUT_INIT=16'b1001100110010110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIFLIH2_6_LC_4_3_2  (
            .in0(N__41771),
            .in1(N__49126),
            .in2(N__36346),
            .in3(N__44330),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIHGIP3_2_LC_4_3_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIHGIP3_2_LC_4_3_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIHGIP3_2_LC_4_3_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIHGIP3_2_LC_4_3_3  (
            .in0(_gnd_net_),
            .in1(N__36343),
            .in2(_gnd_net_),
            .in3(N__43569),
            .lcout(\ppm_encoder_1.init_pulses_RNIHGIP3Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_LC_4_3_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_LC_4_3_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_LC_4_3_5 .LUT_INIT=16'b0000101000000110;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_LC_4_3_5  (
            .in0(N__42071),
            .in1(N__54260),
            .in2(N__71068),
            .in3(N__52741),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94137),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNI1R011_5_LC_4_3_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNI1R011_5_LC_4_3_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNI1R011_5_LC_4_3_6 .LUT_INIT=16'b0000001101000100;
    LogicCell40 \ppm_encoder_1.throttle_RNI1R011_5_LC_4_3_6  (
            .in0(N__36430),
            .in1(N__42067),
            .in2(N__36544),
            .in3(N__44905),
            .lcout(\ppm_encoder_1.un2_throttle_0_0_2_5 ),
            .ltout(\ppm_encoder_1.un2_throttle_0_0_2_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIBLNA2_5_LC_4_3_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIBLNA2_5_LC_4_3_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIBLNA2_5_LC_4_3_7 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \ppm_encoder_1.throttle_RNIBLNA2_5_LC_4_3_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__36337),
            .in3(N__49911),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_9_LC_4_4_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_9_LC_4_4_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_9_LC_4_4_0 .LUT_INIT=16'b0000010100000001;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_9_LC_4_4_0  (
            .in0(N__46927),
            .in1(N__50949),
            .in2(N__44734),
            .in3(N__46531),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94149),
            .ce(N__50384),
            .sr(N__86516));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_1_LC_4_4_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_1_LC_4_4_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_1_LC_4_4_2 .LUT_INIT=16'b1111111110100000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_1_LC_4_4_2  (
            .in0(N__36414),
            .in1(_gnd_net_),
            .in2(N__50599),
            .in3(N__36328),
            .lcout(\ppm_encoder_1.pulses2count_9_0_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIJLS91_1_LC_4_4_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIJLS91_1_LC_4_4_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIJLS91_1_LC_4_4_4 .LUT_INIT=16'b0001111100010001;
    LogicCell40 \ppm_encoder_1.throttle_RNIJLS91_1_LC_4_4_4  (
            .in0(N__47343),
            .in1(N__40692),
            .in2(N__36415),
            .in3(N__44649),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIHI8E1_3_LC_4_4_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIHI8E1_3_LC_4_4_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIHI8E1_3_LC_4_4_5 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \ppm_encoder_1.throttle_RNIHI8E1_3_LC_4_4_5  (
            .in0(N__44650),
            .in1(N__50419),
            .in2(N__50529),
            .in3(N__44570),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIFBLQ_1_LC_4_4_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIFBLQ_1_LC_4_4_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIFBLQ_1_LC_4_4_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_RNIFBLQ_1_LC_4_4_6  (
            .in0(N__44571),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54114),
            .lcout(\ppm_encoder_1.N_529 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_esr_RNIAQM91_5_LC_4_4_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_RNIAQM91_5_LC_4_4_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.rudder_esr_RNIAQM91_5_LC_4_4_7 .LUT_INIT=16'b0000110001011101;
    LogicCell40 \ppm_encoder_1.rudder_esr_RNIAQM91_5_LC_4_4_7  (
            .in0(N__51067),
            .in1(N__38951),
            .in2(N__36373),
            .in3(N__47342),
            .lcout(\ppm_encoder_1.N_307 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI4TGA_2_LC_4_5_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI4TGA_2_LC_4_5_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI4TGA_2_LC_4_5_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI4TGA_2_LC_4_5_0  (
            .in0(_gnd_net_),
            .in1(N__42078),
            .in2(_gnd_net_),
            .in3(N__38948),
            .lcout(\ppm_encoder_1.N_507 ),
            .ltout(\ppm_encoder_1.N_507_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIFG8E1_2_LC_4_5_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIFG8E1_2_LC_4_5_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIFG8E1_2_LC_4_5_1 .LUT_INIT=16'b0111001101010000;
    LogicCell40 \ppm_encoder_1.throttle_RNIFG8E1_2_LC_4_5_1  (
            .in0(N__36450),
            .in1(N__50637),
            .in2(N__36361),
            .in3(N__44572),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNICJSS4_2_LC_4_5_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNICJSS4_2_LC_4_5_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNICJSS4_2_LC_4_5_2 .LUT_INIT=16'b1001100110010110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNICJSS4_2_LC_4_5_2  (
            .in0(N__46644),
            .in1(N__41758),
            .in2(N__36358),
            .in3(N__39004),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_0_axb_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIIIS46_2_LC_4_5_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIIIS46_2_LC_4_5_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIIIS46_2_LC_4_5_3 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIIIS46_2_LC_4_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__36355),
            .in3(N__43562),
            .lcout(\ppm_encoder_1.init_pulses_RNIIIS46Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_0_LC_4_5_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_0_LC_4_5_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.PPM_STATE_0_LC_4_5_4 .LUT_INIT=16'b1100110011011101;
    LogicCell40 \ppm_encoder_1.PPM_STATE_0_LC_4_5_4  (
            .in0(N__49780),
            .in1(N__49740),
            .in2(_gnd_net_),
            .in3(N__49855),
            .lcout(\ppm_encoder_1.PPM_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94160),
            .ce(),
            .sr(N__86515));
    defparam \ppm_encoder_1.init_pulses_RNI6VV71_2_LC_4_5_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI6VV71_2_LC_4_5_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI6VV71_2_LC_4_5_5 .LUT_INIT=16'b1100110001101100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI6VV71_2_LC_4_5_5  (
            .in0(N__42156),
            .in1(N__46643),
            .in2(N__43717),
            .in3(N__52742),
            .lcout(\ppm_encoder_1.N_259_i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_RNIMINS_0_LC_4_5_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNIMINS_0_LC_4_5_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNIMINS_0_LC_4_5_6 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNIMINS_0_LC_4_5_6  (
            .in0(N__49779),
            .in1(N__43701),
            .in2(N__49531),
            .in3(N__42155),
            .lcout(\ppm_encoder_1.PPM_STATE_RNIMINSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI3O6G_2_LC_4_5_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI3O6G_2_LC_4_5_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI3O6G_2_LC_4_5_7 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI3O6G_2_LC_4_5_7  (
            .in0(N__38947),
            .in1(N__44891),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\ppm_encoder_1.N_509 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_LC_4_6_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_LC_4_6_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_LC_4_6_0 .LUT_INIT=16'b1111111011011100;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_LC_4_6_0  (
            .in0(N__52769),
            .in1(N__71029),
            .in2(N__47197),
            .in3(N__44898),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94175),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_rep1_LC_4_6_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_rep1_LC_4_6_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_rep1_LC_4_6_1 .LUT_INIT=16'b0101000000010001;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_3_rep1_LC_4_6_1  (
            .in0(N__71028),
            .in1(N__46894),
            .in2(N__43726),
            .in3(N__52770),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94175),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIE5081_8_LC_4_6_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIE5081_8_LC_4_6_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIE5081_8_LC_4_6_2 .LUT_INIT=16'b1001110011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIE5081_8_LC_4_6_2  (
            .in0(N__52768),
            .in1(N__48963),
            .in2(N__53697),
            .in3(N__53808),
            .lcout(\ppm_encoder_1.N_264_i_i ),
            .ltout(\ppm_encoder_1.N_264_i_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIL76H6_8_LC_4_6_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIL76H6_8_LC_4_6_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIL76H6_8_LC_4_6_3 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIL76H6_8_LC_4_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__36388),
            .in3(N__36379),
            .lcout(\ppm_encoder_1.init_pulses_RNIL76H6Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIFC6O_8_LC_4_6_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIFC6O_8_LC_4_6_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIFC6O_8_LC_4_6_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \ppm_encoder_1.elevator_RNIFC6O_8_LC_4_6_4  (
            .in0(N__44774),
            .in1(N__42079),
            .in2(_gnd_net_),
            .in3(N__44897),
            .lcout(),
            .ltout(\ppm_encoder_1.N_465_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_RNIDD8O2_8_LC_4_6_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_RNIDD8O2_8_LC_4_6_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.rudder_RNIDD8O2_8_LC_4_6_5 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \ppm_encoder_1.rudder_RNIDD8O2_8_LC_4_6_5  (
            .in0(N__44466),
            .in1(N__46995),
            .in2(N__36385),
            .in3(N__53682),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_2_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI72695_8_LC_4_6_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI72695_8_LC_4_6_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI72695_8_LC_4_6_6 .LUT_INIT=16'b0110011001101001;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI72695_8_LC_4_6_6  (
            .in0(N__48962),
            .in1(N__41759),
            .in2(N__36382),
            .in3(N__39049),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_6_LC_4_7_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_6_LC_4_7_0 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.throttle_6_LC_4_7_0 .LUT_INIT=16'b1100001110101010;
    LogicCell40 \ppm_encoder_1.throttle_6_LC_4_7_0  (
            .in0(N__44937),
            .in1(N__36675),
            .in2(N__36472),
            .in3(N__51224),
            .lcout(\ppm_encoder_1.throttleZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94189),
            .ce(),
            .sr(N__86510));
    defparam \ppm_encoder_1.throttle_4_LC_4_7_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_4_LC_4_7_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_4_LC_4_7_1 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.throttle_4_LC_4_7_1  (
            .in0(N__36493),
            .in1(N__39844),
            .in2(N__51323),
            .in3(N__39042),
            .lcout(\ppm_encoder_1.throttleZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94189),
            .ce(),
            .sr(N__86510));
    defparam \ppm_encoder_1.aileron_8_LC_4_7_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_8_LC_4_7_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_8_LC_4_7_2 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.aileron_8_LC_4_7_2  (
            .in0(N__54385),
            .in1(N__47788),
            .in2(N__44814),
            .in3(N__51234),
            .lcout(\ppm_encoder_1.aileronZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94189),
            .ce(),
            .sr(N__86510));
    defparam \ppm_encoder_1.throttle_3_LC_4_7_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_3_LC_4_7_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_3_LC_4_7_3 .LUT_INIT=16'b1101100001110010;
    LogicCell40 \ppm_encoder_1.throttle_3_LC_4_7_3  (
            .in0(N__51222),
            .in1(N__36817),
            .in2(N__50528),
            .in3(N__36505),
            .lcout(\ppm_encoder_1.throttleZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94189),
            .ce(),
            .sr(N__86510));
    defparam \ppm_encoder_1.elevator_8_LC_4_7_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_8_LC_4_7_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_8_LC_4_7_5 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.elevator_8_LC_4_7_5  (
            .in0(N__54544),
            .in1(N__47653),
            .in2(N__51322),
            .in3(N__44778),
            .lcout(\ppm_encoder_1.elevatorZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94189),
            .ce(),
            .sr(N__86510));
    defparam \ppm_encoder_1.throttle_2_LC_4_7_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_2_LC_4_7_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.throttle_2_LC_4_7_6 .LUT_INIT=16'b0010111011100010;
    LogicCell40 \ppm_encoder_1.throttle_2_LC_4_7_6  (
            .in0(N__36449),
            .in1(N__51223),
            .in2(N__36853),
            .in3(N__36517),
            .lcout(\ppm_encoder_1.throttleZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94189),
            .ce(),
            .sr(N__86510));
    defparam \ppm_encoder_1.aileron_5_LC_4_7_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_5_LC_4_7_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_5_LC_4_7_7 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.aileron_5_LC_4_7_7  (
            .in0(N__47830),
            .in1(N__59290),
            .in2(N__51321),
            .in3(N__36429),
            .lcout(\ppm_encoder_1.aileronZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94189),
            .ce(),
            .sr(N__86510));
    defparam \ppm_encoder_1.throttle_1_LC_4_8_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_1_LC_4_8_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_1_LC_4_8_0 .LUT_INIT=16'b1001100111110000;
    LogicCell40 \ppm_encoder_1.throttle_1_LC_4_8_0  (
            .in0(N__36526),
            .in1(N__36871),
            .in2(N__36410),
            .in3(N__51297),
            .lcout(\ppm_encoder_1.throttleZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94204),
            .ce(),
            .sr(N__86508));
    defparam \ppm_encoder_1.throttle_10_LC_4_8_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_10_LC_4_8_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_10_LC_4_8_1 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.throttle_10_LC_4_8_1  (
            .in0(N__36567),
            .in1(N__36610),
            .in2(N__51355),
            .in3(N__46472),
            .lcout(\ppm_encoder_1.throttleZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94204),
            .ce(),
            .sr(N__86508));
    defparam \ppm_encoder_1.throttle_11_LC_4_8_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_11_LC_4_8_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_11_LC_4_8_2 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.throttle_11_LC_4_8_2  (
            .in0(N__36697),
            .in1(N__36598),
            .in2(N__40650),
            .in3(N__51295),
            .lcout(\ppm_encoder_1.throttleZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94204),
            .ce(),
            .sr(N__86508));
    defparam \ppm_encoder_1.throttle_5_LC_4_8_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_5_LC_4_8_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_5_LC_4_8_5 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.throttle_5_LC_4_8_5  (
            .in0(N__36481),
            .in1(N__39808),
            .in2(N__51356),
            .in3(N__36540),
            .lcout(\ppm_encoder_1.throttleZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94204),
            .ce(),
            .sr(N__86508));
    defparam \ppm_encoder_1.throttle_13_LC_4_8_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_13_LC_4_8_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.throttle_13_LC_4_8_6 .LUT_INIT=16'b1001100111110000;
    LogicCell40 \ppm_encoder_1.throttle_13_LC_4_8_6  (
            .in0(N__39628),
            .in1(N__36583),
            .in2(N__39076),
            .in3(N__51296),
            .lcout(\ppm_encoder_1.throttleZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94204),
            .ce(),
            .sr(N__86508));
    defparam \ppm_encoder_1.un1_throttle_cry_0_c_LC_4_9_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_0_c_LC_4_9_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_0_c_LC_4_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_0_c_LC_4_9_0  (
            .in0(_gnd_net_),
            .in1(N__41949),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_9_0_),
            .carryout(\ppm_encoder_1.un1_throttle_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_0_THRU_LUT4_0_LC_4_9_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_0_THRU_LUT4_0_LC_4_9_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_0_THRU_LUT4_0_LC_4_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_0_THRU_LUT4_0_LC_4_9_1  (
            .in0(_gnd_net_),
            .in1(N__36870),
            .in2(N__65866),
            .in3(N__36520),
            .lcout(\ppm_encoder_1.un1_throttle_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_0 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_1_THRU_LUT4_0_LC_4_9_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_1_THRU_LUT4_0_LC_4_9_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_1_THRU_LUT4_0_LC_4_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_1_THRU_LUT4_0_LC_4_9_2  (
            .in0(_gnd_net_),
            .in1(N__36846),
            .in2(_gnd_net_),
            .in3(N__36508),
            .lcout(\ppm_encoder_1.un1_throttle_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_1 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_2_THRU_LUT4_0_LC_4_9_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_2_THRU_LUT4_0_LC_4_9_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_2_THRU_LUT4_0_LC_4_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_2_THRU_LUT4_0_LC_4_9_3  (
            .in0(_gnd_net_),
            .in1(N__36816),
            .in2(N__65867),
            .in3(N__36496),
            .lcout(\ppm_encoder_1.un1_throttle_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_2 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_3_THRU_LUT4_0_LC_4_9_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_3_THRU_LUT4_0_LC_4_9_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_3_THRU_LUT4_0_LC_4_9_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_3_THRU_LUT4_0_LC_4_9_4  (
            .in0(_gnd_net_),
            .in1(N__39843),
            .in2(_gnd_net_),
            .in3(N__36484),
            .lcout(\ppm_encoder_1.un1_throttle_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_3 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_4_THRU_LUT4_0_LC_4_9_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_4_THRU_LUT4_0_LC_4_9_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_4_THRU_LUT4_0_LC_4_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_4_THRU_LUT4_0_LC_4_9_5  (
            .in0(_gnd_net_),
            .in1(N__39804),
            .in2(_gnd_net_),
            .in3(N__36475),
            .lcout(\ppm_encoder_1.un1_throttle_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_4 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_5_THRU_LUT4_0_LC_4_9_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_5_THRU_LUT4_0_LC_4_9_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_5_THRU_LUT4_0_LC_4_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_5_THRU_LUT4_0_LC_4_9_6  (
            .in0(_gnd_net_),
            .in1(N__65822),
            .in2(N__36676),
            .in3(N__36457),
            .lcout(\ppm_encoder_1.un1_throttle_cry_5_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_5 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_6_THRU_LUT4_0_LC_4_9_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_6_THRU_LUT4_0_LC_4_9_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_6_THRU_LUT4_0_LC_4_9_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_6_THRU_LUT4_0_LC_4_9_7  (
            .in0(_gnd_net_),
            .in1(N__45128),
            .in2(_gnd_net_),
            .in3(N__36619),
            .lcout(\ppm_encoder_1.un1_throttle_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_6 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_7_THRU_LUT4_0_LC_4_10_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_7_THRU_LUT4_0_LC_4_10_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_7_THRU_LUT4_0_LC_4_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_7_THRU_LUT4_0_LC_4_10_0  (
            .in0(_gnd_net_),
            .in1(N__45092),
            .in2(_gnd_net_),
            .in3(N__36616),
            .lcout(\ppm_encoder_1.un1_throttle_cry_7_THRU_CO ),
            .ltout(),
            .carryin(bfn_4_10_0_),
            .carryout(\ppm_encoder_1.un1_throttle_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_8_THRU_LUT4_0_LC_4_10_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_8_THRU_LUT4_0_LC_4_10_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_8_THRU_LUT4_0_LC_4_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_8_THRU_LUT4_0_LC_4_10_1  (
            .in0(_gnd_net_),
            .in1(N__45017),
            .in2(_gnd_net_),
            .in3(N__36613),
            .lcout(\ppm_encoder_1.un1_throttle_cry_8_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_8 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_9_THRU_LUT4_0_LC_4_10_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_9_THRU_LUT4_0_LC_4_10_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_9_THRU_LUT4_0_LC_4_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_9_THRU_LUT4_0_LC_4_10_2  (
            .in0(_gnd_net_),
            .in1(N__36560),
            .in2(_gnd_net_),
            .in3(N__36601),
            .lcout(\ppm_encoder_1.un1_throttle_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_9 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_10_THRU_LUT4_0_LC_4_10_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_10_THRU_LUT4_0_LC_4_10_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_10_THRU_LUT4_0_LC_4_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_10_THRU_LUT4_0_LC_4_10_3  (
            .in0(_gnd_net_),
            .in1(N__36692),
            .in2(_gnd_net_),
            .in3(N__36589),
            .lcout(\ppm_encoder_1.un1_throttle_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_10 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_11_THRU_LUT4_0_LC_4_10_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_11_THRU_LUT4_0_LC_4_10_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_11_THRU_LUT4_0_LC_4_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_11_THRU_LUT4_0_LC_4_10_4  (
            .in0(_gnd_net_),
            .in1(N__42027),
            .in2(_gnd_net_),
            .in3(N__36586),
            .lcout(\ppm_encoder_1.un1_throttle_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_11 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_12_THRU_LUT4_0_LC_4_10_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_12_THRU_LUT4_0_LC_4_10_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_12_THRU_LUT4_0_LC_4_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_12_THRU_LUT4_0_LC_4_10_5  (
            .in0(_gnd_net_),
            .in1(N__39627),
            .in2(N__65854),
            .in3(N__36574),
            .lcout(\ppm_encoder_1.un1_throttle_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_12 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_esr_14_LC_4_10_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_esr_14_LC_4_10_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_esr_14_LC_4_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.throttle_esr_14_LC_4_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36571),
            .lcout(\ppm_encoder_1.throttleZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94236),
            .ce(N__47986),
            .sr(N__86502));
    defparam \pid_alt.source_pid_1_10_LC_4_11_0 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_10_LC_4_11_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_10_LC_4_11_0 .LUT_INIT=16'b1111101001110010;
    LogicCell40 \pid_alt.source_pid_1_10_LC_4_11_0  (
            .in0(N__69003),
            .in1(N__36638),
            .in2(N__36568),
            .in3(N__39265),
            .lcout(throttle_order_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94255),
            .ce(),
            .sr(N__39568));
    defparam \pid_alt.pid_prereg_esr_RNIIM6H1_0_6_LC_4_11_1 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIIM6H1_0_6_LC_4_11_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIIM6H1_0_6_LC_4_11_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIIM6H1_0_6_LC_4_11_1  (
            .in0(N__39372),
            .in1(N__39351),
            .in2(N__39331),
            .in3(N__39303),
            .lcout(),
            .ltout(\pid_alt.source_pid_1_sqmuxa_0_a2_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNI4GSA2_10_LC_4_11_2 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNI4GSA2_10_LC_4_11_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNI4GSA2_10_LC_4_11_2 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \pid_alt.pid_prereg_esr_RNI4GSA2_10_LC_4_11_2  (
            .in0(N__69002),
            .in1(N__39285),
            .in2(N__36700),
            .in3(N__39264),
            .lcout(\pid_alt.source_pid_1_sqmuxa_0_a2_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.source_pid_1_11_LC_4_11_3 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_11_LC_4_11_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_11_LC_4_11_3 .LUT_INIT=16'b1010111111001100;
    LogicCell40 \pid_alt.source_pid_1_11_LC_4_11_3  (
            .in0(N__39286),
            .in1(N__36696),
            .in2(N__36648),
            .in3(N__69004),
            .lcout(throttle_order_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94255),
            .ce(),
            .sr(N__39568));
    defparam \pid_alt.source_pid_1_6_LC_4_11_4 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_6_LC_4_11_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_6_LC_4_11_4 .LUT_INIT=16'b1010110011111100;
    LogicCell40 \pid_alt.source_pid_1_6_LC_4_11_4  (
            .in0(N__39304),
            .in1(N__36671),
            .in2(N__69024),
            .in3(N__36642),
            .lcout(throttle_order_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94255),
            .ce(),
            .sr(N__39568));
    defparam \pid_alt.source_pid_1_7_LC_4_11_5 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_7_LC_4_11_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_7_LC_4_11_5 .LUT_INIT=16'b1111110001110100;
    LogicCell40 \pid_alt.source_pid_1_7_LC_4_11_5  (
            .in0(N__36643),
            .in1(N__69008),
            .in2(N__45132),
            .in3(N__39352),
            .lcout(throttle_order_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94255),
            .ce(),
            .sr(N__39568));
    defparam \pid_alt.source_pid_1_8_LC_4_11_6 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_8_LC_4_11_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_8_LC_4_11_6 .LUT_INIT=16'b1111101001110010;
    LogicCell40 \pid_alt.source_pid_1_8_LC_4_11_6  (
            .in0(N__69009),
            .in1(N__36644),
            .in2(N__45102),
            .in3(N__39373),
            .lcout(throttle_order_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94255),
            .ce(),
            .sr(N__39568));
    defparam \pid_alt.source_pid_1_9_LC_4_11_7 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_9_LC_4_11_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_9_LC_4_11_7 .LUT_INIT=16'b1010111111001100;
    LogicCell40 \pid_alt.source_pid_1_9_LC_4_11_7  (
            .in0(N__39329),
            .in1(N__45021),
            .in2(N__36649),
            .in3(N__69010),
            .lcout(throttle_order_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94255),
            .ce(),
            .sr(N__39568));
    defparam \pid_alt.pid_prereg_esr_RNIHKIA2_12_LC_4_12_0 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIHKIA2_12_LC_4_12_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIHKIA2_12_LC_4_12_0 .LUT_INIT=16'b1111011111110000;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIHKIA2_12_LC_4_12_0  (
            .in0(N__40218),
            .in1(N__39715),
            .in2(N__39785),
            .in3(N__39665),
            .lcout(\pid_alt.source_pid_9_0_tz_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIG2382_12_LC_4_12_1 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIG2382_12_LC_4_12_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIG2382_12_LC_4_12_1 .LUT_INIT=16'b0111011101010101;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIG2382_12_LC_4_12_1  (
            .in0(N__39714),
            .in1(N__40217),
            .in2(_gnd_net_),
            .in3(N__39244),
            .lcout(\pid_alt.N_52 ),
            .ltout(\pid_alt.N_52_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNI3BD63_4_LC_4_12_2 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNI3BD63_4_LC_4_12_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNI3BD63_4_LC_4_12_2 .LUT_INIT=16'b1111000011111010;
    LogicCell40 \pid_alt.pid_prereg_esr_RNI3BD63_4_LC_4_12_2  (
            .in0(N__40170),
            .in1(_gnd_net_),
            .in2(N__36622),
            .in3(N__39869),
            .lcout(\pid_alt.N_54 ),
            .ltout(\pid_alt.N_54_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.source_pid_1_esr_0_LC_4_12_3 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_0_LC_4_12_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_0_LC_4_12_3 .LUT_INIT=16'b1110110000000000;
    LogicCell40 \pid_alt.source_pid_1_esr_0_LC_4_12_3  (
            .in0(N__39666),
            .in1(N__39776),
            .in2(N__36874),
            .in3(N__36736),
            .lcout(throttle_order_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94272),
            .ce(N__39594),
            .sr(N__39556));
    defparam \pid_alt.source_pid_1_esr_1_LC_4_12_4 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_1_LC_4_12_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_1_LC_4_12_4 .LUT_INIT=16'b1010100010100000;
    LogicCell40 \pid_alt.source_pid_1_esr_1_LC_4_12_4  (
            .in0(N__36712),
            .in1(N__36827),
            .in2(N__39786),
            .in3(N__39668),
            .lcout(throttle_order_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94272),
            .ce(N__39594),
            .sr(N__39556));
    defparam \pid_alt.source_pid_1_esr_2_LC_4_12_5 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_2_LC_4_12_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_2_LC_4_12_5 .LUT_INIT=16'b1110110000000000;
    LogicCell40 \pid_alt.source_pid_1_esr_2_LC_4_12_5  (
            .in0(N__39667),
            .in1(N__39780),
            .in2(N__36832),
            .in3(N__37042),
            .lcout(throttle_order_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94272),
            .ce(N__39594),
            .sr(N__39556));
    defparam \pid_alt.source_pid_1_esr_3_LC_4_12_6 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_3_LC_4_12_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_3_LC_4_12_6 .LUT_INIT=16'b1110000010100000;
    LogicCell40 \pid_alt.source_pid_1_esr_3_LC_4_12_6  (
            .in0(N__39781),
            .in1(N__36831),
            .in2(N__36985),
            .in3(N__39669),
            .lcout(throttle_order_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94272),
            .ce(N__39594),
            .sr(N__39556));
    defparam \pid_alt.pid_prereg_esr_RNIQT5H1_0_LC_4_12_7 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIQT5H1_0_LC_4_12_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIQT5H1_0_LC_4_12_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIQT5H1_0_LC_4_12_7  (
            .in0(N__37041),
            .in1(N__36711),
            .in2(N__36984),
            .in3(N__36735),
            .lcout(\pid_alt.source_pid_1_sqmuxa_0_a2_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_4_13_0 .C_ON=1'b1;
    defparam \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_4_13_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_4_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_4_13_0  (
            .in0(_gnd_net_),
            .in1(N__36795),
            .in2(N__36802),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_13_0_),
            .carryout(\pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_0_LC_4_13_1 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_0_LC_4_13_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_0_LC_4_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_0_LC_4_13_1  (
            .in0(_gnd_net_),
            .in1(N__36775),
            .in2(N__36763),
            .in3(N__36727),
            .lcout(\pid_alt.pid_preregZ0Z_0 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CO ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_0 ),
            .clk(N__94288),
            .ce(N__40511),
            .sr(N__86485));
    defparam \pid_alt.pid_prereg_esr_1_LC_4_13_2 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_1_LC_4_13_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_1_LC_4_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_1_LC_4_13_2  (
            .in0(_gnd_net_),
            .in1(N__36724),
            .in2(N__38866),
            .in3(N__36703),
            .lcout(\pid_alt.pid_preregZ0Z_1 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_0 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_1 ),
            .clk(N__94288),
            .ce(N__40511),
            .sr(N__86485));
    defparam \pid_alt.pid_prereg_esr_2_LC_4_13_3 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_2_LC_4_13_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_2_LC_4_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_2_LC_4_13_3  (
            .in0(_gnd_net_),
            .in1(N__37084),
            .in2(N__37075),
            .in3(N__37030),
            .lcout(\pid_alt.pid_preregZ0Z_2 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_1 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_2 ),
            .clk(N__94288),
            .ce(N__40511),
            .sr(N__86485));
    defparam \pid_alt.pid_prereg_esr_3_LC_4_13_4 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_3_LC_4_13_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_3_LC_4_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_3_LC_4_13_4  (
            .in0(_gnd_net_),
            .in1(N__37027),
            .in2(N__37021),
            .in3(N__36967),
            .lcout(\pid_alt.pid_preregZ0Z_3 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_2 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_3 ),
            .clk(N__94288),
            .ce(N__40511),
            .sr(N__86485));
    defparam \pid_alt.pid_prereg_esr_4_LC_4_13_5 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_4_LC_4_13_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_4_LC_4_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_4_LC_4_13_5  (
            .in0(_gnd_net_),
            .in1(N__36957),
            .in2(N__36946),
            .in3(N__36937),
            .lcout(\pid_alt.pid_preregZ0Z_4 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_3 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_4 ),
            .clk(N__94288),
            .ce(N__40511),
            .sr(N__86485));
    defparam \pid_alt.pid_prereg_esr_5_LC_4_13_6 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_5_LC_4_13_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_5_LC_4_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_5_LC_4_13_6  (
            .in0(_gnd_net_),
            .in1(N__36934),
            .in2(N__36928),
            .in3(N__36913),
            .lcout(\pid_alt.pid_preregZ0Z_5 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_4 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_5 ),
            .clk(N__94288),
            .ce(N__40511),
            .sr(N__86485));
    defparam \pid_alt.pid_prereg_esr_6_LC_4_13_7 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_6_LC_4_13_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_6_LC_4_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_6_LC_4_13_7  (
            .in0(_gnd_net_),
            .in1(N__36910),
            .in2(N__36903),
            .in3(N__36886),
            .lcout(\pid_alt.pid_preregZ0Z_6 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_5 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_6 ),
            .clk(N__94288),
            .ce(N__40511),
            .sr(N__86485));
    defparam \pid_alt.pid_prereg_esr_7_LC_4_14_0 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_7_LC_4_14_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_7_LC_4_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_7_LC_4_14_0  (
            .in0(_gnd_net_),
            .in1(N__39931),
            .in2(N__39993),
            .in3(N__36883),
            .lcout(\pid_alt.pid_preregZ0Z_7 ),
            .ltout(),
            .carryin(bfn_4_14_0_),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_7 ),
            .clk(N__94303),
            .ce(N__40508),
            .sr(N__86478));
    defparam \pid_alt.pid_prereg_esr_8_LC_4_14_1 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_8_LC_4_14_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_8_LC_4_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_8_LC_4_14_1  (
            .in0(_gnd_net_),
            .in1(N__39523),
            .in2(N__40078),
            .in3(N__36880),
            .lcout(\pid_alt.pid_preregZ0Z_8 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_7 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_8 ),
            .clk(N__94303),
            .ce(N__40508),
            .sr(N__86478));
    defparam \pid_alt.pid_prereg_esr_9_LC_4_14_2 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_9_LC_4_14_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_9_LC_4_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_9_LC_4_14_2  (
            .in0(_gnd_net_),
            .in1(N__37711),
            .in2(N__39402),
            .in3(N__36877),
            .lcout(\pid_alt.pid_preregZ0Z_9 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_8 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_9 ),
            .clk(N__94303),
            .ce(N__40508),
            .sr(N__86478));
    defparam \pid_alt.pid_prereg_esr_10_LC_4_14_3 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_10_LC_4_14_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_10_LC_4_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_10_LC_4_14_3  (
            .in0(_gnd_net_),
            .in1(N__37336),
            .in2(N__37668),
            .in3(N__37324),
            .lcout(\pid_alt.pid_preregZ0Z_10 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_9 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_10 ),
            .clk(N__94303),
            .ce(N__40508),
            .sr(N__86478));
    defparam \pid_alt.pid_prereg_esr_11_LC_4_14_4 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_11_LC_4_14_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_11_LC_4_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_11_LC_4_14_4  (
            .in0(_gnd_net_),
            .in1(N__37321),
            .in2(N__37309),
            .in3(N__37285),
            .lcout(\pid_alt.pid_preregZ0Z_11 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_10 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_11 ),
            .clk(N__94303),
            .ce(N__40508),
            .sr(N__86478));
    defparam \pid_alt.pid_prereg_esr_12_LC_4_14_5 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_12_LC_4_14_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_12_LC_4_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_12_LC_4_14_5  (
            .in0(_gnd_net_),
            .in1(N__37282),
            .in2(N__37276),
            .in3(N__37249),
            .lcout(\pid_alt.pid_preregZ0Z_12 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_11 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_12 ),
            .clk(N__94303),
            .ce(N__40508),
            .sr(N__86478));
    defparam \pid_alt.pid_prereg_esr_13_LC_4_14_6 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_13_LC_4_14_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_13_LC_4_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_13_LC_4_14_6  (
            .in0(_gnd_net_),
            .in1(N__37246),
            .in2(N__37239),
            .in3(N__37222),
            .lcout(\pid_alt.pid_preregZ0Z_13 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_12 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_13 ),
            .clk(N__94303),
            .ce(N__40508),
            .sr(N__86478));
    defparam \pid_alt.pid_prereg_esr_14_LC_4_14_7 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_14_LC_4_14_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_14_LC_4_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_14_LC_4_14_7  (
            .in0(_gnd_net_),
            .in1(N__37219),
            .in2(N__37210),
            .in3(N__37195),
            .lcout(\pid_alt.pid_preregZ0Z_14 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_13 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_14 ),
            .clk(N__94303),
            .ce(N__40508),
            .sr(N__86478));
    defparam \pid_alt.pid_prereg_esr_15_LC_4_15_0 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_15_LC_4_15_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_15_LC_4_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_15_LC_4_15_0  (
            .in0(_gnd_net_),
            .in1(N__37192),
            .in2(N__37182),
            .in3(N__37165),
            .lcout(\pid_alt.pid_preregZ0Z_15 ),
            .ltout(),
            .carryin(bfn_4_15_0_),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_15 ),
            .clk(N__94321),
            .ce(N__40504),
            .sr(N__86468));
    defparam \pid_alt.pid_prereg_esr_16_LC_4_15_1 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_16_LC_4_15_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_16_LC_4_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_16_LC_4_15_1  (
            .in0(_gnd_net_),
            .in1(N__37162),
            .in2(N__37143),
            .in3(N__37126),
            .lcout(\pid_alt.pid_preregZ0Z_16 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_15 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_16 ),
            .clk(N__94321),
            .ce(N__40504),
            .sr(N__86468));
    defparam \pid_alt.pid_prereg_esr_17_LC_4_15_2 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_17_LC_4_15_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_17_LC_4_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_17_LC_4_15_2  (
            .in0(_gnd_net_),
            .in1(N__37123),
            .in2(N__37102),
            .in3(N__37087),
            .lcout(\pid_alt.pid_preregZ0Z_17 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_16 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_17 ),
            .clk(N__94321),
            .ce(N__40504),
            .sr(N__86468));
    defparam \pid_alt.pid_prereg_esr_18_LC_4_15_3 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_18_LC_4_15_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_18_LC_4_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_18_LC_4_15_3  (
            .in0(_gnd_net_),
            .in1(N__37579),
            .in2(N__37567),
            .in3(N__37540),
            .lcout(\pid_alt.pid_preregZ0Z_18 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_17 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_18 ),
            .clk(N__94321),
            .ce(N__40504),
            .sr(N__86468));
    defparam \pid_alt.pid_prereg_esr_19_LC_4_15_4 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_19_LC_4_15_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_19_LC_4_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_19_LC_4_15_4  (
            .in0(_gnd_net_),
            .in1(N__37537),
            .in2(N__37528),
            .in3(N__37507),
            .lcout(\pid_alt.pid_preregZ0Z_19 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_18 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_19 ),
            .clk(N__94321),
            .ce(N__40504),
            .sr(N__86468));
    defparam \pid_alt.pid_prereg_esr_20_LC_4_15_5 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_20_LC_4_15_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_20_LC_4_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_20_LC_4_15_5  (
            .in0(_gnd_net_),
            .in1(N__37504),
            .in2(N__37495),
            .in3(N__37477),
            .lcout(\pid_alt.pid_preregZ0Z_20 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_19 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_20 ),
            .clk(N__94321),
            .ce(N__40504),
            .sr(N__86468));
    defparam \pid_alt.pid_prereg_esr_21_LC_4_15_6 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_21_LC_4_15_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_21_LC_4_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_21_LC_4_15_6  (
            .in0(_gnd_net_),
            .in1(N__37474),
            .in2(N__37462),
            .in3(N__37450),
            .lcout(\pid_alt.pid_preregZ0Z_21 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_20 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_21 ),
            .clk(N__94321),
            .ce(N__40504),
            .sr(N__86468));
    defparam \pid_alt.pid_prereg_esr_22_LC_4_15_7 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_22_LC_4_15_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_22_LC_4_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_22_LC_4_15_7  (
            .in0(_gnd_net_),
            .in1(N__37447),
            .in2(N__37432),
            .in3(N__37435),
            .lcout(\pid_alt.pid_preregZ0Z_22 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_21 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_22 ),
            .clk(N__94321),
            .ce(N__40504),
            .sr(N__86468));
    defparam \pid_alt.pid_prereg_esr_23_LC_4_16_0 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_23_LC_4_16_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_23_LC_4_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_23_LC_4_16_0  (
            .in0(_gnd_net_),
            .in1(N__37431),
            .in2(N__37405),
            .in3(N__37390),
            .lcout(\pid_alt.pid_preregZ0Z_23 ),
            .ltout(),
            .carryin(bfn_4_16_0_),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_23 ),
            .clk(N__94336),
            .ce(N__40502),
            .sr(N__86464));
    defparam \pid_alt.pid_prereg_esr_24_LC_4_16_1 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_24_LC_4_16_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_24_LC_4_16_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_alt.pid_prereg_esr_24_LC_4_16_1  (
            .in0(_gnd_net_),
            .in1(N__37387),
            .in2(_gnd_net_),
            .in3(N__37375),
            .lcout(\pid_alt.pid_preregZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94336),
            .ce(N__40502),
            .sr(N__86464));
    defparam \pid_alt.error_i_acumm_prereg_esr_14_LC_4_16_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_14_LC_4_16_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_14_LC_4_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_14_LC_4_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37372),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94336),
            .ce(N__40502),
            .sr(N__86464));
    defparam \pid_alt.error_i_acumm_prereg_esr_6_LC_4_16_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_6_LC_4_16_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_6_LC_4_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_6_LC_4_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37765),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94336),
            .ce(N__40502),
            .sr(N__86464));
    defparam \pid_alt.error_i_acumm_prereg_esr_19_LC_4_16_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_19_LC_4_16_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_19_LC_4_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_19_LC_4_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37744),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94336),
            .ce(N__40502),
            .sr(N__86464));
    defparam \pid_alt.error_d_reg_prev_esr_RNIN49Q5_8_LC_4_17_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIN49Q5_8_LC_4_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIN49Q5_8_LC_4_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIN49Q5_8_LC_4_17_0  (
            .in0(N__37678),
            .in1(N__37644),
            .in2(N__39406),
            .in3(N__37592),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIN49Q5Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIL8611_0_9_LC_4_17_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIL8611_0_9_LC_4_17_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIL8611_0_9_LC_4_17_1 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIL8611_0_9_LC_4_17_1  (
            .in0(N__37702),
            .in1(N__37605),
            .in2(_gnd_net_),
            .in3(N__37634),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIG75T2_8_LC_4_17_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIG75T2_8_LC_4_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIG75T2_8_LC_4_17_2 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIG75T2_8_LC_4_17_2  (
            .in0(_gnd_net_),
            .in1(N__37645),
            .in2(N__37672),
            .in3(N__37593),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIG75T2Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNII5611_8_LC_4_17_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNII5611_8_LC_4_17_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNII5611_8_LC_4_17_3 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNII5611_8_LC_4_17_3  (
            .in0(N__39516),
            .in1(N__39486),
            .in2(_gnd_net_),
            .in3(N__39471),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNII5611Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_8_LC_4_17_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_8_LC_4_17_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_8_LC_4_17_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_8_LC_4_17_4  (
            .in0(N__39472),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94351),
            .ce(N__40500),
            .sr(N__86459));
    defparam \pid_alt.error_d_reg_prev_esr_9_LC_4_17_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_9_LC_4_17_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_9_LC_4_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_9_LC_4_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37635),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94351),
            .ce(N__40500),
            .sr(N__86459));
    defparam \pid_alt.error_i_acumm_prereg_esr_9_LC_4_17_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_9_LC_4_17_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_9_LC_4_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_9_LC_4_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37594),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94351),
            .ce(N__40500),
            .sr(N__86459));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIPNRC1_11_LC_4_17_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIPNRC1_11_LC_4_17_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIPNRC1_11_LC_4_17_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNIPNRC1_11_LC_4_17_7  (
            .in0(N__38123),
            .in1(N__38107),
            .in2(N__38082),
            .in3(N__38675),
            .lcout(\pid_alt.m21_e_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_0_c_LC_4_18_0 .C_ON=1'b1;
    defparam \pid_alt.error_cry_0_c_LC_4_18_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_0_c_LC_4_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_alt.error_cry_0_c_LC_4_18_0  (
            .in0(_gnd_net_),
            .in1(N__46231),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_18_0_),
            .carryout(\pid_alt.error_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_0_c_RNI1N2F_LC_4_18_1 .C_ON=1'b1;
    defparam \pid_alt.error_cry_0_c_RNI1N2F_LC_4_18_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_0_c_RNI1N2F_LC_4_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_cry_0_c_RNI1N2F_LC_4_18_1  (
            .in0(_gnd_net_),
            .in1(N__48430),
            .in2(_gnd_net_),
            .in3(N__37996),
            .lcout(\pid_alt.error_1 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_0 ),
            .carryout(\pid_alt.error_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_1_c_RNI3Q3F_LC_4_18_2 .C_ON=1'b1;
    defparam \pid_alt.error_cry_1_c_RNI3Q3F_LC_4_18_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_1_c_RNI3Q3F_LC_4_18_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_cry_1_c_RNI3Q3F_LC_4_18_2  (
            .in0(_gnd_net_),
            .in1(N__52300),
            .in2(_gnd_net_),
            .in3(N__37954),
            .lcout(\pid_alt.error_2 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_1 ),
            .carryout(\pid_alt.error_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_2_c_RNI5T4F_LC_4_18_3 .C_ON=1'b1;
    defparam \pid_alt.error_cry_2_c_RNI5T4F_LC_4_18_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_2_c_RNI5T4F_LC_4_18_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_cry_2_c_RNI5T4F_LC_4_18_3  (
            .in0(_gnd_net_),
            .in1(N__52285),
            .in2(_gnd_net_),
            .in3(N__37906),
            .lcout(\pid_alt.error_3 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_2 ),
            .carryout(\pid_alt.error_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_3_c_RNIKE1T_LC_4_18_4 .C_ON=1'b1;
    defparam \pid_alt.error_cry_3_c_RNIKE1T_LC_4_18_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_3_c_RNIKE1T_LC_4_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_3_c_RNIKE1T_LC_4_18_4  (
            .in0(_gnd_net_),
            .in1(N__46162),
            .in2(N__40093),
            .in3(N__37858),
            .lcout(\pid_alt.error_4 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_3 ),
            .carryout(\pid_alt.error_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_4_c_RNINI2T_LC_4_18_5 .C_ON=1'b1;
    defparam \pid_alt.error_cry_4_c_RNINI2T_LC_4_18_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_4_c_RNINI2T_LC_4_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_4_c_RNINI2T_LC_4_18_5  (
            .in0(_gnd_net_),
            .in1(N__46153),
            .in2(N__40129),
            .in3(N__37813),
            .lcout(\pid_alt.error_5 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_4 ),
            .carryout(\pid_alt.error_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_5_c_RNIQM3T_LC_4_18_6 .C_ON=1'b1;
    defparam \pid_alt.error_cry_5_c_RNIQM3T_LC_4_18_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_5_c_RNIQM3T_LC_4_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_5_c_RNIQM3T_LC_4_18_6  (
            .in0(_gnd_net_),
            .in1(N__40363),
            .in2(N__46144),
            .in3(N__37768),
            .lcout(\pid_alt.error_6 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_5 ),
            .carryout(\pid_alt.error_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_6_c_RNITQ4T_LC_4_18_7 .C_ON=1'b1;
    defparam \pid_alt.error_cry_6_c_RNITQ4T_LC_4_18_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_6_c_RNITQ4T_LC_4_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_6_c_RNITQ4T_LC_4_18_7  (
            .in0(_gnd_net_),
            .in1(N__40104),
            .in2(N__46129),
            .in3(N__38509),
            .lcout(\pid_alt.error_7 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_6 ),
            .carryout(\pid_alt.error_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_7_c_RNI9LEM_LC_4_19_0 .C_ON=1'b1;
    defparam \pid_alt.error_cry_7_c_RNI9LEM_LC_4_19_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_7_c_RNI9LEM_LC_4_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_7_c_RNI9LEM_LC_4_19_0  (
            .in0(_gnd_net_),
            .in1(N__40303),
            .in2(N__40345),
            .in3(N__38464),
            .lcout(\pid_alt.error_8 ),
            .ltout(),
            .carryin(bfn_4_19_0_),
            .carryout(\pid_alt.error_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_8_c_RNICPFM_LC_4_19_1 .C_ON=1'b1;
    defparam \pid_alt.error_cry_8_c_RNICPFM_LC_4_19_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_8_c_RNICPFM_LC_4_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_8_c_RNICPFM_LC_4_19_1  (
            .in0(_gnd_net_),
            .in1(N__46375),
            .in2(N__40336),
            .in3(N__38419),
            .lcout(\pid_alt.error_9 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_8 ),
            .carryout(\pid_alt.error_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_9_c_RNIMMUJ_LC_4_19_2 .C_ON=1'b1;
    defparam \pid_alt.error_cry_9_c_RNIMMUJ_LC_4_19_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_9_c_RNIMMUJ_LC_4_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_9_c_RNIMMUJ_LC_4_19_2  (
            .in0(_gnd_net_),
            .in1(N__48640),
            .in2(N__40327),
            .in3(N__38374),
            .lcout(\pid_alt.error_10 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_9 ),
            .carryout(\pid_alt.error_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_10_c_RNI0SDO_LC_4_19_3 .C_ON=1'b1;
    defparam \pid_alt.error_cry_10_c_RNI0SDO_LC_4_19_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_10_c_RNI0SDO_LC_4_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_10_c_RNI0SDO_LC_4_19_3  (
            .in0(_gnd_net_),
            .in1(N__52483),
            .in2(N__40432),
            .in3(N__38326),
            .lcout(\pid_alt.error_11 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_10 ),
            .carryout(\pid_alt.error_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_11_c_RNI5JAH_LC_4_19_4 .C_ON=1'b1;
    defparam \pid_alt.error_cry_11_c_RNI5JAH_LC_4_19_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_11_c_RNI5JAH_LC_4_19_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_cry_11_c_RNI5JAH_LC_4_19_4  (
            .in0(_gnd_net_),
            .in1(N__48415),
            .in2(_gnd_net_),
            .in3(N__38278),
            .lcout(\pid_alt.error_12 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_11 ),
            .carryout(\pid_alt.error_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_12_c_RNI7MBH_LC_4_19_5 .C_ON=1'b1;
    defparam \pid_alt.error_cry_12_c_RNI7MBH_LC_4_19_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_12_c_RNI7MBH_LC_4_19_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_cry_12_c_RNI7MBH_LC_4_19_5  (
            .in0(_gnd_net_),
            .in1(N__52372),
            .in2(_gnd_net_),
            .in3(N__38230),
            .lcout(\pid_alt.error_13 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_12 ),
            .carryout(\pid_alt.error_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_13_c_RNI9PCH_LC_4_19_6 .C_ON=1'b1;
    defparam \pid_alt.error_cry_13_c_RNI9PCH_LC_4_19_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_13_c_RNI9PCH_LC_4_19_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_cry_13_c_RNI9PCH_LC_4_19_6  (
            .in0(_gnd_net_),
            .in1(N__52351),
            .in2(_gnd_net_),
            .in3(N__38185),
            .lcout(\pid_alt.error_14 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_13 ),
            .carryout(\pid_alt.error_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_14_c_RNIBSDH_LC_4_19_7 .C_ON=1'b0;
    defparam \pid_alt.error_cry_14_c_RNIBSDH_LC_4_19_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_14_c_RNIBSDH_LC_4_19_7 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \pid_alt.error_cry_14_c_RNIBSDH_LC_4_19_7  (
            .in0(N__48451),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38182),
            .lcout(\pid_alt.error_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_1_LC_4_20_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_1_LC_4_20_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_1_LC_4_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_1_LC_4_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38865),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94380),
            .ce(N__40497),
            .sr(N__86446));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI935T_0_LC_4_20_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI935T_0_LC_4_20_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI935T_0_LC_4_20_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNI935T_0_LC_4_20_1  (
            .in0(_gnd_net_),
            .in1(N__38823),
            .in2(_gnd_net_),
            .in3(N__38721),
            .lcout(),
            .ltout(\pid_alt.m21_e_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI57T82_7_LC_4_20_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI57T82_7_LC_4_20_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI57T82_7_LC_4_20_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNI57T82_7_LC_4_20_2  (
            .in0(N__38699),
            .in1(N__38580),
            .in2(N__38812),
            .in3(N__38804),
            .lcout(\pid_alt.m21_e_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_0_LC_4_20_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_0_LC_4_20_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_0_LC_4_20_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_0_LC_4_20_3  (
            .in0(_gnd_net_),
            .in1(N__38776),
            .in2(_gnd_net_),
            .in3(N__38743),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94380),
            .ce(N__40497),
            .sr(N__86446));
    defparam \pid_alt.error_i_acumm_prereg_esr_7_LC_4_20_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_7_LC_4_20_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_7_LC_4_20_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_7_LC_4_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39961),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94380),
            .ce(N__40497),
            .sr(N__86446));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNILF5T_6_LC_4_20_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNILF5T_6_LC_4_20_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNILF5T_6_LC_4_20_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNILF5T_6_LC_4_20_5  (
            .in0(_gnd_net_),
            .in1(N__38700),
            .in2(_gnd_net_),
            .in3(N__38682),
            .lcout(\pid_alt.m35_e_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_5_LC_4_20_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_5_LC_4_20_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_5_LC_4_20_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_5_LC_4_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38641),
            .lcout(\pid_alt.error_i_acumm7lto5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94380),
            .ce(N__40497),
            .sr(N__86446));
    defparam \pid_front.error_p_reg_esr_16_LC_4_23_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_16_LC_4_23_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_16_LC_4_23_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_16_LC_4_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38563),
            .lcout(\pid_front.error_p_regZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94399),
            .ce(N__93386),
            .sr(N__92987));
    defparam \ppm_encoder_1.PPM_STATE_fast_0_LC_5_1_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_fast_0_LC_5_1_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.PPM_STATE_fast_0_LC_5_1_2 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \ppm_encoder_1.PPM_STATE_fast_0_LC_5_1_2  (
            .in0(N__49741),
            .in1(N__49854),
            .in2(_gnd_net_),
            .in3(N__49783),
            .lcout(\ppm_encoder_1.PPM_STATE_fastZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94115),
            .ce(),
            .sr(N__86519));
    defparam \ppm_encoder_1.init_pulses_RNI70081_3_LC_5_2_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI70081_3_LC_5_2_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI70081_3_LC_5_2_0 .LUT_INIT=16'b1111000001111000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI70081_3_LC_5_2_0  (
            .in0(N__42197),
            .in1(N__43727),
            .in2(N__44851),
            .in3(N__52711),
            .lcout(\ppm_encoder_1.N_256_i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_3_LC_5_2_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_3_LC_5_2_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_3_LC_5_2_2 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \ppm_encoder_1.init_pulses_3_LC_5_2_2  (
            .in0(N__49390),
            .in1(N__41449),
            .in2(N__49504),
            .in3(N__43507),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94123),
            .ce(),
            .sr(N__86518));
    defparam \ppm_encoder_1.init_pulses_1_LC_5_2_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_1_LC_5_2_4 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_1_LC_5_2_4 .LUT_INIT=16'b0010001100100000;
    LogicCell40 \ppm_encoder_1.init_pulses_1_LC_5_2_4  (
            .in0(N__41488),
            .in1(N__49499),
            .in2(N__49395),
            .in3(N__43609),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94123),
            .ce(),
            .sr(N__86518));
    defparam \ppm_encoder_1.init_pulses_4_LC_5_2_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_4_LC_5_2_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_4_LC_5_2_6 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \ppm_encoder_1.init_pulses_4_LC_5_2_6  (
            .in0(N__49495),
            .in1(N__41428),
            .in2(N__49396),
            .in3(N__43975),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94123),
            .ce(),
            .sr(N__86518));
    defparam \ppm_encoder_1.init_pulses_RNIA2081_5_LC_5_2_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIA2081_5_LC_5_2_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIA2081_5_LC_5_2_7 .LUT_INIT=16'b1001110011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIA2081_5_LC_5_2_7  (
            .in0(N__52712),
            .in1(N__49967),
            .in2(N__43736),
            .in3(N__53695),
            .lcout(\ppm_encoder_1.N_261_i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI58QQ_3_LC_5_3_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI58QQ_3_LC_5_3_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI58QQ_3_LC_5_3_0 .LUT_INIT=16'b1111111111101011;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI58QQ_3_LC_5_3_0  (
            .in0(N__49765),
            .in1(N__41983),
            .in2(N__42206),
            .in3(N__49532),
            .lcout(\ppm_encoder_1.init_pulses_4_sqmuxa_i_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_1_LC_5_3_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_1_LC_5_3_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.PPM_STATE_1_LC_5_3_1 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \ppm_encoder_1.PPM_STATE_1_LC_5_3_1  (
            .in0(N__49533),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49733),
            .lcout(\ppm_encoder_1.PPM_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94131),
            .ce(),
            .sr(N__86517));
    defparam \ppm_encoder_1.PPM_STATE_fast_RNICIAB_0_LC_5_3_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_fast_RNICIAB_0_LC_5_3_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_fast_RNICIAB_0_LC_5_3_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \ppm_encoder_1.PPM_STATE_fast_RNICIAB_0_LC_5_3_3  (
            .in0(_gnd_net_),
            .in1(N__38878),
            .in2(_gnd_net_),
            .in3(N__49764),
            .lcout(\ppm_encoder_1.PPM_STATE_fast_RNICIABZ0Z_0 ),
            .ltout(\ppm_encoder_1.PPM_STATE_fast_RNICIABZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_RNI7E8E1_1_LC_5_3_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_RNI7E8E1_1_LC_5_3_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.aileron_RNI7E8E1_1_LC_5_3_4 .LUT_INIT=16'b1111110111111100;
    LogicCell40 \ppm_encoder_1.aileron_RNI7E8E1_1_LC_5_3_4  (
            .in0(N__50241),
            .in1(N__41984),
            .in2(N__38869),
            .in3(N__44593),
            .lcout(),
            .ltout(\ppm_encoder_1.aileron_RNI7E8E1Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNII4422_0_LC_5_3_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNII4422_0_LC_5_3_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNII4422_0_LC_5_3_5 .LUT_INIT=16'b1111101011111001;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNII4422_0_LC_5_3_5  (
            .in0(N__38953),
            .in1(N__38917),
            .in2(N__38968),
            .in3(N__38899),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNITALE4_1_LC_5_3_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNITALE4_1_LC_5_3_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNITALE4_1_LC_5_3_6 .LUT_INIT=16'b1001100110010110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNITALE4_1_LC_5_3_6  (
            .in0(N__40411),
            .in1(N__41788),
            .in2(N__38965),
            .in3(N__38962),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_0_axb_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI29LM5_1_LC_5_3_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI29LM5_1_LC_5_3_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI29LM5_1_LC_5_3_7 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI29LM5_1_LC_5_3_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38956),
            .in3(N__43626),
            .lcout(\ppm_encoder_1.init_pulses_RNI29LM5Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_2_LC_5_4_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_2_LC_5_4_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_2_LC_5_4_0 .LUT_INIT=16'b0100010000000101;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_2_LC_5_4_0  (
            .in0(N__71046),
            .in1(N__38950),
            .in2(N__47149),
            .in3(N__52680),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94138),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_0_i_o2_LC_5_4_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_0_i_o2_LC_5_4_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_0_i_o2_LC_5_4_1 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_0_i_o2_LC_5_4_1  (
            .in0(_gnd_net_),
            .in1(N__38914),
            .in2(_gnd_net_),
            .in3(N__38896),
            .lcout(\ppm_encoder_1.N_300 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_0_LC_5_4_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_0_LC_5_4_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_0_LC_5_4_2 .LUT_INIT=16'b1111101011111100;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_0_LC_5_4_2  (
            .in0(N__38898),
            .in1(N__47193),
            .in2(N__71062),
            .in3(N__52679),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94138),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_1_LC_5_4_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_1_LC_5_4_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_1_LC_5_4_3 .LUT_INIT=16'b0000000010011100;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_1_LC_5_4_3  (
            .in0(N__52678),
            .in1(N__38916),
            .in2(N__54262),
            .in3(N__71051),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94138),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_3_LC_5_4_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_3_LC_5_4_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_3_LC_5_4_4 .LUT_INIT=16'b0100010000000101;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_3_LC_5_4_4  (
            .in0(N__71047),
            .in1(N__41982),
            .in2(N__46912),
            .in3(N__52681),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94138),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI6LFQ_0_LC_5_4_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI6LFQ_0_LC_5_4_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI6LFQ_0_LC_5_4_5 .LUT_INIT=16'b1111101011111001;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI6LFQ_0_LC_5_4_5  (
            .in0(N__38949),
            .in1(N__38915),
            .in2(N__41988),
            .in3(N__38897),
            .lcout(),
            .ltout(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI6LFQZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNII7Q51_0_LC_5_4_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNII7Q51_0_LC_5_4_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNII7Q51_0_LC_5_4_6 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNII7Q51_0_LC_5_4_6  (
            .in0(N__65792),
            .in1(_gnd_net_),
            .in2(N__38881),
            .in3(N__52677),
            .lcout(\ppm_encoder_1.N_303 ),
            .ltout(\ppm_encoder_1.N_303_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNI4HVB2_2_LC_5_4_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI4HVB2_2_LC_5_4_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI4HVB2_2_LC_5_4_7 .LUT_INIT=16'b1111110011111101;
    LogicCell40 \ppm_encoder_1.elevator_RNI4HVB2_2_LC_5_4_7  (
            .in0(N__40809),
            .in1(N__42179),
            .in2(N__39007),
            .in3(N__47354),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_RNIM1KQ_12_LC_5_5_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_RNIM1KQ_12_LC_5_5_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.rudder_RNIM1KQ_12_LC_5_5_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \ppm_encoder_1.rudder_RNIM1KQ_12_LC_5_5_1  (
            .in0(_gnd_net_),
            .in1(N__42452),
            .in2(_gnd_net_),
            .in3(N__42170),
            .lcout(),
            .ltout(\ppm_encoder_1.N_448_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNI0PME2_12_LC_5_5_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI0PME2_12_LC_5_5_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI0PME2_12_LC_5_5_2 .LUT_INIT=16'b1111101011111011;
    LogicCell40 \ppm_encoder_1.elevator_RNI0PME2_12_LC_5_5_2  (
            .in0(N__44457),
            .in1(N__47355),
            .in2(N__38998),
            .in3(N__38990),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_2_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_12_LC_5_5_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_12_LC_5_5_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_12_LC_5_5_3 .LUT_INIT=16'b1000100011111000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_12_LC_5_5_3  (
            .in0(N__47508),
            .in1(N__42453),
            .in2(N__38995),
            .in3(N__47357),
            .lcout(\ppm_encoder_1.pulses2count_9_0_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_12_LC_5_5_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_12_LC_5_5_4 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_12_LC_5_5_4 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.elevator_12_LC_5_5_4  (
            .in0(N__55705),
            .in1(N__47602),
            .in2(N__51368),
            .in3(N__38994),
            .lcout(\ppm_encoder_1.elevatorZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94150),
            .ce(),
            .sr(N__86512));
    defparam \ppm_encoder_1.elevator_RNI5IVB2_3_LC_5_5_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI5IVB2_3_LC_5_5_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI5IVB2_3_LC_5_5_5 .LUT_INIT=16'b1110111011111110;
    LogicCell40 \ppm_encoder_1.elevator_RNI5IVB2_3_LC_5_5_5  (
            .in0(N__42172),
            .in1(N__44458),
            .in2(N__47554),
            .in3(N__47356),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIGNSS4_3_LC_5_5_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIGNSS4_3_LC_5_5_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIGNSS4_3_LC_5_5_6 .LUT_INIT=16'b0110011001101001;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIGNSS4_3_LC_5_5_6  (
            .in0(N__44852),
            .in1(N__41760),
            .in2(N__38980),
            .in3(N__38977),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_0_axb_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNINNS46_3_LC_5_5_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNINNS46_3_LC_5_5_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNINNS46_3_LC_5_5_7 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNINNS46_3_LC_5_5_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38971),
            .in3(N__43524),
            .lcout(\ppm_encoder_1.init_pulses_RNINNS46Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI5UV71_1_LC_5_6_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI5UV71_1_LC_5_6_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI5UV71_1_LC_5_6_0 .LUT_INIT=16'b1111000001111000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI5UV71_1_LC_5_6_0  (
            .in0(N__43711),
            .in1(N__42162),
            .in2(N__40416),
            .in3(N__52764),
            .lcout(\ppm_encoder_1.N_258_i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIRS8E1_8_LC_5_6_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIRS8E1_8_LC_5_6_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIRS8E1_8_LC_5_6_1 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \ppm_encoder_1.throttle_RNIRS8E1_8_LC_5_6_1  (
            .in0(N__44574),
            .in1(N__45060),
            .in2(N__44668),
            .in3(N__44804),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_1_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIJK8E1_4_LC_5_6_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIJK8E1_4_LC_5_6_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIJK8E1_4_LC_5_6_2 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \ppm_encoder_1.throttle_RNIJK8E1_4_LC_5_6_2  (
            .in0(N__46741),
            .in1(N__44648),
            .in2(N__39043),
            .in3(N__44573),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI81081_4_LC_5_6_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI81081_4_LC_5_6_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI81081_4_LC_5_6_3 .LUT_INIT=16'b1001110011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI81081_4_LC_5_6_3  (
            .in0(N__52765),
            .in1(N__50008),
            .in2(N__42192),
            .in3(N__43712),
            .lcout(\ppm_encoder_1.N_260_i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI81081_0_4_LC_5_6_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI81081_0_4_LC_5_6_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI81081_0_4_LC_5_6_4 .LUT_INIT=16'b0000111110000111;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI81081_0_4_LC_5_6_4  (
            .in0(N__43713),
            .in1(N__42166),
            .in2(N__50013),
            .in3(N__52766),
            .lcout(),
            .ltout(\ppm_encoder_1.N_260_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI7SCD5_4_LC_5_6_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI7SCD5_4_LC_5_6_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI7SCD5_4_LC_5_6_5 .LUT_INIT=16'b1111000011100001;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI7SCD5_4_LC_5_6_5  (
            .in0(N__39022),
            .in1(N__40723),
            .in2(N__39016),
            .in3(N__44467),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_0_axb_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIFTCL6_4_LC_5_6_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIFTCL6_4_LC_5_6_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIFTCL6_4_LC_5_6_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIFTCL6_4_LC_5_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__39013),
            .in3(N__43986),
            .lcout(\ppm_encoder_1.init_pulses_RNIFTCL6Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_LC_5_6_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_LC_5_6_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_LC_5_6_7 .LUT_INIT=16'b0000000010110001;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_LC_5_6_7  (
            .in0(N__52767),
            .in1(N__47142),
            .in2(N__42193),
            .in3(N__71017),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94161),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNICE0O2_9_LC_5_7_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNICE0O2_9_LC_5_7_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNICE0O2_9_LC_5_7_0 .LUT_INIT=16'b1110111011111110;
    LogicCell40 \ppm_encoder_1.elevator_RNICE0O2_9_LC_5_7_0  (
            .in0(N__39088),
            .in1(N__44478),
            .in2(N__44716),
            .in3(N__47431),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_2_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI96U85_9_LC_5_7_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI96U85_9_LC_5_7_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI96U85_9_LC_5_7_1 .LUT_INIT=16'b0110011001101001;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI96U85_9_LC_5_7_1  (
            .in0(N__46527),
            .in1(N__41776),
            .in2(N__39010),
            .in3(N__39082),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_0_axb_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIOCUG6_9_LC_5_7_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIOCUG6_9_LC_5_7_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIOCUG6_9_LC_5_7_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIOCUG6_9_LC_5_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__39091),
            .in3(N__43845),
            .lcout(\ppm_encoder_1.init_pulses_RNIOCUG6Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_RNICQ7Q_9_LC_5_7_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_RNICQ7Q_9_LC_5_7_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.rudder_RNICQ7Q_9_LC_5_7_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ppm_encoder_1.rudder_RNICQ7Q_9_LC_5_7_3  (
            .in0(_gnd_net_),
            .in1(N__46962),
            .in2(_gnd_net_),
            .in3(N__42171),
            .lcout(\ppm_encoder_1.N_454 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNITU8E1_9_LC_5_7_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNITU8E1_9_LC_5_7_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNITU8E1_9_LC_5_7_4 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \ppm_encoder_1.throttle_RNITU8E1_9_LC_5_7_4  (
            .in0(N__44758),
            .in1(N__44681),
            .in2(N__44986),
            .in3(N__44597),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_1_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIV7N11_13_LC_5_8_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIV7N11_13_LC_5_8_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIV7N11_13_LC_5_8_6 .LUT_INIT=16'b0010001011000000;
    LogicCell40 \ppm_encoder_1.throttle_RNIV7N11_13_LC_5_8_6  (
            .in0(N__51402),
            .in1(N__44907),
            .in2(N__39075),
            .in3(N__42089),
            .lcout(\ppm_encoder_1.un2_throttle_0_2_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.source_data_valid_esr_LC_5_10_0 .C_ON=1'b0;
    defparam \pid_alt.source_data_valid_esr_LC_5_10_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_data_valid_esr_LC_5_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.source_data_valid_esr_LC_5_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69011),
            .lcout(pid_altitude_dv),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94220),
            .ce(N__40144),
            .sr(N__86496));
    defparam \pid_alt.source_pid_1_esr_12_LC_5_11_0 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_12_LC_5_11_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_12_LC_5_11_0 .LUT_INIT=16'b1100010011000000;
    LogicCell40 \pid_alt.source_pid_1_esr_12_LC_5_11_0  (
            .in0(N__39723),
            .in1(N__40219),
            .in2(N__39787),
            .in3(N__39676),
            .lcout(throttle_order_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94237),
            .ce(N__39593),
            .sr(N__39566));
    defparam \pid_alt.pid_prereg_esr_RNIP29I1_4_LC_5_12_0 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIP29I1_4_LC_5_12_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIP29I1_4_LC_5_12_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIP29I1_4_LC_5_12_0  (
            .in0(N__39868),
            .in1(N__68958),
            .in2(N__39724),
            .in3(N__40163),
            .lcout(),
            .ltout(\pid_alt.source_pid_1_sqmuxa_0_a2_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIVVFP6_4_LC_5_12_1 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIVVFP6_4_LC_5_12_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIVVFP6_4_LC_5_12_1 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIVVFP6_4_LC_5_12_1  (
            .in0(N__39228),
            .in1(N__39243),
            .in2(N__39058),
            .in3(N__39663),
            .lcout(),
            .ltout(\pid_alt.N_57_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNI4AMM7_24_LC_5_12_2 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNI4AMM7_24_LC_5_12_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNI4AMM7_24_LC_5_12_2 .LUT_INIT=16'b0000000100000101;
    LogicCell40 \pid_alt.pid_prereg_esr_RNI4AMM7_24_LC_5_12_2  (
            .in0(N__70838),
            .in1(N__39772),
            .in2(N__39055),
            .in3(N__68959),
            .lcout(),
            .ltout(\pid_alt.un1_reset_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNI3A6GE_13_LC_5_12_3 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNI3A6GE_13_LC_5_12_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNI3A6GE_13_LC_5_12_3 .LUT_INIT=16'b0100111100001111;
    LogicCell40 \pid_alt.pid_prereg_esr_RNI3A6GE_13_LC_5_12_3  (
            .in0(N__39722),
            .in1(N__39214),
            .in2(N__39052),
            .in3(N__39664),
            .lcout(\pid_alt.un1_reset_0_i ),
            .ltout(\pid_alt.un1_reset_0_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.state_RNIOVDUE_1_LC_5_12_4 .C_ON=1'b0;
    defparam \pid_alt.state_RNIOVDUE_1_LC_5_12_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.state_RNIOVDUE_1_LC_5_12_4 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \pid_alt.state_RNIOVDUE_1_LC_5_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__39376),
            .in3(N__68960),
            .lcout(\pid_alt.N_72_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIIM6H1_6_LC_5_12_5 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIIM6H1_6_LC_5_12_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIIM6H1_6_LC_5_12_5 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIIM6H1_6_LC_5_12_5  (
            .in0(N__39371),
            .in1(N__39350),
            .in2(N__39330),
            .in3(N__39297),
            .lcout(),
            .ltout(\pid_alt.source_pid_1_sqmuxa_0_o2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIFQKS1_10_LC_5_12_6 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIFQKS1_10_LC_5_12_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIFQKS1_10_LC_5_12_6 .LUT_INIT=16'b1111001111111111;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIFQKS1_10_LC_5_12_6  (
            .in0(_gnd_net_),
            .in1(N__39284),
            .in2(N__39268),
            .in3(N__39263),
            .lcout(\pid_alt.N_51 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIHMCQ4_4_LC_5_12_7 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIHMCQ4_4_LC_5_12_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIHMCQ4_4_LC_5_12_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIHMCQ4_4_LC_5_12_7  (
            .in0(N__40162),
            .in1(N__39867),
            .in2(N__39232),
            .in3(N__39220),
            .lcout(\pid_alt.source_pid_1_sqmuxa_0_a2_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNICSUM_17_LC_5_13_0 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNICSUM_17_LC_5_13_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNICSUM_17_LC_5_13_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_alt.pid_prereg_esr_RNICSUM_17_LC_5_13_0  (
            .in0(N__39208),
            .in1(N__39196),
            .in2(N__39187),
            .in3(N__39172),
            .lcout(\pid_alt.source_pid_1_sqmuxa_0_a2_2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIBRUM_15_LC_5_13_1 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIBRUM_15_LC_5_13_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIBRUM_15_LC_5_13_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIBRUM_15_LC_5_13_1  (
            .in0(N__39163),
            .in1(N__39154),
            .in2(N__39145),
            .in3(N__39130),
            .lcout(),
            .ltout(\pid_alt.source_pid_1_sqmuxa_0_a2_2_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIT4CP1_14_LC_5_13_2 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIT4CP1_14_LC_5_13_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIT4CP1_14_LC_5_13_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIT4CP1_14_LC_5_13_2  (
            .in0(N__39121),
            .in1(N__39109),
            .in2(N__39103),
            .in3(N__39100),
            .lcout(\pid_alt.N_539 ),
            .ltout(\pid_alt.N_539_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.source_pid_1_esr_RNO_0_4_LC_5_13_3 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_RNO_0_4_LC_5_13_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.source_pid_1_esr_RNO_0_4_LC_5_13_3 .LUT_INIT=16'b0101010001000100;
    LogicCell40 \pid_alt.source_pid_1_esr_RNO_0_4_LC_5_13_3  (
            .in0(N__39870),
            .in1(N__39766),
            .in2(N__39094),
            .in3(N__40171),
            .lcout(),
            .ltout(\pid_alt.source_pid_9_0_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.source_pid_1_esr_4_LC_5_13_4 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_4_LC_5_13_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_4_LC_5_13_4 .LUT_INIT=16'b0000110100001111;
    LogicCell40 \pid_alt.source_pid_1_esr_4_LC_5_13_4  (
            .in0(N__39822),
            .in1(N__39871),
            .in2(N__39847),
            .in3(N__39675),
            .lcout(throttle_order_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94273),
            .ce(N__39604),
            .sr(N__39567));
    defparam \pid_alt.source_pid_1_esr_5_LC_5_13_5 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_5_LC_5_13_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_5_LC_5_13_5 .LUT_INIT=16'b1110000011000000;
    LogicCell40 \pid_alt.source_pid_1_esr_5_LC_5_13_5  (
            .in0(N__39673),
            .in1(N__39768),
            .in2(N__40191),
            .in3(N__39823),
            .lcout(throttle_order_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94273),
            .ce(N__39604),
            .sr(N__39567));
    defparam \pid_alt.source_pid_1_esr_13_LC_5_13_6 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_13_LC_5_13_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_13_LC_5_13_6 .LUT_INIT=16'b1100110011011101;
    LogicCell40 \pid_alt.source_pid_1_esr_13_LC_5_13_6  (
            .in0(N__39767),
            .in1(N__39707),
            .in2(_gnd_net_),
            .in3(N__39674),
            .lcout(throttle_order_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94273),
            .ce(N__39604),
            .sr(N__39567));
    defparam \pid_alt.error_d_reg_prev_esr_RNI5G6Q5_7_LC_5_14_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI5G6Q5_7_LC_5_14_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI5G6Q5_7_LC_5_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI5G6Q5_7_LC_5_14_0  (
            .in0(N__39442),
            .in1(N__39384),
            .in2(N__40077),
            .in3(N__39431),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI5G6Q5Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNII5611_0_8_LC_5_14_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNII5611_0_8_LC_5_14_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNII5611_0_8_LC_5_14_1 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNII5611_0_8_LC_5_14_1  (
            .in0(N__39517),
            .in1(N__39487),
            .in2(_gnd_net_),
            .in3(N__39465),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNII5611_0Z0Z_8 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNII5611_0Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI7T3T2_7_LC_5_14_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI7T3T2_7_LC_5_14_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI7T3T2_7_LC_5_14_2 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI7T3T2_7_LC_5_14_2  (
            .in0(_gnd_net_),
            .in1(N__39385),
            .in2(N__39436),
            .in3(N__39432),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI7T3T2Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIF2611_7_LC_5_14_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIF2611_7_LC_5_14_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIF2611_7_LC_5_14_3 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIF2611_7_LC_5_14_3  (
            .in0(N__40020),
            .in1(N__40029),
            .in2(_gnd_net_),
            .in3(N__40055),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIF2611Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_7_LC_5_14_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_7_LC_5_14_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_7_LC_5_14_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_7_LC_5_14_4  (
            .in0(N__40057),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94289),
            .ce(N__40505),
            .sr(N__86469));
    defparam \pid_alt.error_d_reg_prev_esr_RNIUI2T2_6_LC_5_14_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIUI2T2_6_LC_5_14_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIUI2T2_6_LC_5_14_5 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIUI2T2_6_LC_5_14_5  (
            .in0(N__40000),
            .in1(N__39976),
            .in2(_gnd_net_),
            .in3(N__39957),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIUI2T2Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIF2611_0_7_LC_5_14_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIF2611_0_7_LC_5_14_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIF2611_0_7_LC_5_14_6 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIF2611_0_7_LC_5_14_6  (
            .in0(N__40056),
            .in1(_gnd_net_),
            .in2(N__40033),
            .in3(N__40021),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIF2611_0Z0Z_7 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIF2611_0Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIJR3Q5_6_LC_5_14_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIJR3Q5_6_LC_5_14_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIJR3Q5_6_LC_5_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIJR3Q5_6_LC_5_14_7  (
            .in0(N__39994),
            .in1(N__39975),
            .in2(N__39964),
            .in3(N__39956),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIJR3Q5Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_17_LC_5_15_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_17_LC_5_15_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_17_LC_5_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_17_LC_5_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39922),
            .lcout(\pid_front.error_p_regZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94304),
            .ce(N__93316),
            .sr(N__92974));
    defparam \pid_front.error_p_reg_esr_3_LC_5_15_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_3_LC_5_15_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_3_LC_5_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_3_LC_5_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39907),
            .lcout(\pid_front.error_p_regZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94304),
            .ce(N__93316),
            .sr(N__92974));
    defparam \pid_front.error_p_reg_esr_7_LC_5_15_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_7_LC_5_15_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_7_LC_5_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_7_LC_5_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39898),
            .lcout(\pid_front.error_p_regZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94304),
            .ce(N__93316),
            .sr(N__92974));
    defparam \pid_front.error_p_reg_esr_8_LC_5_15_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_8_LC_5_15_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_8_LC_5_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_8_LC_5_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39886),
            .lcout(\pid_front.error_p_regZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94304),
            .ce(N__93316),
            .sr(N__92974));
    defparam \uart_pc.state_1_LC_5_16_0 .C_ON=1'b0;
    defparam \uart_pc.state_1_LC_5_16_0 .SEQ_MODE=4'b1000;
    defparam \uart_pc.state_1_LC_5_16_0 .LUT_INIT=16'b0000000011001000;
    LogicCell40 \uart_pc.state_1_LC_5_16_0  (
            .in0(N__41019),
            .in1(N__52242),
            .in2(N__41182),
            .in3(N__70938),
            .lcout(\uart_pc.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94322),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc_sync.aux_1__0__0_LC_5_16_4 .C_ON=1'b0;
    defparam \uart_pc_sync.aux_1__0__0_LC_5_16_4 .SEQ_MODE=4'b1000;
    defparam \uart_pc_sync.aux_1__0__0_LC_5_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_pc_sync.aux_1__0__0_LC_5_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40225),
            .lcout(\uart_pc_sync.aux_1__0_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94322),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc_sync.aux_0__0__0_LC_5_16_5 .C_ON=1'b0;
    defparam \uart_pc_sync.aux_0__0__0_LC_5_16_5 .SEQ_MODE=4'b1000;
    defparam \uart_pc_sync.aux_0__0__0_LC_5_16_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart_pc_sync.aux_0__0__0_LC_5_16_5  (
            .in0(N__40246),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uart_pc_sync.aux_0__0_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94322),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIIM0I_5_LC_5_16_6 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIIM0I_5_LC_5_16_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIIM0I_5_LC_5_16_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIIM0I_5_LC_5_16_6  (
            .in0(_gnd_net_),
            .in1(N__40216),
            .in2(_gnd_net_),
            .in3(N__40192),
            .lcout(\pid_alt.N_154 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.source_data_valid_esr_RNO_LC_5_16_7 .C_ON=1'b0;
    defparam \pid_alt.source_data_valid_esr_RNO_LC_5_16_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.source_data_valid_esr_RNO_LC_5_16_7 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \pid_alt.source_data_valid_esr_RNO_LC_5_16_7  (
            .in0(_gnd_net_),
            .in1(N__69078),
            .in2(_gnd_net_),
            .in3(N__86583),
            .lcout(\pid_alt.state_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH1data8lto7_LC_5_17_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data8lto7_LC_5_17_0 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.source_CH1data8lto7_LC_5_17_0 .LUT_INIT=16'b0001000011110000;
    LogicCell40 \Commands_frame_decoder.source_CH1data8lto7_LC_5_17_0  (
            .in0(N__85480),
            .in1(N__92431),
            .in2(N__40114),
            .in3(N__92234),
            .lcout(\Commands_frame_decoder.source_CH1data8 ),
            .ltout(\Commands_frame_decoder.source_CH1data8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH1data_1_LC_5_17_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_1_LC_5_17_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_1_LC_5_17_1 .LUT_INIT=16'b0000110010101010;
    LogicCell40 \Commands_frame_decoder.source_CH1data_1_LC_5_17_1  (
            .in0(N__40128),
            .in1(N__85481),
            .in2(N__40132),
            .in3(N__52461),
            .lcout(alt_command_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94337),
            .ce(),
            .sr(N__86454));
    defparam \Commands_frame_decoder.source_CH1data8lto7_2_LC_5_17_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data8lto7_2_LC_5_17_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.source_CH1data8lto7_2_LC_5_17_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Commands_frame_decoder.source_CH1data8lto7_2_LC_5_17_2  (
            .in0(N__88798),
            .in1(N__88641),
            .in2(N__92101),
            .in3(N__88425),
            .lcout(\Commands_frame_decoder.source_CH1data8lto7Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH1data_3_LC_5_17_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_3_LC_5_17_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_3_LC_5_17_3 .LUT_INIT=16'b0011101100001000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_3_LC_5_17_3  (
            .in0(N__92235),
            .in1(N__52463),
            .in2(N__40381),
            .in3(N__40105),
            .lcout(alt_command_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94337),
            .ce(),
            .sr(N__86454));
    defparam \Commands_frame_decoder.source_CH1data_0_LC_5_17_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_0_LC_5_17_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_0_LC_5_17_4 .LUT_INIT=16'b0010111100100000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_0_LC_5_17_4  (
            .in0(N__88263),
            .in1(N__40373),
            .in2(N__52465),
            .in3(N__40092),
            .lcout(alt_command_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94337),
            .ce(),
            .sr(N__86454));
    defparam \Commands_frame_decoder.source_CH1data_2_LC_5_17_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_2_LC_5_17_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_2_LC_5_17_5 .LUT_INIT=16'b0011101100001000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_2_LC_5_17_5  (
            .in0(N__92432),
            .in1(N__52462),
            .in2(N__40380),
            .in3(N__40362),
            .lcout(alt_command_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94337),
            .ce(),
            .sr(N__86454));
    defparam \Commands_frame_decoder.state_RNO_3_0_LC_5_17_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_3_0_LC_5_17_6 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_3_0_LC_5_17_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Commands_frame_decoder.state_RNO_3_0_LC_5_17_6  (
            .in0(N__88262),
            .in1(N__88642),
            .in2(N__92102),
            .in3(N__92430),
            .lcout(),
            .ltout(\Commands_frame_decoder.state_ns_i_a2_0_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNO_2_0_LC_5_17_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_2_0_LC_5_17_7 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_2_0_LC_5_17_7 .LUT_INIT=16'b1110110000000000;
    LogicCell40 \Commands_frame_decoder.state_RNO_2_0_LC_5_17_7  (
            .in0(N__41092),
            .in1(N__45960),
            .in2(N__40348),
            .in3(N__43159),
            .lcout(\Commands_frame_decoder.N_371 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH1data_esr_4_LC_5_18_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_esr_4_LC_5_18_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_esr_4_LC_5_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_esr_4_LC_5_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88828),
            .lcout(alt_command_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94352),
            .ce(N__45495),
            .sr(N__86450));
    defparam \Commands_frame_decoder.source_CH1data_esr_5_LC_5_18_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_esr_5_LC_5_18_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_esr_5_LC_5_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_esr_5_LC_5_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88666),
            .lcout(alt_command_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94352),
            .ce(N__45495),
            .sr(N__86450));
    defparam \Commands_frame_decoder.source_CH1data_esr_6_LC_5_18_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_esr_6_LC_5_18_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_esr_6_LC_5_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_esr_6_LC_5_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88470),
            .lcout(alt_command_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94352),
            .ce(N__45495),
            .sr(N__86450));
    defparam \Commands_frame_decoder.source_alt_kp_e_0_2_LC_5_19_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_2_LC_5_19_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_2_LC_5_19_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_e_0_2_LC_5_19_2  (
            .in0(_gnd_net_),
            .in1(N__92474),
            .in2(_gnd_net_),
            .in3(N__93149),
            .lcout(alt_kp_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94363),
            .ce(N__48691),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNILMDC_8_LC_5_19_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNILMDC_8_LC_5_19_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNILMDC_8_LC_5_19_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNILMDC_8_LC_5_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48442),
            .lcout(drone_altitude_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNISPHM_15_LC_5_20_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNISPHM_15_LC_5_20_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNISPHM_15_LC_5_20_0 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNISPHM_15_LC_5_20_0  (
            .in0(N__40296),
            .in1(N__40530),
            .in2(_gnd_net_),
            .in3(N__40563),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNISPHMZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_15_LC_5_20_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_15_LC_5_20_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_15_LC_5_20_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_15_LC_5_20_1  (
            .in0(N__40564),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94372),
            .ce(N__40495),
            .sr(N__86443));
    defparam \pid_alt.state_RNIAAPN5_1_LC_5_20_2 .C_ON=1'b0;
    defparam \pid_alt.state_RNIAAPN5_1_LC_5_20_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.state_RNIAAPN5_1_LC_5_20_2 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \pid_alt.state_RNIAAPN5_1_LC_5_20_2  (
            .in0(N__71026),
            .in1(N__69012),
            .in2(_gnd_net_),
            .in3(N__40444),
            .lcout(\pid_alt.un1_reset_1_0_i ),
            .ltout(\pid_alt.un1_reset_1_0_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.state_RNIVV066_1_LC_5_20_3 .C_ON=1'b0;
    defparam \pid_alt.state_RNIVV066_1_LC_5_20_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.state_RNIVV066_1_LC_5_20_3 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \pid_alt.state_RNIVV066_1_LC_5_20_3  (
            .in0(N__69013),
            .in1(_gnd_net_),
            .in2(N__40435),
            .in3(_gnd_net_),
            .lcout(\pid_alt.N_72_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_data_valid_2_sqmuxa_i_LC_5_20_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_data_valid_2_sqmuxa_i_LC_5_20_4 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_data_valid_2_sqmuxa_i_LC_5_20_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \dron_frame_decoder_1.source_data_valid_2_sqmuxa_i_LC_5_20_4  (
            .in0(N__71027),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48557),
            .lcout(\dron_frame_decoder_1.source_data_valid_2_sqmuxa_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNIB78K_2_LC_5_20_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNIB78K_2_LC_5_20_6 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNIB78K_2_LC_5_20_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \dron_frame_decoder_1.state_RNIB78K_2_LC_5_20_6  (
            .in0(_gnd_net_),
            .in1(N__46365),
            .in2(_gnd_net_),
            .in3(N__86588),
            .lcout(\dron_frame_decoder_1.N_708_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNI6P6K_4_LC_5_20_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNI6P6K_4_LC_5_20_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNI6P6K_4_LC_5_20_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \dron_frame_decoder_1.state_RNI6P6K_4_LC_5_20_7  (
            .in0(N__48556),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46339),
            .lcout(\dron_frame_decoder_1.state_RNI6P6KZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH1data_esr_7_LC_5_21_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_esr_7_LC_5_21_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_esr_7_LC_5_21_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_esr_7_LC_5_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__92103),
            .lcout(alt_command_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94381),
            .ce(N__45499),
            .sr(N__86441));
    defparam \ppm_encoder_1.init_pulses_RNI90081_3_LC_7_1_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI90081_3_LC_7_1_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI90081_3_LC_7_1_0 .LUT_INIT=16'b1111000001111000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI90081_3_LC_7_1_0  (
            .in0(N__53806),
            .in1(N__53691),
            .in2(N__44865),
            .in3(N__52878),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_fast_RNIJ2CB_0_LC_7_1_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_fast_RNIJ2CB_0_LC_7_1_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_fast_RNIJ2CB_0_LC_7_1_1 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \ppm_encoder_1.PPM_STATE_fast_RNIJ2CB_0_LC_7_1_1  (
            .in0(N__52879),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86584),
            .lcout(\ppm_encoder_1.N_295_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI7UV71_1_LC_7_1_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI7UV71_1_LC_7_1_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI7UV71_1_LC_7_1_2 .LUT_INIT=16'b1111000001111000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI7UV71_1_LC_7_1_2  (
            .in0(N__53805),
            .in1(N__53690),
            .in2(N__40420),
            .in3(N__52877),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone_sync.aux_0__0__0_LC_7_1_5 .C_ON=1'b0;
    defparam \uart_drone_sync.aux_0__0__0_LC_7_1_5 .SEQ_MODE=4'b1000;
    defparam \uart_drone_sync.aux_0__0__0_LC_7_1_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone_sync.aux_0__0__0_LC_7_1_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40579),
            .lcout(\uart_drone_sync.aux_0__0__0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94101),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5I0L2_3_LC_7_1_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5I0L2_3_LC_7_1_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5I0L2_3_LC_7_1_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5I0L2_3_LC_7_1_6  (
            .in0(N__44280),
            .in1(N__44343),
            .in2(_gnd_net_),
            .in3(N__47512),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5I0L2Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNICI741_5_LC_7_2_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNICI741_5_LC_7_2_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNICI741_5_LC_7_2_0 .LUT_INIT=16'b1011010011110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNICI741_5_LC_7_2_0  (
            .in0(N__52859),
            .in1(N__56305),
            .in2(N__49969),
            .in3(N__53793),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIA1081_4_LC_7_2_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIA1081_4_LC_7_2_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIA1081_4_LC_7_2_1 .LUT_INIT=16'b1010101001101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIA1081_4_LC_7_2_1  (
            .in0(N__50009),
            .in1(N__53696),
            .in2(N__53807),
            .in3(N__52860),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNITK131_0_14_LC_7_2_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNITK131_0_14_LC_7_2_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNITK131_0_14_LC_7_2_2 .LUT_INIT=16'b1011010011110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNITK131_0_14_LC_7_2_2  (
            .in0(N__52862),
            .in1(N__49648),
            .in2(N__48771),
            .in3(N__56308),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIOHJF3_13_LC_7_2_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIOHJF3_13_LC_7_2_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIOHJF3_13_LC_7_2_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIOHJF3_13_LC_7_2_3  (
            .in0(_gnd_net_),
            .in1(N__40573),
            .in2(_gnd_net_),
            .in3(N__44114),
            .lcout(\ppm_encoder_1.init_pulses_RNIOHJF3Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIEK741_7_LC_7_2_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIEK741_7_LC_7_2_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIEK741_7_LC_7_2_4 .LUT_INIT=16'b1011010011110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIEK741_7_LC_7_2_4  (
            .in0(N__52861),
            .in1(N__56306),
            .in2(N__49075),
            .in3(N__53794),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIUL131_0_15_LC_7_2_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIUL131_0_15_LC_7_2_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIUL131_0_15_LC_7_2_7 .LUT_INIT=16'b1100110001101100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIUL131_0_15_LC_7_2_7  (
            .in0(N__56307),
            .in1(N__48800),
            .in2(N__49676),
            .in3(N__52863),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI0O131_0_17_LC_7_3_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI0O131_0_17_LC_7_3_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI0O131_0_17_LC_7_3_0 .LUT_INIT=16'b1001110011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI0O131_0_17_LC_7_3_0  (
            .in0(N__52805),
            .in1(N__49172),
            .in2(N__56326),
            .in3(N__49644),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIPG131_10_LC_7_3_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIPG131_10_LC_7_3_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIPG131_10_LC_7_3_1 .LUT_INIT=16'b1111000001111000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIPG131_10_LC_7_3_1  (
            .in0(N__49641),
            .in1(N__56316),
            .in2(N__50118),
            .in3(N__52803),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIFL741_8_LC_7_3_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIFL741_8_LC_7_3_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIFL741_8_LC_7_3_2 .LUT_INIT=16'b1001110011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIFL741_8_LC_7_3_2  (
            .in0(N__52801),
            .in1(N__48961),
            .in2(N__56323),
            .in3(N__53789),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIF6081_9_LC_7_3_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIF6081_9_LC_7_3_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIF6081_9_LC_7_3_3 .LUT_INIT=16'b1111000001111000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIF6081_9_LC_7_3_3  (
            .in0(N__53787),
            .in1(N__53686),
            .in2(N__46520),
            .in3(N__52799),
            .lcout(\ppm_encoder_1.N_265_i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIH2561_9_LC_7_3_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIH2561_9_LC_7_3_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIH2561_9_LC_7_3_4 .LUT_INIT=16'b1001110011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIH2561_9_LC_7_3_4  (
            .in0(N__52802),
            .in1(N__46513),
            .in2(N__56324),
            .in3(N__49642),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIRI131_12_LC_7_3_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIRI131_12_LC_7_3_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIRI131_12_LC_7_3_6 .LUT_INIT=16'b1011111101000000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIRI131_12_LC_7_3_6  (
            .in0(N__52804),
            .in1(N__49643),
            .in2(N__56325),
            .in3(N__50850),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIR7411_13_LC_7_3_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIR7411_13_LC_7_3_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIR7411_13_LC_7_3_7 .LUT_INIT=16'b1111000001111000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIR7411_13_LC_7_3_7  (
            .in0(N__53788),
            .in1(N__56309),
            .in2(N__41873),
            .in3(N__52800),
            .lcout(\ppm_encoder_1.N_268_i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIGRJA2_13_LC_7_4_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIGRJA2_13_LC_7_4_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIGRJA2_13_LC_7_4_0 .LUT_INIT=16'b1110111011111110;
    LogicCell40 \ppm_encoder_1.elevator_RNIGRJA2_13_LC_7_4_0  (
            .in0(N__50739),
            .in1(N__40603),
            .in2(N__42379),
            .in3(N__47397),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_0_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIDDVF4_13_LC_7_4_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIDDVF4_13_LC_7_4_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIDDVF4_13_LC_7_4_1 .LUT_INIT=16'b0110011001101001;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIDDVF4_13_LC_7_4_1  (
            .in0(N__41858),
            .in1(N__41790),
            .in2(N__40606),
            .in3(N__44509),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_RNIO2KQ_13_LC_7_4_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_RNIO2KQ_13_LC_7_4_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.rudder_RNIO2KQ_13_LC_7_4_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ppm_encoder_1.rudder_RNIO2KQ_13_LC_7_4_4  (
            .in0(_gnd_net_),
            .in1(N__42298),
            .in2(_gnd_net_),
            .in3(N__53660),
            .lcout(\ppm_encoder_1.N_516 ),
            .ltout(\ppm_encoder_1.N_516_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_13_LC_7_4_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_13_LC_7_4_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_13_LC_7_4_5 .LUT_INIT=16'b1111110111111100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_13_LC_7_4_5  (
            .in0(N__47398),
            .in1(N__40597),
            .in2(N__40582),
            .in3(N__42378),
            .lcout(\ppm_encoder_1.pulses2count_9_0_1_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIFVUE1_11_LC_7_5_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIFVUE1_11_LC_7_5_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIFVUE1_11_LC_7_5_0 .LUT_INIT=16'b0101110100001100;
    LogicCell40 \ppm_encoder_1.throttle_RNIFVUE1_11_LC_7_5_0  (
            .in0(N__50174),
            .in1(N__44679),
            .in2(N__40651),
            .in3(N__44595),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_1_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_8_LC_7_5_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_8_LC_7_5_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_8_LC_7_5_1 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_8_LC_7_5_1  (
            .in0(N__54245),
            .in1(N__45061),
            .in2(_gnd_net_),
            .in3(N__54109),
            .lcout(\ppm_encoder_1.N_420 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIQ6411_12_LC_7_5_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIQ6411_12_LC_7_5_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIQ6411_12_LC_7_5_2 .LUT_INIT=16'b0000111110000111;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIQ6411_12_LC_7_5_2  (
            .in0(N__56274),
            .in1(N__53781),
            .in2(N__50848),
            .in3(N__52864),
            .lcout(\ppm_encoder_1.N_267_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_LC_7_5_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_LC_7_5_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_LC_7_5_3 .LUT_INIT=16'b0010001100000001;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_3_LC_7_5_3  (
            .in0(N__52866),
            .in1(N__71038),
            .in2(N__46907),
            .in3(N__49623),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94132),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_rep2_LC_7_5_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_rep2_LC_7_5_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_rep2_LC_7_5_5 .LUT_INIT=16'b0010001100000001;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_3_rep2_LC_7_5_5  (
            .in0(N__52867),
            .in1(N__71039),
            .in2(N__46908),
            .in3(N__53772),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94132),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIPMS41_12_LC_7_5_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIPMS41_12_LC_7_5_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIPMS41_12_LC_7_5_6 .LUT_INIT=16'b1111000001111000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIPMS41_12_LC_7_5_6  (
            .in0(N__53771),
            .in1(N__53656),
            .in2(N__50849),
            .in3(N__52865),
            .lcout(\ppm_encoder_1.N_267_i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone_sync.aux_1__0__0_LC_7_5_7 .C_ON=1'b0;
    defparam \uart_drone_sync.aux_1__0__0_LC_7_5_7 .SEQ_MODE=4'b1000;
    defparam \uart_drone_sync.aux_1__0__0_LC_7_5_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone_sync.aux_1__0__0_LC_7_5_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40663),
            .lcout(\uart_drone_sync.aux_1__0__0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94132),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_11_LC_7_6_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_11_LC_7_6_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_11_LC_7_6_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_11_LC_7_6_3  (
            .in0(_gnd_net_),
            .in1(N__50559),
            .in2(_gnd_net_),
            .in3(N__40649),
            .lcout(\ppm_encoder_1.N_431 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIDFS81_11_LC_7_6_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIDFS81_11_LC_7_6_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIDFS81_11_LC_7_6_4 .LUT_INIT=16'b0001111100010001;
    LogicCell40 \ppm_encoder_1.elevator_RNIDFS81_11_LC_7_6_4  (
            .in0(N__47410),
            .in1(N__40830),
            .in2(N__40775),
            .in3(N__53626),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_0_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNI6CI25_11_LC_7_6_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI6CI25_11_LC_7_6_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI6CI25_11_LC_7_6_5 .LUT_INIT=16'b0011001100110110;
    LogicCell40 \ppm_encoder_1.elevator_RNI6CI25_11_LC_7_6_5  (
            .in0(N__40615),
            .in1(N__42277),
            .in2(N__40609),
            .in3(N__44514),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_11_LC_7_6_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_11_LC_7_6_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_11_LC_7_6_6 .LUT_INIT=16'b1111010001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_11_LC_7_6_6  (
            .in0(N__47411),
            .in1(N__40831),
            .in2(N__40776),
            .in3(N__47516),
            .lcout(\ppm_encoder_1.pulses2count_9_0_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_esr_RNIQU9H1_4_LC_7_6_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_RNIQU9H1_4_LC_7_6_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.rudder_esr_RNIQU9H1_4_LC_7_6_7 .LUT_INIT=16'b1010000011101100;
    LogicCell40 \ppm_encoder_1.rudder_esr_RNIQU9H1_4_LC_7_6_7  (
            .in0(N__53625),
            .in1(N__46705),
            .in2(N__47029),
            .in3(N__47409),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNISKME2_10_LC_7_7_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNISKME2_10_LC_7_7_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNISKME2_10_LC_7_7_0 .LUT_INIT=16'b1111101011111110;
    LogicCell40 \ppm_encoder_1.elevator_RNISKME2_10_LC_7_7_0  (
            .in0(N__40708),
            .in1(N__42419),
            .in2(N__44518),
            .in3(N__47432),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_2_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIHP6T4_10_LC_7_7_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIHP6T4_10_LC_7_7_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIHP6T4_10_LC_7_7_1 .LUT_INIT=16'b0110011001101001;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIHP6T4_10_LC_7_7_1  (
            .in0(N__41794),
            .in1(N__50110),
            .in2(N__40714),
            .in3(N__40702),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_0_axb_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI8E326_10_LC_7_7_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI8E326_10_LC_7_7_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI8E326_10_LC_7_7_2 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI8E326_10_LC_7_7_2  (
            .in0(_gnd_net_),
            .in1(N__43803),
            .in2(N__40711),
            .in3(_gnd_net_),
            .lcout(\ppm_encoder_1.init_pulses_RNI8E326Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_RNIKVJQ_10_LC_7_7_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_RNIKVJQ_10_LC_7_7_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.rudder_RNIKVJQ_10_LC_7_7_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ppm_encoder_1.rudder_RNIKVJQ_10_LC_7_7_3  (
            .in0(_gnd_net_),
            .in1(N__47085),
            .in2(_gnd_net_),
            .in3(N__42198),
            .lcout(\ppm_encoder_1.N_458 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIDTUE1_10_LC_7_7_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIDTUE1_10_LC_7_7_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIDTUE1_10_LC_7_7_4 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \ppm_encoder_1.throttle_RNIDTUE1_10_LC_7_7_4  (
            .in0(N__44682),
            .in1(N__42224),
            .in2(N__46479),
            .in3(N__44607),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_1_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_10_LC_7_7_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_10_LC_7_7_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_10_LC_7_7_6 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.aileron_10_LC_7_7_6  (
            .in0(N__53458),
            .in1(N__47758),
            .in2(N__42234),
            .in3(N__51320),
            .lcout(\ppm_encoder_1.aileronZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94151),
            .ce(),
            .sr(N__86503));
    defparam \ppm_encoder_1.elevator_1_LC_7_8_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_1_LC_7_8_0 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_1_LC_7_8_0 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \ppm_encoder_1.elevator_1_LC_7_8_0  (
            .in0(N__47290),
            .in1(N__55000),
            .in2(N__51371),
            .in3(N__40685),
            .lcout(\ppm_encoder_1.elevatorZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94162),
            .ce(),
            .sr(N__86497));
    defparam \ppm_encoder_1.elevator_11_LC_7_8_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_11_LC_7_8_2 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_11_LC_7_8_2 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.elevator_11_LC_7_8_2  (
            .in0(N__54646),
            .in1(N__47614),
            .in2(N__51370),
            .in3(N__40829),
            .lcout(\ppm_encoder_1.elevatorZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94162),
            .ce(),
            .sr(N__86497));
    defparam \ppm_encoder_1.elevator_2_LC_7_8_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_2_LC_7_8_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_2_LC_7_8_3 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.elevator_2_LC_7_8_3  (
            .in0(N__60226),
            .in1(N__47275),
            .in2(N__40808),
            .in3(N__51344),
            .lcout(\ppm_encoder_1.elevatorZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94162),
            .ce(),
            .sr(N__86497));
    defparam \ppm_encoder_1.rudder_7_LC_7_8_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_7_LC_7_8_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_7_LC_7_8_4 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.rudder_7_LC_7_8_4  (
            .in0(N__40747),
            .in1(N__40855),
            .in2(N__51372),
            .in3(N__44163),
            .lcout(\ppm_encoder_1.rudderZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94162),
            .ce(),
            .sr(N__86497));
    defparam \ppm_encoder_1.rudder_11_LC_7_8_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_11_LC_7_8_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.rudder_11_LC_7_8_5 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.rudder_11_LC_7_8_5  (
            .in0(N__40876),
            .in1(N__40920),
            .in2(N__40777),
            .in3(N__51345),
            .lcout(\ppm_encoder_1.rudderZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94162),
            .ce(),
            .sr(N__86497));
    defparam \ppm_encoder_1.rudder_9_LC_7_8_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_9_LC_7_8_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_9_LC_7_8_6 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.rudder_9_LC_7_8_6  (
            .in0(N__40942),
            .in1(N__40735),
            .in2(N__51373),
            .in3(N__46955),
            .lcout(\ppm_encoder_1.rudderZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94162),
            .ce(),
            .sr(N__86497));
    defparam \ppm_encoder_1.un1_rudder_cry_6_c_LC_7_9_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_6_c_LC_7_9_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_6_c_LC_7_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_6_c_LC_7_9_0  (
            .in0(_gnd_net_),
            .in1(N__43764),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_9_0_),
            .carryout(\ppm_encoder_1.un1_rudder_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_6_THRU_LUT4_0_LC_7_9_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_6_THRU_LUT4_0_LC_7_9_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_6_THRU_LUT4_0_LC_7_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_6_THRU_LUT4_0_LC_7_9_1  (
            .in0(_gnd_net_),
            .in1(N__40854),
            .in2(_gnd_net_),
            .in3(N__40741),
            .lcout(\ppm_encoder_1.un1_rudder_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_6 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_7_THRU_LUT4_0_LC_7_9_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_7_THRU_LUT4_0_LC_7_9_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_7_THRU_LUT4_0_LC_7_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_7_THRU_LUT4_0_LC_7_9_2  (
            .in0(_gnd_net_),
            .in1(N__42396),
            .in2(_gnd_net_),
            .in3(N__40738),
            .lcout(\ppm_encoder_1.un1_rudder_cry_7_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_7 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_8_THRU_LUT4_0_LC_7_9_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_8_THRU_LUT4_0_LC_7_9_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_8_THRU_LUT4_0_LC_7_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_8_THRU_LUT4_0_LC_7_9_3  (
            .in0(_gnd_net_),
            .in1(N__40941),
            .in2(_gnd_net_),
            .in3(N__40729),
            .lcout(\ppm_encoder_1.un1_rudder_cry_8_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_8 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_9_THRU_LUT4_0_LC_7_9_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_9_THRU_LUT4_0_LC_7_9_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_9_THRU_LUT4_0_LC_7_9_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_9_THRU_LUT4_0_LC_7_9_4  (
            .in0(_gnd_net_),
            .in1(N__42339),
            .in2(_gnd_net_),
            .in3(N__40726),
            .lcout(\ppm_encoder_1.un1_rudder_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_9 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_10_THRU_LUT4_0_LC_7_9_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_10_THRU_LUT4_0_LC_7_9_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_10_THRU_LUT4_0_LC_7_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_10_THRU_LUT4_0_LC_7_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__40921),
            .in3(N__40870),
            .lcout(\ppm_encoder_1.un1_rudder_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_10 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_11_THRU_LUT4_0_LC_7_9_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_11_THRU_LUT4_0_LC_7_9_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_11_THRU_LUT4_0_LC_7_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_11_THRU_LUT4_0_LC_7_9_6  (
            .in0(_gnd_net_),
            .in1(N__42474),
            .in2(_gnd_net_),
            .in3(N__40867),
            .lcout(\ppm_encoder_1.un1_rudder_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_11 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_12_THRU_LUT4_0_LC_7_9_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_12_THRU_LUT4_0_LC_7_9_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_12_THRU_LUT4_0_LC_7_9_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_12_THRU_LUT4_0_LC_7_9_7  (
            .in0(_gnd_net_),
            .in1(N__42315),
            .in2(N__65788),
            .in3(N__40864),
            .lcout(\ppm_encoder_1.un1_rudder_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_12 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_esr_14_LC_7_10_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_14_LC_7_10_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_esr_14_LC_7_10_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.rudder_esr_14_LC_7_10_0  (
            .in0(_gnd_net_),
            .in1(N__40888),
            .in2(_gnd_net_),
            .in3(N__40861),
            .lcout(\ppm_encoder_1.rudderZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94190),
            .ce(N__47985),
            .sr(N__86486));
    defparam \scaler_4.un2_source_data_0_cry_1_c_LC_7_11_0 .C_ON=1'b1;
    defparam \scaler_4.un2_source_data_0_cry_1_c_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un2_source_data_0_cry_1_c_LC_7_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \scaler_4.un2_source_data_0_cry_1_c_LC_7_11_0  (
            .in0(_gnd_net_),
            .in1(N__45259),
            .in2(N__45214),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_11_0_),
            .carryout(\scaler_4.un2_source_data_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.source_data_1_esr_6_LC_7_11_1 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_6_LC_7_11_1 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_6_LC_7_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_6_LC_7_11_1  (
            .in0(_gnd_net_),
            .in1(N__42600),
            .in2(N__45267),
            .in3(N__40858),
            .lcout(scaler_4_data_6),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_1 ),
            .carryout(\scaler_4.un2_source_data_0_cry_2 ),
            .clk(N__94205),
            .ce(N__48067),
            .sr(N__86479));
    defparam \scaler_4.source_data_1_esr_7_LC_7_11_2 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_7_LC_7_11_2 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_7_LC_7_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_7_LC_7_11_2  (
            .in0(_gnd_net_),
            .in1(N__42579),
            .in2(N__42604),
            .in3(N__40837),
            .lcout(scaler_4_data_7),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_2 ),
            .carryout(\scaler_4.un2_source_data_0_cry_3 ),
            .clk(N__94205),
            .ce(N__48067),
            .sr(N__86479));
    defparam \scaler_4.source_data_1_esr_8_LC_7_11_3 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_8_LC_7_11_3 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_8_LC_7_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_8_LC_7_11_3  (
            .in0(_gnd_net_),
            .in1(N__42558),
            .in2(N__42583),
            .in3(N__40834),
            .lcout(scaler_4_data_8),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_3 ),
            .carryout(\scaler_4.un2_source_data_0_cry_4 ),
            .clk(N__94205),
            .ce(N__48067),
            .sr(N__86479));
    defparam \scaler_4.source_data_1_esr_9_LC_7_11_4 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_9_LC_7_11_4 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_9_LC_7_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_9_LC_7_11_4  (
            .in0(_gnd_net_),
            .in1(N__42537),
            .in2(N__42562),
            .in3(N__40927),
            .lcout(scaler_4_data_9),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_4 ),
            .carryout(\scaler_4.un2_source_data_0_cry_5 ),
            .clk(N__94205),
            .ce(N__48067),
            .sr(N__86479));
    defparam \scaler_4.source_data_1_esr_10_LC_7_11_5 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_10_LC_7_11_5 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_10_LC_7_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_10_LC_7_11_5  (
            .in0(_gnd_net_),
            .in1(N__42516),
            .in2(N__42541),
            .in3(N__40924),
            .lcout(scaler_4_data_10),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_5 ),
            .carryout(\scaler_4.un2_source_data_0_cry_6 ),
            .clk(N__94205),
            .ce(N__48067),
            .sr(N__86479));
    defparam \scaler_4.source_data_1_esr_11_LC_7_11_6 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_11_LC_7_11_6 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_11_LC_7_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_11_LC_7_11_6  (
            .in0(_gnd_net_),
            .in1(N__42501),
            .in2(N__42520),
            .in3(N__40900),
            .lcout(scaler_4_data_11),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_6 ),
            .carryout(\scaler_4.un2_source_data_0_cry_7 ),
            .clk(N__94205),
            .ce(N__48067),
            .sr(N__86479));
    defparam \scaler_4.source_data_1_esr_12_LC_7_11_7 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_12_LC_7_11_7 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_12_LC_7_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_12_LC_7_11_7  (
            .in0(_gnd_net_),
            .in1(N__42489),
            .in2(N__42505),
            .in3(N__40897),
            .lcout(scaler_4_data_12),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_7 ),
            .carryout(\scaler_4.un2_source_data_0_cry_8 ),
            .clk(N__94205),
            .ce(N__48067),
            .sr(N__86479));
    defparam \scaler_4.source_data_1_esr_13_LC_7_12_0 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_13_LC_7_12_0 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_13_LC_7_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_13_LC_7_12_0  (
            .in0(_gnd_net_),
            .in1(N__42490),
            .in2(N__42748),
            .in3(N__40894),
            .lcout(scaler_4_data_13),
            .ltout(),
            .carryin(bfn_7_12_0_),
            .carryout(\scaler_4.un2_source_data_0_cry_9 ),
            .clk(N__94221),
            .ce(N__48063),
            .sr(N__86470));
    defparam \scaler_4.source_data_1_esr_14_LC_7_12_1 .C_ON=1'b0;
    defparam \scaler_4.source_data_1_esr_14_LC_7_12_1 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_14_LC_7_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \scaler_4.source_data_1_esr_14_LC_7_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40891),
            .lcout(scaler_4_data_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94221),
            .ce(N__48063),
            .sr(N__86470));
    defparam \Commands_frame_decoder.preinit_RNIHOV81_LC_7_13_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.preinit_RNIHOV81_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.preinit_RNIHOV81_LC_7_13_0 .LUT_INIT=16'b0000000001011111;
    LogicCell40 \Commands_frame_decoder.preinit_RNIHOV81_LC_7_13_0  (
            .in0(N__48286),
            .in1(_gnd_net_),
            .in2(N__48327),
            .in3(N__40976),
            .lcout(),
            .ltout(\Commands_frame_decoder.preinit_RNIHOVZ0Z81_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNIATE75_13_LC_7_13_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNIATE75_13_LC_7_13_1 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNIATE75_13_LC_7_13_1 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \Commands_frame_decoder.WDT_RNIATE75_13_LC_7_13_1  (
            .in0(N__42771),
            .in1(N__48321),
            .in2(N__40879),
            .in3(N__40984),
            .lcout(\Commands_frame_decoder.state_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNIET8A1_0_4_LC_7_13_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNIET8A1_0_4_LC_7_13_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNIET8A1_0_4_LC_7_13_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Commands_frame_decoder.WDT_RNIET8A1_0_4_LC_7_13_3  (
            .in0(N__42929),
            .in1(N__42635),
            .in2(N__42909),
            .in3(N__42656),
            .lcout(\Commands_frame_decoder.WDT_RNIET8A1_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNIHV6P_11_LC_7_13_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNIHV6P_11_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNIHV6P_11_LC_7_13_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Commands_frame_decoder.WDT_RNIHV6P_11_LC_7_13_4  (
            .in0(_gnd_net_),
            .in1(N__42793),
            .in2(_gnd_net_),
            .in3(N__42820),
            .lcout(),
            .ltout(\Commands_frame_decoder.WDT_RNIHV6PZ0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNI30853_10_LC_7_13_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNI30853_10_LC_7_13_5 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNI30853_10_LC_7_13_5 .LUT_INIT=16'b0010111110101111;
    LogicCell40 \Commands_frame_decoder.WDT_RNI30853_10_LC_7_13_5  (
            .in0(N__42843),
            .in1(N__41041),
            .in2(N__40993),
            .in3(N__40990),
            .lcout(\Commands_frame_decoder.WDT_RNI30853Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.preinit_LC_7_13_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.preinit_LC_7_13_6 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.preinit_LC_7_13_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Commands_frame_decoder.preinit_LC_7_13_6  (
            .in0(N__55281),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40977),
            .lcout(\Commands_frame_decoder.preinitZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94238),
            .ce(),
            .sr(N__86465));
    defparam \Commands_frame_decoder.source_data_valid_LC_7_13_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_data_valid_LC_7_13_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_data_valid_LC_7_13_7 .LUT_INIT=16'b1110111011100010;
    LogicCell40 \Commands_frame_decoder.source_data_valid_LC_7_13_7  (
            .in0(N__40978),
            .in1(N__55282),
            .in2(N__48103),
            .in3(N__41128),
            .lcout(debug_CH3_20A_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94238),
            .ce(),
            .sr(N__86465));
    defparam \Commands_frame_decoder.WDT_RNIHV6P_0_11_LC_7_14_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNIHV6P_0_11_LC_7_14_0 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNIHV6P_0_11_LC_7_14_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Commands_frame_decoder.WDT_RNIHV6P_0_11_LC_7_14_0  (
            .in0(_gnd_net_),
            .in1(N__42794),
            .in2(_gnd_net_),
            .in3(N__42821),
            .lcout(\Commands_frame_decoder.WDT_RNIHV6P_0Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNI2VDI1_10_LC_7_14_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNI2VDI1_10_LC_7_14_1 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNI2VDI1_10_LC_7_14_1 .LUT_INIT=16'b0011001100110111;
    LogicCell40 \Commands_frame_decoder.WDT_RNI2VDI1_10_LC_7_14_1  (
            .in0(N__42822),
            .in1(N__42770),
            .in2(N__42799),
            .in3(N__42842),
            .lcout(\Commands_frame_decoder.WDT_RNI2VDI1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNITK4L_0_8_LC_7_14_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNITK4L_0_8_LC_7_14_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNITK4L_0_8_LC_7_14_2 .LUT_INIT=16'b0000010100000101;
    LogicCell40 \Commands_frame_decoder.WDT_RNITK4L_0_8_LC_7_14_2  (
            .in0(N__42882),
            .in1(_gnd_net_),
            .in2(N__42865),
            .in3(_gnd_net_),
            .lcout(\Commands_frame_decoder.WDT_RNITK4L_0Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNIET8A1_4_LC_7_14_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNIET8A1_4_LC_7_14_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNIET8A1_4_LC_7_14_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Commands_frame_decoder.WDT_RNIET8A1_4_LC_7_14_3  (
            .in0(N__42930),
            .in1(N__42636),
            .in2(N__42910),
            .in3(N__42657),
            .lcout(),
            .ltout(\Commands_frame_decoder.WDT_RNIET8A1Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNIUG2B4_4_LC_7_14_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNIUG2B4_4_LC_7_14_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNIUG2B4_4_LC_7_14_4 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \Commands_frame_decoder.WDT_RNIUG2B4_4_LC_7_14_4  (
            .in0(N__40966),
            .in1(N__40960),
            .in2(N__40954),
            .in3(N__40951),
            .lcout(\Commands_frame_decoder.WDT8lt14_0 ),
            .ltout(\Commands_frame_decoder.WDT8lt14_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNIPRJG5_14_LC_7_14_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNIPRJG5_14_LC_7_14_5 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNIPRJG5_14_LC_7_14_5 .LUT_INIT=16'b0100010001000000;
    LogicCell40 \Commands_frame_decoder.WDT_RNIPRJG5_14_LC_7_14_5  (
            .in0(N__55267),
            .in1(N__48325),
            .in2(N__40945),
            .in3(N__48287),
            .lcout(\Commands_frame_decoder.N_365_0 ),
            .ltout(\Commands_frame_decoder.N_365_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNO_0_0_LC_7_14_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_0_0_LC_7_14_6 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_0_0_LC_7_14_6 .LUT_INIT=16'b0000001000001010;
    LogicCell40 \Commands_frame_decoder.state_RNO_0_0_LC_7_14_6  (
            .in0(N__41226),
            .in1(N__55268),
            .in2(N__41044),
            .in3(N__41629),
            .lcout(\Commands_frame_decoder.N_372 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNITK4L_8_LC_7_14_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNITK4L_8_LC_7_14_7 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNITK4L_8_LC_7_14_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Commands_frame_decoder.WDT_RNITK4L_8_LC_7_14_7  (
            .in0(_gnd_net_),
            .in1(N__42860),
            .in2(_gnd_net_),
            .in3(N__42881),
            .lcout(\Commands_frame_decoder.WDT_RNITK4LZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_9_LC_7_15_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_9_LC_7_15_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_9_LC_7_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_9_LC_7_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41035),
            .lcout(\pid_front.error_p_regZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94274),
            .ce(N__93315),
            .sr(N__92975));
    defparam \uart_pc.state_RNO_0_2_LC_7_16_0 .C_ON=1'b0;
    defparam \uart_pc.state_RNO_0_2_LC_7_16_0 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNO_0_2_LC_7_16_0 .LUT_INIT=16'b0000000000111010;
    LogicCell40 \uart_pc.state_RNO_0_2_LC_7_16_0  (
            .in0(N__41117),
            .in1(N__52229),
            .in2(N__41020),
            .in3(N__70961),
            .lcout(),
            .ltout(\uart_pc.state_srsts_i_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_2_LC_7_16_1 .C_ON=1'b0;
    defparam \uart_pc.state_2_LC_7_16_1 .SEQ_MODE=4'b1000;
    defparam \uart_pc.state_2_LC_7_16_1 .LUT_INIT=16'b1101000011110000;
    LogicCell40 \uart_pc.state_2_LC_7_16_1  (
            .in0(N__41349),
            .in1(N__41018),
            .in2(N__40999),
            .in3(N__41400),
            .lcout(\uart_pc.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94290),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIGRIF1_2_LC_7_16_2 .C_ON=1'b0;
    defparam \uart_pc.state_RNIGRIF1_2_LC_7_16_2 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIGRIF1_2_LC_7_16_2 .LUT_INIT=16'b0101010011111100;
    LogicCell40 \uart_pc.state_RNIGRIF1_2_LC_7_16_2  (
            .in0(N__41398),
            .in1(N__41116),
            .in2(N__45794),
            .in3(N__41348),
            .lcout(\uart_pc.timer_Count_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNI5UFA2_3_LC_7_16_3 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNI5UFA2_3_LC_7_16_3 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNI5UFA2_3_LC_7_16_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uart_pc.timer_Count_RNI5UFA2_3_LC_7_16_3  (
            .in0(N__41347),
            .in1(N__45536),
            .in2(_gnd_net_),
            .in3(N__41397),
            .lcout(\uart_pc.N_144_1 ),
            .ltout(\uart_pc.N_144_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_3_LC_7_16_4 .C_ON=1'b0;
    defparam \uart_pc.state_3_LC_7_16_4 .SEQ_MODE=4'b1000;
    defparam \uart_pc.state_3_LC_7_16_4 .LUT_INIT=16'b0000000000100011;
    LogicCell40 \uart_pc.state_3_LC_7_16_4  (
            .in0(N__41118),
            .in1(N__41098),
            .in2(N__40996),
            .in3(N__70962),
            .lcout(\uart_pc.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94290),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIITIF1_4_LC_7_16_5 .C_ON=1'b0;
    defparam \uart_pc.state_RNIITIF1_4_LC_7_16_5 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIITIF1_4_LC_7_16_5 .LUT_INIT=16'b0101000100010001;
    LogicCell40 \uart_pc.state_RNIITIF1_4_LC_7_16_5  (
            .in0(N__45843),
            .in1(N__45780),
            .in2(N__41350),
            .in3(N__41396),
            .lcout(\uart_pc.un1_state_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_data_valid_RNO_0_LC_7_16_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_data_valid_RNO_0_LC_7_16_6 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.source_data_valid_RNO_0_LC_7_16_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.source_data_valid_RNO_0_LC_7_16_6  (
            .in0(_gnd_net_),
            .in1(N__41623),
            .in2(_gnd_net_),
            .in3(N__41219),
            .lcout(\Commands_frame_decoder.count_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNO_0_3_LC_7_16_7 .C_ON=1'b0;
    defparam \uart_pc.state_RNO_0_3_LC_7_16_7 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNO_0_3_LC_7_16_7 .LUT_INIT=16'b0001001100110011;
    LogicCell40 \uart_pc.state_RNO_0_3_LC_7_16_7  (
            .in0(N__41346),
            .in1(N__45781),
            .in2(N__41119),
            .in3(N__41399),
            .lcout(\uart_pc.N_145 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_1_LC_7_17_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_1_LC_7_17_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_1_LC_7_17_0 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \Commands_frame_decoder.state_1_LC_7_17_0  (
            .in0(N__45980),
            .in1(N__69408),
            .in2(N__41533),
            .in3(N__43157),
            .lcout(\Commands_frame_decoder.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94305),
            .ce(),
            .sr(N__86447));
    defparam \Commands_frame_decoder.state_RNI6QPK_1_LC_7_17_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNI6QPK_1_LC_7_17_1 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNI6QPK_1_LC_7_17_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Commands_frame_decoder.state_RNI6QPK_1_LC_7_17_1  (
            .in0(_gnd_net_),
            .in1(N__41217),
            .in2(_gnd_net_),
            .in3(N__45979),
            .lcout(\Commands_frame_decoder.N_370_2 ),
            .ltout(\Commands_frame_decoder.N_370_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNO_1_0_LC_7_17_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_1_0_LC_7_17_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_1_0_LC_7_17_2 .LUT_INIT=16'b0011001100100011;
    LogicCell40 \Commands_frame_decoder.state_RNO_1_0_LC_7_17_2  (
            .in0(N__41547),
            .in1(N__41083),
            .in2(N__41074),
            .in3(N__41055),
            .lcout(),
            .ltout(\Commands_frame_decoder.state_ns_i_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_0_LC_7_17_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_0_LC_7_17_3 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.state_0_LC_7_17_3 .LUT_INIT=16'b0000000001110000;
    LogicCell40 \Commands_frame_decoder.state_0_LC_7_17_3  (
            .in0(N__45984),
            .in1(N__69410),
            .in2(N__41071),
            .in3(N__41068),
            .lcout(\Commands_frame_decoder.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94305),
            .ce(),
            .sr(N__86447));
    defparam \Commands_frame_decoder.state_2_LC_7_17_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_2_LC_7_17_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_2_LC_7_17_4 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \Commands_frame_decoder.state_2_LC_7_17_4  (
            .in0(N__69409),
            .in1(N__45961),
            .in2(N__41197),
            .in3(N__43158),
            .lcout(\Commands_frame_decoder.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94305),
            .ce(),
            .sr(N__86447));
    defparam \Commands_frame_decoder.state_RNO_0_14_LC_7_17_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_0_14_LC_7_17_5 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_0_14_LC_7_17_5 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \Commands_frame_decoder.state_RNO_0_14_LC_7_17_5  (
            .in0(N__41627),
            .in1(N__55206),
            .in2(_gnd_net_),
            .in3(N__41218),
            .lcout(),
            .ltout(\Commands_frame_decoder.state_RNO_0Z0Z_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_14_LC_7_17_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_14_LC_7_17_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_14_LC_7_17_6 .LUT_INIT=16'b1000100011111000;
    LogicCell40 \Commands_frame_decoder.state_14_LC_7_17_6  (
            .in0(N__55207),
            .in1(N__48625),
            .in2(N__41059),
            .in3(N__41056),
            .lcout(\Commands_frame_decoder.stateZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94305),
            .ce(),
            .sr(N__86447));
    defparam \Commands_frame_decoder.state_RNIEI1J_2_LC_7_17_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIEI1J_2_LC_7_17_7 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIEI1J_2_LC_7_17_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_RNIEI1J_2_LC_7_17_7  (
            .in0(_gnd_net_),
            .in1(N__41193),
            .in2(_gnd_net_),
            .in3(N__55205),
            .lcout(\Commands_frame_decoder.un1_sink_data_valid_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNIPD2K1_2_LC_7_18_0 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNIPD2K1_2_LC_7_18_0 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNIPD2K1_2_LC_7_18_0 .LUT_INIT=16'b1100110010000000;
    LogicCell40 \uart_pc.timer_Count_RNIPD2K1_2_LC_7_18_0  (
            .in0(N__41330),
            .in1(N__45840),
            .in2(N__41157),
            .in3(N__41390),
            .lcout(\uart_pc.data_rdyc_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIFJ1J_3_LC_7_18_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIFJ1J_3_LC_7_18_1 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIFJ1J_3_LC_7_18_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_RNIFJ1J_3_LC_7_18_1  (
            .in0(_gnd_net_),
            .in1(N__52423),
            .in2(_gnd_net_),
            .in3(N__55263),
            .lcout(\Commands_frame_decoder.source_CH2data_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNO_0_0_LC_7_18_3 .C_ON=1'b0;
    defparam \uart_pc.state_RNO_0_0_LC_7_18_3 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNO_0_0_LC_7_18_3 .LUT_INIT=16'b0101010100010001;
    LogicCell40 \uart_pc.state_RNO_0_0_LC_7_18_3  (
            .in0(N__70978),
            .in1(N__41172),
            .in2(_gnd_net_),
            .in3(N__52241),
            .lcout(),
            .ltout(\uart_pc.state_srsts_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_0_LC_7_18_4 .C_ON=1'b0;
    defparam \uart_pc.state_0_LC_7_18_4 .SEQ_MODE=4'b1000;
    defparam \uart_pc.state_0_LC_7_18_4 .LUT_INIT=16'b1100111110001111;
    LogicCell40 \uart_pc.state_0_LC_7_18_4  (
            .in0(N__45870),
            .in1(N__45841),
            .in2(N__41185),
            .in3(N__41391),
            .lcout(\uart_pc.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94323),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_2_LC_7_18_5 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_2_LC_7_18_5 .SEQ_MODE=4'b1000;
    defparam \uart_pc.timer_Count_2_LC_7_18_5 .LUT_INIT=16'b0100010001000000;
    LogicCell40 \uart_pc.timer_Count_2_LC_7_18_5  (
            .in0(N__70979),
            .in1(N__41137),
            .in2(N__41283),
            .in3(N__41579),
            .lcout(\uart_pc.timer_CountZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94323),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNIVT8S_2_LC_7_18_6 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNIVT8S_2_LC_7_18_6 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNIVT8S_2_LC_7_18_6 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \uart_pc.timer_Count_RNIVT8S_2_LC_7_18_6  (
            .in0(N__41331),
            .in1(_gnd_net_),
            .in2(N__41158),
            .in3(_gnd_net_),
            .lcout(\uart_pc.N_126_li ),
            .ltout(\uart_pc.N_126_li_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIMQ8T1_4_LC_7_18_7 .C_ON=1'b0;
    defparam \uart_pc.state_RNIMQ8T1_4_LC_7_18_7 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIMQ8T1_4_LC_7_18_7 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \uart_pc.state_RNIMQ8T1_4_LC_7_18_7  (
            .in0(N__70977),
            .in1(N__41401),
            .in2(N__41161),
            .in3(N__45842),
            .lcout(\uart_pc.N_143 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNIRP8S_1_LC_7_19_0 .C_ON=1'b1;
    defparam \uart_pc.timer_Count_RNIRP8S_1_LC_7_19_0 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNIRP8S_1_LC_7_19_0 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \uart_pc.timer_Count_RNIRP8S_1_LC_7_19_0  (
            .in0(N__41305),
            .in1(N__41238),
            .in2(N__41308),
            .in3(_gnd_net_),
            .lcout(\uart_pc.un1_state_2_0_a3_0 ),
            .ltout(),
            .carryin(bfn_7_19_0_),
            .carryout(\uart_pc.un4_timer_Count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNO_0_2_LC_7_19_1 .C_ON=1'b1;
    defparam \uart_pc.timer_Count_RNO_0_2_LC_7_19_1 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNO_0_2_LC_7_19_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_pc.timer_Count_RNO_0_2_LC_7_19_1  (
            .in0(_gnd_net_),
            .in1(N__41156),
            .in2(_gnd_net_),
            .in3(N__41131),
            .lcout(\uart_pc.timer_Count_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\uart_pc.un4_timer_Count_1_cry_1 ),
            .carryout(\uart_pc.un4_timer_Count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNO_0_3_LC_7_19_2 .C_ON=1'b1;
    defparam \uart_pc.timer_Count_RNO_0_3_LC_7_19_2 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNO_0_3_LC_7_19_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_pc.timer_Count_RNO_0_3_LC_7_19_2  (
            .in0(_gnd_net_),
            .in1(N__41329),
            .in2(_gnd_net_),
            .in3(N__41413),
            .lcout(\uart_pc.timer_Count_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\uart_pc.un4_timer_Count_1_cry_2 ),
            .carryout(\uart_pc.un4_timer_Count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNO_0_4_LC_7_19_3 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNO_0_4_LC_7_19_3 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNO_0_4_LC_7_19_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uart_pc.timer_Count_RNO_0_4_LC_7_19_3  (
            .in0(_gnd_net_),
            .in1(N__41395),
            .in2(_gnd_net_),
            .in3(N__41410),
            .lcout(\uart_pc.timer_Count_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_0_LC_7_19_5 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_0_LC_7_19_5 .SEQ_MODE=4'b1000;
    defparam \uart_pc.timer_Count_0_LC_7_19_5 .LUT_INIT=16'b0000000001010100;
    LogicCell40 \uart_pc.timer_Count_0_LC_7_19_5  (
            .in0(N__70982),
            .in1(N__41571),
            .in2(N__41284),
            .in3(N__41306),
            .lcout(\uart_pc.timer_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94338),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_4_LC_7_19_6 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_4_LC_7_19_6 .SEQ_MODE=4'b1000;
    defparam \uart_pc.timer_Count_4_LC_7_19_6 .LUT_INIT=16'b0000000011001000;
    LogicCell40 \uart_pc.timer_Count_4_LC_7_19_6  (
            .in0(N__41573),
            .in1(N__41407),
            .in2(N__41286),
            .in3(N__70984),
            .lcout(\uart_pc.timer_CountZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94338),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_3_LC_7_19_7 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_3_LC_7_19_7 .SEQ_MODE=4'b1000;
    defparam \uart_pc.timer_Count_3_LC_7_19_7 .LUT_INIT=16'b0100010001000000;
    LogicCell40 \uart_pc.timer_Count_3_LC_7_19_7  (
            .in0(N__70983),
            .in1(N__41356),
            .in2(N__41285),
            .in3(N__41572),
            .lcout(\uart_pc.timer_CountZ1Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94338),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNO_0_1_LC_7_20_1 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNO_0_1_LC_7_20_1 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNO_0_1_LC_7_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_pc.timer_Count_RNO_0_1_LC_7_20_1  (
            .in0(_gnd_net_),
            .in1(N__41307),
            .in2(_gnd_net_),
            .in3(N__41239),
            .lcout(),
            .ltout(\uart_pc.timer_Count_RNO_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_1_LC_7_20_2 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_1_LC_7_20_2 .SEQ_MODE=4'b1000;
    defparam \uart_pc.timer_Count_1_LC_7_20_2 .LUT_INIT=16'b0101000001000000;
    LogicCell40 \uart_pc.timer_Count_1_LC_7_20_2  (
            .in0(N__71023),
            .in1(N__41287),
            .in2(N__41242),
            .in3(N__41583),
            .lcout(\uart_pc.timer_CountZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94353),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNI4N6K_2_LC_7_20_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNI4N6K_2_LC_7_20_5 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNI4N6K_2_LC_7_20_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \dron_frame_decoder_1.state_RNI4N6K_2_LC_7_20_5  (
            .in0(N__48558),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43409),
            .lcout(\dron_frame_decoder_1.state_RNI4N6KZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.count_0_LC_7_20_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.count_0_LC_7_20_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.count_0_LC_7_20_6 .LUT_INIT=16'b0001010001010000;
    LogicCell40 \Commands_frame_decoder.count_0_LC_7_20_6  (
            .in0(N__71024),
            .in1(N__55279),
            .in2(N__41628),
            .in3(N__41227),
            .lcout(\Commands_frame_decoder.countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94353),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_4_LC_7_20_7 .C_ON=1'b0;
    defparam \uart_pc.state_4_LC_7_20_7 .SEQ_MODE=4'b1000;
    defparam \uart_pc.state_4_LC_7_20_7 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \uart_pc.state_4_LC_7_20_7  (
            .in0(N__41596),
            .in1(N__45796),
            .in2(N__41584),
            .in3(N__71025),
            .lcout(\uart_pc.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94353),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNO_0_1_LC_7_21_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_0_1_LC_7_21_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_0_1_LC_7_21_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Commands_frame_decoder.state_RNO_0_1_LC_7_21_3  (
            .in0(N__46402),
            .in1(N__88646),
            .in2(N__41551),
            .in3(N__92475),
            .lcout(\Commands_frame_decoder.state_ns_0_a3_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.state_RNI3OO4_0_LC_7_25_0 .C_ON=1'b0;
    defparam \pid_front.state_RNI3OO4_0_LC_7_25_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.state_RNI3OO4_0_LC_7_25_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pid_front.state_RNI3OO4_0_LC_7_25_0  (
            .in0(_gnd_net_),
            .in1(N__70606),
            .in2(_gnd_net_),
            .in3(N__86581),
            .lcout(\pid_front.state_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIO43R3_0_LC_8_1_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNIO43R3_0_LC_8_1_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIO43R3_0_LC_8_1_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIO43R3_0_LC_8_1_0  (
            .in0(_gnd_net_),
            .in1(N__44278),
            .in2(N__41503),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_1_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_1_LC_8_1_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_1_LC_8_1_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_1_LC_8_1_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_1_LC_8_1_1  (
            .in0(_gnd_net_),
            .in1(N__41494),
            .in2(_gnd_net_),
            .in3(N__41476),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_1 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_0 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_2_LC_8_1_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_2_LC_8_1_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_2_LC_8_1_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_2_LC_8_1_2  (
            .in0(_gnd_net_),
            .in1(N__43584),
            .in2(N__41473),
            .in3(N__41458),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_2 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_1 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_3_LC_8_1_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_3_LC_8_1_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_3_LC_8_1_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_3_LC_8_1_3  (
            .in0(_gnd_net_),
            .in1(N__41455),
            .in2(_gnd_net_),
            .in3(N__41437),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_3 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_2 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_4_LC_8_1_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_4_LC_8_1_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_4_LC_8_1_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_4_LC_8_1_4  (
            .in0(_gnd_net_),
            .in1(N__41434),
            .in2(_gnd_net_),
            .in3(N__41416),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_4 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_3 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_5_LC_8_1_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_5_LC_8_1_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_5_LC_8_1_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_5_LC_8_1_5  (
            .in0(_gnd_net_),
            .in1(N__41689),
            .in2(_gnd_net_),
            .in3(N__41683),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_5 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_4 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_6_LC_8_1_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_6_LC_8_1_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_6_LC_8_1_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_6_LC_8_1_6  (
            .in0(_gnd_net_),
            .in1(N__43924),
            .in2(N__43654),
            .in3(N__41680),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_6 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_5 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_7_LC_8_1_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_7_LC_8_1_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_7_LC_8_1_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_7_LC_8_1_7  (
            .in0(_gnd_net_),
            .in1(N__41677),
            .in2(_gnd_net_),
            .in3(N__41671),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_7 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_6 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_8_LC_8_2_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_8_LC_8_2_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_8_LC_8_2_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_8_LC_8_2_0  (
            .in0(_gnd_net_),
            .in1(N__41668),
            .in2(_gnd_net_),
            .in3(N__41662),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_8 ),
            .ltout(),
            .carryin(bfn_8_2_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_9_LC_8_2_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_9_LC_8_2_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_9_LC_8_2_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_9_LC_8_2_1  (
            .in0(_gnd_net_),
            .in1(N__41659),
            .in2(_gnd_net_),
            .in3(N__41653),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_9 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_8 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_10_LC_8_2_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_10_LC_8_2_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_10_LC_8_2_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_10_LC_8_2_2  (
            .in0(_gnd_net_),
            .in1(N__41650),
            .in2(_gnd_net_),
            .in3(N__41644),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_10 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_9 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_11_LC_8_2_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_11_LC_8_2_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_11_LC_8_2_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_11_LC_8_2_3  (
            .in0(_gnd_net_),
            .in1(N__41701),
            .in2(_gnd_net_),
            .in3(N__41641),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_11 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_10 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_12_LC_8_2_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_12_LC_8_2_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_12_LC_8_2_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_12_LC_8_2_4  (
            .in0(_gnd_net_),
            .in1(N__41638),
            .in2(_gnd_net_),
            .in3(N__41632),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_12 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_11 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_13_LC_8_2_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_13_LC_8_2_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_13_LC_8_2_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_13_LC_8_2_5  (
            .in0(_gnd_net_),
            .in1(N__44118),
            .in2(N__41830),
            .in3(N__41821),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_13 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_12 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_14_LC_8_2_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_14_LC_8_2_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_14_LC_8_2_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_14_LC_8_2_6  (
            .in0(_gnd_net_),
            .in1(N__41818),
            .in2(_gnd_net_),
            .in3(N__41812),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_14 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_13 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_15_LC_8_2_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_15_LC_8_2_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_15_LC_8_2_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_15_LC_8_2_7  (
            .in0(_gnd_net_),
            .in1(N__41809),
            .in2(_gnd_net_),
            .in3(N__41803),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_15 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_14 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_16_LC_8_3_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_16_LC_8_3_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_16_LC_8_3_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_16_LC_8_3_0  (
            .in0(_gnd_net_),
            .in1(N__46855),
            .in2(_gnd_net_),
            .in3(N__41800),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_16 ),
            .ltout(),
            .carryin(bfn_8_3_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_17_LC_8_3_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_17_LC_8_3_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_17_LC_8_3_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_17_LC_8_3_1  (
            .in0(_gnd_net_),
            .in1(N__41929),
            .in2(_gnd_net_),
            .in3(N__41797),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_17 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_16 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_18_LC_8_3_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNO_1_18_LC_8_3_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_18_LC_8_3_2 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_18_LC_8_3_2  (
            .in0(N__41789),
            .in1(N__49005),
            .in2(_gnd_net_),
            .in3(N__41704),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIQH131_11_LC_8_3_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIQH131_11_LC_8_3_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIQH131_11_LC_8_3_3 .LUT_INIT=16'b1111000001111000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIQH131_11_LC_8_3_3  (
            .in0(N__49645),
            .in1(N__56301),
            .in2(N__46807),
            .in3(N__52891),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI8L3H5_13_LC_8_3_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI8L3H5_13_LC_8_3_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI8L3H5_13_LC_8_3_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI8L3H5_13_LC_8_3_4  (
            .in0(N__44113),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41695),
            .lcout(\ppm_encoder_1.init_pulses_RNI8L3H5Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIUL131_15_LC_8_3_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIUL131_15_LC_8_3_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIUL131_15_LC_8_3_5 .LUT_INIT=16'b1111000001111000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIUL131_15_LC_8_3_5  (
            .in0(N__49646),
            .in1(N__56302),
            .in2(N__48804),
            .in3(N__52892),
            .lcout(\ppm_encoder_1.N_254_i_i ),
            .ltout(\ppm_encoder_1.N_254_i_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNILFR51_15_LC_8_3_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNILFR51_15_LC_8_3_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNILFR51_15_LC_8_3_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNILFR51_15_LC_8_3_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__41932),
            .in3(N__48799),
            .lcout(\ppm_encoder_1.init_pulses_RNILFR51Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI0O131_17_LC_8_3_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI0O131_17_LC_8_3_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI0O131_17_LC_8_3_7 .LUT_INIT=16'b1111000001111000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI0O131_17_LC_8_3_7  (
            .in0(N__49647),
            .in1(N__56303),
            .in2(N__49179),
            .in3(N__52893),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_16_LC_8_4_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_16_LC_8_4_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_16_LC_8_4_0 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \ppm_encoder_1.init_pulses_16_LC_8_4_0  (
            .in0(N__49482),
            .in1(N__49306),
            .in2(N__41923),
            .in3(N__44050),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94116),
            .ce(),
            .sr(N__86509));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNITL7J1_2_LC_8_4_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNITL7J1_2_LC_8_4_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNITL7J1_2_LC_8_4_1 .LUT_INIT=16'b1111111101100110;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_RNITL7J1_2_LC_8_4_1  (
            .in0(N__44692),
            .in1(N__56304),
            .in2(_gnd_net_),
            .in3(N__52868),
            .lcout(\ppm_encoder_1.N_298 ),
            .ltout(\ppm_encoder_1.N_298_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_10_LC_8_4_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_10_LC_8_4_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_10_LC_8_4_2 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \ppm_encoder_1.init_pulses_10_LC_8_4_2  (
            .in0(N__49480),
            .in1(N__41914),
            .in2(N__41905),
            .in3(N__43792),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94116),
            .ce(),
            .sr(N__86509));
    defparam \ppm_encoder_1.init_pulses_17_LC_8_4_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_17_LC_8_4_3 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_17_LC_8_4_3 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \ppm_encoder_1.init_pulses_17_LC_8_4_3  (
            .in0(N__49307),
            .in1(N__41902),
            .in2(N__49503),
            .in3(N__44029),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94116),
            .ce(),
            .sr(N__86509));
    defparam \ppm_encoder_1.init_pulses_18_LC_8_4_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_18_LC_8_4_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_18_LC_8_4_4 .LUT_INIT=16'b0000101100001000;
    LogicCell40 \ppm_encoder_1.init_pulses_18_LC_8_4_4  (
            .in0(N__41896),
            .in1(N__49308),
            .in2(N__49500),
            .in3(N__44017),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94116),
            .ce(),
            .sr(N__86509));
    defparam \ppm_encoder_1.init_pulses_13_LC_8_4_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_13_LC_8_4_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_13_LC_8_4_5 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \ppm_encoder_1.init_pulses_13_LC_8_4_5  (
            .in0(N__49303),
            .in1(N__41890),
            .in2(N__49501),
            .in3(N__44092),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94116),
            .ce(),
            .sr(N__86509));
    defparam \ppm_encoder_1.init_pulses_14_LC_8_4_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_14_LC_8_4_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_14_LC_8_4_6 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \ppm_encoder_1.init_pulses_14_LC_8_4_6  (
            .in0(N__49481),
            .in1(N__49304),
            .in2(N__41842),
            .in3(N__44083),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94116),
            .ce(),
            .sr(N__86509));
    defparam \ppm_encoder_1.init_pulses_15_LC_8_4_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_15_LC_8_4_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_15_LC_8_4_7 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \ppm_encoder_1.init_pulses_15_LC_8_4_7  (
            .in0(N__49305),
            .in1(N__42004),
            .in2(N__49502),
            .in3(N__44059),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94116),
            .ce(),
            .sr(N__86509));
    defparam \ppm_encoder_1.init_pulses_RNIJI261_0_LC_8_5_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIJI261_0_LC_8_5_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIJI261_0_LC_8_5_1 .LUT_INIT=16'b1111000001111000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIJI261_0_LC_8_5_1  (
            .in0(N__42205),
            .in1(N__41995),
            .in2(N__49246),
            .in3(N__52887),
            .lcout(\ppm_encoder_1.N_257_i_i ),
            .ltout(\ppm_encoder_1.N_257_i_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_0_LC_8_5_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNO_0_0_LC_8_5_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_0_LC_8_5_2 .LUT_INIT=16'b0000111100011110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_0_LC_8_5_2  (
            .in0(N__44305),
            .in1(N__44293),
            .in2(N__41959),
            .in3(N__44512),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIBC8E1_0_LC_8_5_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIBC8E1_0_LC_8_5_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIBC8E1_0_LC_8_5_3 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \ppm_encoder_1.throttle_RNIBC8E1_0_LC_8_5_3  (
            .in0(N__44678),
            .in1(N__42269),
            .in2(N__42255),
            .in3(N__44596),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIG7561_0_LC_8_5_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIG7561_0_LC_8_5_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIG7561_0_LC_8_5_5 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \ppm_encoder_1.elevator_RNIG7561_0_LC_8_5_5  (
            .in0(N__47230),
            .in1(N__42204),
            .in2(_gnd_net_),
            .in3(N__47437),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_0_LC_8_5_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_0_LC_8_5_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_0_LC_8_5_6 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \ppm_encoder_1.aileron_0_LC_8_5_6  (
            .in0(N__42270),
            .in1(N__51346),
            .in2(_gnd_net_),
            .in3(N__59175),
            .lcout(\ppm_encoder_1.aileronZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94124),
            .ce(),
            .sr(N__86506));
    defparam \ppm_encoder_1.throttle_0_LC_8_5_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_0_LC_8_5_7 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.throttle_0_LC_8_5_7 .LUT_INIT=16'b0000101011111010;
    LogicCell40 \ppm_encoder_1.throttle_0_LC_8_5_7  (
            .in0(N__42251),
            .in1(_gnd_net_),
            .in2(N__51374),
            .in3(N__41956),
            .lcout(\ppm_encoder_1.throttleZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94124),
            .ce(),
            .sr(N__86506));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNIUTMR_LC_8_6_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNIUTMR_LC_8_6_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNIUTMR_LC_8_6_0 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNIUTMR_LC_8_6_0  (
            .in0(N__42208),
            .in1(N__42091),
            .in2(_gnd_net_),
            .in3(N__44923),
            .lcout(\ppm_encoder_1.N_514 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNINKS41_10_LC_8_6_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNINKS41_10_LC_8_6_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNINKS41_10_LC_8_6_1 .LUT_INIT=16'b1111000001111000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNINKS41_10_LC_8_6_1  (
            .in0(N__53780),
            .in1(N__53644),
            .in2(N__50117),
            .in3(N__52883),
            .lcout(\ppm_encoder_1.N_255_i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep2_LC_8_6_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep2_LC_8_6_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep2_LC_8_6_2 .LUT_INIT=16'b0000000010110001;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_2_rep2_LC_8_6_2  (
            .in0(N__52884),
            .in1(N__47135),
            .in2(N__53681),
            .in3(N__71037),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94133),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIOLS41_0_11_LC_8_6_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIOLS41_0_11_LC_8_6_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIOLS41_0_11_LC_8_6_3 .LUT_INIT=16'b0000111110000111;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIOLS41_0_11_LC_8_6_3  (
            .in0(N__53779),
            .in1(N__53643),
            .in2(N__46803),
            .in3(N__52882),
            .lcout(\ppm_encoder_1.N_266_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_0_LC_8_6_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_0_LC_8_6_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_0_LC_8_6_4 .LUT_INIT=16'b0010001011000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_0_LC_8_6_4  (
            .in0(N__42271),
            .in1(N__54194),
            .in2(N__42256),
            .in3(N__54074),
            .lcout(\ppm_encoder_1.pulses2count_9_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_10_LC_8_6_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_10_LC_8_6_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_10_LC_8_6_5 .LUT_INIT=16'b0010001000001010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_10_LC_8_6_5  (
            .in0(N__54075),
            .in1(N__42430),
            .in2(N__42235),
            .in3(N__54195),
            .lcout(\ppm_encoder_1.pulses2count_9_i_0_1_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNIUTMR_0_LC_8_6_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNIUTMR_0_LC_8_6_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNIUTMR_0_LC_8_6_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNIUTMR_0_LC_8_6_6  (
            .in0(N__42207),
            .in1(N__42090),
            .in2(_gnd_net_),
            .in3(N__44922),
            .lcout(\ppm_encoder_1.N_508 ),
            .ltout(\ppm_encoder_1.N_508_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_0_LC_8_6_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_0_LC_8_6_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_0_LC_8_6_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_0_LC_8_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42037),
            .in3(N__49245),
            .lcout(\ppm_encoder_1.N_393 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_11_LC_8_7_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_11_LC_8_7_0 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_11_LC_8_7_0 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.aileron_11_LC_8_7_0  (
            .in0(N__54483),
            .in1(N__48022),
            .in2(N__50184),
            .in3(N__51317),
            .lcout(\ppm_encoder_1.aileronZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94139),
            .ce(),
            .sr(N__86498));
    defparam \ppm_encoder_1.elevator_3_LC_8_7_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_3_LC_8_7_1 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_3_LC_8_7_1 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \ppm_encoder_1.elevator_3_LC_8_7_1  (
            .in0(N__47260),
            .in1(N__60061),
            .in2(N__51366),
            .in3(N__47549),
            .lcout(\ppm_encoder_1.elevatorZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94139),
            .ce(),
            .sr(N__86498));
    defparam \ppm_encoder_1.throttle_12_LC_8_7_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_12_LC_8_7_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_12_LC_8_7_3 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.throttle_12_LC_8_7_3  (
            .in0(N__42034),
            .in1(N__42016),
            .in2(N__51367),
            .in3(N__47720),
            .lcout(\ppm_encoder_1.throttleZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94139),
            .ce(),
            .sr(N__86498));
    defparam \ppm_encoder_1.aileron_12_LC_8_7_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_12_LC_8_7_4 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_12_LC_8_7_4 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.aileron_12_LC_8_7_4  (
            .in0(N__53184),
            .in1(N__48007),
            .in2(N__50700),
            .in3(N__51318),
            .lcout(\ppm_encoder_1.aileronZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94139),
            .ce(),
            .sr(N__86498));
    defparam \ppm_encoder_1.aileron_2_LC_8_7_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_2_LC_8_7_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_2_LC_8_7_5 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.aileron_2_LC_8_7_5  (
            .in0(N__47686),
            .in1(N__56035),
            .in2(N__51365),
            .in3(N__50630),
            .lcout(\ppm_encoder_1.aileronZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94139),
            .ce(),
            .sr(N__86498));
    defparam \ppm_encoder_1.aileron_1_LC_8_7_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_1_LC_8_7_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_1_LC_8_7_6 .LUT_INIT=16'b1001100111110000;
    LogicCell40 \ppm_encoder_1.aileron_1_LC_8_7_6  (
            .in0(N__56059),
            .in1(N__47701),
            .in2(N__50234),
            .in3(N__51319),
            .lcout(\ppm_encoder_1.aileronZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94139),
            .ce(),
            .sr(N__86498));
    defparam \ppm_encoder_1.elevator_10_LC_8_8_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_10_LC_8_8_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_10_LC_8_8_0 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.elevator_10_LC_8_8_0  (
            .in0(N__54676),
            .in1(N__47626),
            .in2(N__42429),
            .in3(N__51261),
            .lcout(\ppm_encoder_1.elevatorZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94152),
            .ce(),
            .sr(N__86492));
    defparam \ppm_encoder_1.aileron_3_LC_8_8_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_3_LC_8_8_7 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_3_LC_8_8_7 .LUT_INIT=16'b1101100001110010;
    LogicCell40 \ppm_encoder_1.aileron_3_LC_8_8_7  (
            .in0(N__51260),
            .in1(N__56008),
            .in2(N__50414),
            .in3(N__47854),
            .lcout(\ppm_encoder_1.aileronZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94152),
            .ce(),
            .sr(N__86492));
    defparam \ppm_encoder_1.aileron_9_LC_8_9_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_9_LC_8_9_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_9_LC_8_9_0 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.aileron_9_LC_8_9_0  (
            .in0(N__54349),
            .in1(N__47773),
            .in2(N__51353),
            .in3(N__44754),
            .lcout(\ppm_encoder_1.aileronZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94163),
            .ce(),
            .sr(N__86487));
    defparam \ppm_encoder_1.rudder_8_LC_8_9_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_8_LC_8_9_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_8_LC_8_9_1 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.rudder_8_LC_8_9_1  (
            .in0(N__42403),
            .in1(N__42397),
            .in2(N__46994),
            .in3(N__51288),
            .lcout(\ppm_encoder_1.rudderZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94163),
            .ce(),
            .sr(N__86487));
    defparam \ppm_encoder_1.elevator_13_LC_8_9_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_13_LC_8_9_3 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_13_LC_8_9_3 .LUT_INIT=16'b1001100111110000;
    LogicCell40 \ppm_encoder_1.elevator_13_LC_8_9_3  (
            .in0(N__55750),
            .in1(N__47584),
            .in2(N__42374),
            .in3(N__51285),
            .lcout(\ppm_encoder_1.elevatorZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94163),
            .ce(),
            .sr(N__86487));
    defparam \ppm_encoder_1.rudder_10_LC_8_9_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_10_LC_8_9_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_10_LC_8_9_4 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.rudder_10_LC_8_9_4  (
            .in0(N__42346),
            .in1(N__42340),
            .in2(N__51354),
            .in3(N__47084),
            .lcout(\ppm_encoder_1.rudderZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94163),
            .ce(),
            .sr(N__86487));
    defparam \ppm_encoder_1.rudder_13_LC_8_9_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_13_LC_8_9_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.rudder_13_LC_8_9_5 .LUT_INIT=16'b1001100111110000;
    LogicCell40 \ppm_encoder_1.rudder_13_LC_8_9_5  (
            .in0(N__42325),
            .in1(N__42319),
            .in2(N__42297),
            .in3(N__51287),
            .lcout(\ppm_encoder_1.rudderZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94163),
            .ce(),
            .sr(N__86487));
    defparam \ppm_encoder_1.rudder_12_LC_8_9_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_12_LC_8_9_7 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.rudder_12_LC_8_9_7 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.rudder_12_LC_8_9_7  (
            .in0(N__42475),
            .in1(N__42460),
            .in2(N__42454),
            .in3(N__51286),
            .lcout(\ppm_encoder_1.rudderZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94163),
            .ce(),
            .sr(N__86487));
    defparam \Commands_frame_decoder.source_CH4data_esr_0_LC_8_10_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_0_LC_8_10_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_0_LC_8_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_0_LC_8_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88281),
            .lcout(frame_decoder_CH4data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94176),
            .ce(N__45886),
            .sr(N__86480));
    defparam \Commands_frame_decoder.source_CH4data_esr_1_LC_8_10_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_1_LC_8_10_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_1_LC_8_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_1_LC_8_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85509),
            .lcout(frame_decoder_CH4data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94176),
            .ce(N__45886),
            .sr(N__86480));
    defparam \Commands_frame_decoder.source_CH4data_esr_2_LC_8_10_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_2_LC_8_10_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_2_LC_8_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_2_LC_8_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__92515),
            .lcout(frame_decoder_CH4data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94176),
            .ce(N__45886),
            .sr(N__86480));
    defparam \Commands_frame_decoder.source_CH4data_esr_3_LC_8_10_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_3_LC_8_10_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_3_LC_8_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_3_LC_8_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__92283),
            .lcout(frame_decoder_CH4data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94176),
            .ce(N__45886),
            .sr(N__86480));
    defparam \Commands_frame_decoder.source_CH4data_esr_4_LC_8_10_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_4_LC_8_10_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_4_LC_8_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_4_LC_8_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88813),
            .lcout(frame_decoder_CH4data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94176),
            .ce(N__45886),
            .sr(N__86480));
    defparam \Commands_frame_decoder.source_CH4data_esr_5_LC_8_10_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_5_LC_8_10_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_5_LC_8_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_5_LC_8_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88664),
            .lcout(frame_decoder_CH4data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94176),
            .ce(N__45886),
            .sr(N__86480));
    defparam \Commands_frame_decoder.source_CH4data_esr_6_LC_8_10_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_6_LC_8_10_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_6_LC_8_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_6_LC_8_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88481),
            .lcout(frame_decoder_CH4data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94176),
            .ce(N__45886),
            .sr(N__86480));
    defparam \Commands_frame_decoder.source_CH4data_ess_7_LC_8_10_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_ess_7_LC_8_10_7 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_CH4data_ess_7_LC_8_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_ess_7_LC_8_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__92065),
            .lcout(frame_decoder_CH4data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94176),
            .ce(N__45886),
            .sr(N__86480));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_LC_8_11_0 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_LC_8_11_0 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_LC_8_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_LC_8_11_0  (
            .in0(_gnd_net_),
            .in1(N__45235),
            .in2(N__45184),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_11_0_),
            .carryout(\scaler_4.un3_source_data_0_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_RNI40BL_LC_8_11_1 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_RNI40BL_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_RNI40BL_LC_8_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_RNI40BL_LC_8_11_1  (
            .in0(_gnd_net_),
            .in1(N__42619),
            .in2(N__45451),
            .in3(N__42613),
            .lcout(\scaler_4.un2_source_data_0 ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_0 ),
            .carryout(\scaler_4.un3_source_data_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_1_c_RNI74CL_LC_8_11_2 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_1_c_RNI74CL_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_1_c_RNI74CL_LC_8_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_1_c_RNI74CL_LC_8_11_2  (
            .in0(_gnd_net_),
            .in1(N__42610),
            .in2(N__45439),
            .in3(N__42592),
            .lcout(\scaler_4.un3_source_data_0_cry_1_c_RNI74CL ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_1 ),
            .carryout(\scaler_4.un3_source_data_0_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_2_c_RNIA8DL_LC_8_11_3 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_2_c_RNIA8DL_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_2_c_RNIA8DL_LC_8_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_2_c_RNIA8DL_LC_8_11_3  (
            .in0(_gnd_net_),
            .in1(N__42589),
            .in2(N__45427),
            .in3(N__42571),
            .lcout(\scaler_4.un3_source_data_0_cry_2_c_RNIA8DL ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_2 ),
            .carryout(\scaler_4.un3_source_data_0_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_3_c_RNIDCEL_LC_8_11_4 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_3_c_RNIDCEL_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_3_c_RNIDCEL_LC_8_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_3_c_RNIDCEL_LC_8_11_4  (
            .in0(_gnd_net_),
            .in1(N__42568),
            .in2(N__45415),
            .in3(N__42550),
            .lcout(\scaler_4.un3_source_data_0_cry_3_c_RNIDCEL ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_3 ),
            .carryout(\scaler_4.un3_source_data_0_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_4_c_RNIGGFL_LC_8_11_5 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_4_c_RNIGGFL_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_4_c_RNIGGFL_LC_8_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_4_c_RNIGGFL_LC_8_11_5  (
            .in0(_gnd_net_),
            .in1(N__42547),
            .in2(N__45403),
            .in3(N__42529),
            .lcout(\scaler_4.un3_source_data_0_cry_4_c_RNIGGFL ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_4 ),
            .carryout(\scaler_4.un3_source_data_0_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_5_c_RNIJKGL_LC_8_11_6 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_5_c_RNIJKGL_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_5_c_RNIJKGL_LC_8_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_5_c_RNIJKGL_LC_8_11_6  (
            .in0(_gnd_net_),
            .in1(N__42526),
            .in2(N__45391),
            .in3(N__42508),
            .lcout(\scaler_4.un3_source_data_0_cry_5_c_RNIJKGL ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_5 ),
            .carryout(\scaler_4.un3_source_data_0_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_6_c_RNIOUNN_LC_8_11_7 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_6_c_RNIOUNN_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_6_c_RNIOUNN_LC_8_11_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_6_c_RNIOUNN_LC_8_11_7  (
            .in0(_gnd_net_),
            .in1(N__42715),
            .in2(_gnd_net_),
            .in3(N__42493),
            .lcout(\scaler_4.un3_source_data_0_cry_6_c_RNIOUNN ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_6 ),
            .carryout(\scaler_4.un3_source_data_0_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_7_c_RNIP0PN_LC_8_12_0 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_7_c_RNIP0PN_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_7_c_RNIP0PN_LC_8_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_7_c_RNIP0PN_LC_8_12_0  (
            .in0(_gnd_net_),
            .in1(N__46174),
            .in2(N__65858),
            .in3(N__42478),
            .lcout(\scaler_4.un3_source_data_0_cry_7_c_RNIP0PN ),
            .ltout(),
            .carryin(bfn_8_12_0_),
            .carryout(\scaler_4.un3_source_data_0_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_8_c_RNIS918_LC_8_12_1 .C_ON=1'b0;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_8_c_RNIS918_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_8_c_RNIS918_LC_8_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_8_c_RNIS918_LC_8_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42751),
            .lcout(\scaler_4.un3_source_data_0_cry_8_c_RNIS918 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIQRI31_10_LC_8_12_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIQRI31_10_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIQRI31_10_LC_8_12_2 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \Commands_frame_decoder.state_RNIQRI31_10_LC_8_12_2  (
            .in0(N__48261),
            .in1(N__55280),
            .in2(_gnd_net_),
            .in3(N__70843),
            .lcout(\Commands_frame_decoder.state_RNIQRI31Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_axb_7_LC_8_12_6 .C_ON=1'b0;
    defparam \scaler_4.un3_source_data_un3_source_data_0_axb_7_LC_8_12_6 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_axb_7_LC_8_12_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_axb_7_LC_8_12_6  (
            .in0(_gnd_net_),
            .in1(N__46206),
            .in2(_gnd_net_),
            .in3(N__46191),
            .lcout(\scaler_4.un3_source_data_0_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_0_LC_8_13_0 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_0_LC_8_13_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_0_LC_8_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_0_LC_8_13_0  (
            .in0(_gnd_net_),
            .in1(N__42691),
            .in2(N__42708),
            .in3(N__42709),
            .lcout(\Commands_frame_decoder.WDTZ0Z_0 ),
            .ltout(),
            .carryin(bfn_8_13_0_),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_0 ),
            .clk(N__94222),
            .ce(),
            .sr(N__55101));
    defparam \Commands_frame_decoder.WDT_1_LC_8_13_1 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_1_LC_8_13_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_1_LC_8_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_1_LC_8_13_1  (
            .in0(_gnd_net_),
            .in1(N__42685),
            .in2(_gnd_net_),
            .in3(N__42679),
            .lcout(\Commands_frame_decoder.WDTZ0Z_1 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_0 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_1 ),
            .clk(N__94222),
            .ce(),
            .sr(N__55101));
    defparam \Commands_frame_decoder.WDT_2_LC_8_13_2 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_2_LC_8_13_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_2_LC_8_13_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_2_LC_8_13_2  (
            .in0(_gnd_net_),
            .in1(N__42676),
            .in2(_gnd_net_),
            .in3(N__42670),
            .lcout(\Commands_frame_decoder.WDTZ0Z_2 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_1 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_2 ),
            .clk(N__94222),
            .ce(),
            .sr(N__55101));
    defparam \Commands_frame_decoder.WDT_3_LC_8_13_3 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_3_LC_8_13_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_3_LC_8_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_3_LC_8_13_3  (
            .in0(_gnd_net_),
            .in1(N__42667),
            .in2(_gnd_net_),
            .in3(N__42661),
            .lcout(\Commands_frame_decoder.WDTZ0Z_3 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_2 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_3 ),
            .clk(N__94222),
            .ce(),
            .sr(N__55101));
    defparam \Commands_frame_decoder.WDT_4_LC_8_13_4 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_4_LC_8_13_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_4_LC_8_13_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_4_LC_8_13_4  (
            .in0(_gnd_net_),
            .in1(N__42658),
            .in2(_gnd_net_),
            .in3(N__42640),
            .lcout(\Commands_frame_decoder.WDTZ0Z_4 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_3 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_4 ),
            .clk(N__94222),
            .ce(),
            .sr(N__55101));
    defparam \Commands_frame_decoder.WDT_5_LC_8_13_5 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_5_LC_8_13_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_5_LC_8_13_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_5_LC_8_13_5  (
            .in0(_gnd_net_),
            .in1(N__42637),
            .in2(_gnd_net_),
            .in3(N__42934),
            .lcout(\Commands_frame_decoder.WDTZ0Z_5 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_4 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_5 ),
            .clk(N__94222),
            .ce(),
            .sr(N__55101));
    defparam \Commands_frame_decoder.WDT_6_LC_8_13_6 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_6_LC_8_13_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_6_LC_8_13_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_6_LC_8_13_6  (
            .in0(_gnd_net_),
            .in1(N__42931),
            .in2(_gnd_net_),
            .in3(N__42913),
            .lcout(\Commands_frame_decoder.WDTZ0Z_6 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_5 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_6 ),
            .clk(N__94222),
            .ce(),
            .sr(N__55101));
    defparam \Commands_frame_decoder.WDT_7_LC_8_13_7 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_7_LC_8_13_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_7_LC_8_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_7_LC_8_13_7  (
            .in0(_gnd_net_),
            .in1(N__42908),
            .in2(_gnd_net_),
            .in3(N__42886),
            .lcout(\Commands_frame_decoder.WDTZ0Z_7 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_6 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_7 ),
            .clk(N__94222),
            .ce(),
            .sr(N__55101));
    defparam \Commands_frame_decoder.WDT_8_LC_8_14_0 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_8_LC_8_14_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_8_LC_8_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_8_LC_8_14_0  (
            .in0(_gnd_net_),
            .in1(N__42883),
            .in2(_gnd_net_),
            .in3(N__42868),
            .lcout(\Commands_frame_decoder.WDTZ0Z_8 ),
            .ltout(),
            .carryin(bfn_8_14_0_),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_8 ),
            .clk(N__94239),
            .ce(),
            .sr(N__55105));
    defparam \Commands_frame_decoder.WDT_9_LC_8_14_1 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_9_LC_8_14_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_9_LC_8_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_9_LC_8_14_1  (
            .in0(_gnd_net_),
            .in1(N__42864),
            .in2(_gnd_net_),
            .in3(N__42847),
            .lcout(\Commands_frame_decoder.WDTZ0Z_9 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_8 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_9 ),
            .clk(N__94239),
            .ce(),
            .sr(N__55105));
    defparam \Commands_frame_decoder.WDT_10_LC_8_14_2 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_10_LC_8_14_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_10_LC_8_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_10_LC_8_14_2  (
            .in0(_gnd_net_),
            .in1(N__42844),
            .in2(_gnd_net_),
            .in3(N__42826),
            .lcout(\Commands_frame_decoder.WDTZ0Z_10 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_9 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_10 ),
            .clk(N__94239),
            .ce(),
            .sr(N__55105));
    defparam \Commands_frame_decoder.WDT_11_LC_8_14_3 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_11_LC_8_14_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_11_LC_8_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_11_LC_8_14_3  (
            .in0(_gnd_net_),
            .in1(N__42823),
            .in2(_gnd_net_),
            .in3(N__42802),
            .lcout(\Commands_frame_decoder.WDTZ0Z_11 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_10 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_11 ),
            .clk(N__94239),
            .ce(),
            .sr(N__55105));
    defparam \Commands_frame_decoder.WDT_12_LC_8_14_4 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_12_LC_8_14_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_12_LC_8_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_12_LC_8_14_4  (
            .in0(_gnd_net_),
            .in1(N__42798),
            .in2(_gnd_net_),
            .in3(N__42775),
            .lcout(\Commands_frame_decoder.WDTZ0Z_12 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_11 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_12 ),
            .clk(N__94239),
            .ce(),
            .sr(N__55105));
    defparam \Commands_frame_decoder.WDT_13_LC_8_14_5 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_13_LC_8_14_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_13_LC_8_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_13_LC_8_14_5  (
            .in0(_gnd_net_),
            .in1(N__42772),
            .in2(_gnd_net_),
            .in3(N__42754),
            .lcout(\Commands_frame_decoder.WDTZ0Z_13 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_12 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_13 ),
            .clk(N__94239),
            .ce(),
            .sr(N__55105));
    defparam \Commands_frame_decoder.WDT_14_LC_8_14_6 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_14_LC_8_14_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_14_LC_8_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_14_LC_8_14_6  (
            .in0(_gnd_net_),
            .in1(N__48291),
            .in2(_gnd_net_),
            .in3(N__42961),
            .lcout(\Commands_frame_decoder.WDTZ0Z_14 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_13 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_14 ),
            .clk(N__94239),
            .ce(),
            .sr(N__55105));
    defparam \Commands_frame_decoder.WDT_15_LC_8_14_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_15_LC_8_14_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_15_LC_8_14_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Commands_frame_decoder.WDT_15_LC_8_14_7  (
            .in0(_gnd_net_),
            .in1(N__48326),
            .in2(_gnd_net_),
            .in3(N__42958),
            .lcout(\Commands_frame_decoder.WDTZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94239),
            .ce(),
            .sr(N__55105));
    defparam \scaler_4.source_data_1_esr_5_LC_8_15_0 .C_ON=1'b0;
    defparam \scaler_4.source_data_1_esr_5_LC_8_15_0 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_5_LC_8_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \scaler_4.source_data_1_esr_5_LC_8_15_0  (
            .in0(N__45183),
            .in1(N__45268),
            .in2(_gnd_net_),
            .in3(N__45241),
            .lcout(scaler_4_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94256),
            .ce(N__48062),
            .sr(N__86451));
    defparam \uart_pc.bit_Count_RNI4U6E1_2_LC_8_15_1 .C_ON=1'b0;
    defparam \uart_pc.bit_Count_RNI4U6E1_2_LC_8_15_1 .SEQ_MODE=4'b0000;
    defparam \uart_pc.bit_Count_RNI4U6E1_2_LC_8_15_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uart_pc.bit_Count_RNI4U6E1_2_LC_8_15_1  (
            .in0(N__42989),
            .in1(N__43074),
            .in2(_gnd_net_),
            .in3(N__43024),
            .lcout(\uart_pc.N_152 ),
            .ltout(\uart_pc.N_152_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIUPE73_3_LC_8_15_2 .C_ON=1'b0;
    defparam \uart_pc.state_RNIUPE73_3_LC_8_15_2 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIUPE73_3_LC_8_15_2 .LUT_INIT=16'b1111001100000000;
    LogicCell40 \uart_pc.state_RNIUPE73_3_LC_8_15_2  (
            .in0(_gnd_net_),
            .in1(N__45785),
            .in2(N__42937),
            .in3(N__43099),
            .lcout(\uart_pc.un1_state_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_0_LC_8_15_3 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_0_LC_8_15_3 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_0_LC_8_15_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \uart_pc.data_Aux_RNO_0_0_LC_8_15_3  (
            .in0(N__42992),
            .in1(N__43075),
            .in2(_gnd_net_),
            .in3(N__43025),
            .lcout(\uart_pc.data_Auxce_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_1_LC_8_15_4 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_1_LC_8_15_4 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_1_LC_8_15_4 .LUT_INIT=16'b0000000000001010;
    LogicCell40 \uart_pc.data_Aux_RNO_0_1_LC_8_15_4  (
            .in0(N__43076),
            .in1(_gnd_net_),
            .in2(N__43042),
            .in3(N__42991),
            .lcout(\uart_pc.data_Auxce_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_2_LC_8_15_5 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_2_LC_8_15_5 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_2_LC_8_15_5 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \uart_pc.data_Aux_RNO_0_2_LC_8_15_5  (
            .in0(N__42993),
            .in1(N__43077),
            .in2(_gnd_net_),
            .in3(N__43029),
            .lcout(\uart_pc.data_Auxce_0_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_3_LC_8_15_6 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_3_LC_8_15_6 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_3_LC_8_15_6 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \uart_pc.data_Aux_RNO_0_3_LC_8_15_6  (
            .in0(N__43078),
            .in1(_gnd_net_),
            .in2(N__43043),
            .in3(N__42990),
            .lcout(\uart_pc.data_Auxce_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_4_LC_8_15_7 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_4_LC_8_15_7 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_4_LC_8_15_7 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \uart_pc.data_Aux_RNO_0_4_LC_8_15_7  (
            .in0(N__42994),
            .in1(N__43079),
            .in2(_gnd_net_),
            .in3(N__43033),
            .lcout(\uart_pc.data_Auxce_0_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.bit_Count_0_LC_8_16_0 .C_ON=1'b0;
    defparam \uart_pc.bit_Count_0_LC_8_16_0 .SEQ_MODE=4'b1000;
    defparam \uart_pc.bit_Count_0_LC_8_16_0 .LUT_INIT=16'b0100011001000100;
    LogicCell40 \uart_pc.bit_Count_0_LC_8_16_0  (
            .in0(N__43101),
            .in1(N__43083),
            .in2(N__45541),
            .in3(N__45790),
            .lcout(\uart_pc.bit_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94275),
            .ce(),
            .sr(N__86448));
    defparam \uart_pc.bit_Count_RNO_0_2_LC_8_16_1 .C_ON=1'b0;
    defparam \uart_pc.bit_Count_RNO_0_2_LC_8_16_1 .SEQ_MODE=4'b0000;
    defparam \uart_pc.bit_Count_RNO_0_2_LC_8_16_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uart_pc.bit_Count_RNO_0_2_LC_8_16_1  (
            .in0(N__43082),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43100),
            .lcout(),
            .ltout(\uart_pc.CO0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.bit_Count_2_LC_8_16_2 .C_ON=1'b0;
    defparam \uart_pc.bit_Count_2_LC_8_16_2 .SEQ_MODE=4'b1000;
    defparam \uart_pc.bit_Count_2_LC_8_16_2 .LUT_INIT=16'b0001010001000100;
    LogicCell40 \uart_pc.bit_Count_2_LC_8_16_2  (
            .in0(N__43111),
            .in1(N__42997),
            .in2(N__43114),
            .in3(N__43041),
            .lcout(\uart_pc.bit_CountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94275),
            .ce(),
            .sr(N__86448));
    defparam \uart_pc.bit_Count_1_LC_8_16_3 .C_ON=1'b0;
    defparam \uart_pc.bit_Count_1_LC_8_16_3 .SEQ_MODE=4'b1000;
    defparam \uart_pc.bit_Count_1_LC_8_16_3 .LUT_INIT=16'b0001001000110000;
    LogicCell40 \uart_pc.bit_Count_1_LC_8_16_3  (
            .in0(N__43084),
            .in1(N__43110),
            .in2(N__43045),
            .in3(N__43102),
            .lcout(\uart_pc.bit_CountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94275),
            .ce(),
            .sr(N__86448));
    defparam \uart_pc.data_Aux_RNO_0_5_LC_8_16_4 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_5_LC_8_16_4 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_5_LC_8_16_4 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \uart_pc.data_Aux_RNO_0_5_LC_8_16_4  (
            .in0(N__42995),
            .in1(N__43034),
            .in2(_gnd_net_),
            .in3(N__43080),
            .lcout(\uart_pc.data_Auxce_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_6_LC_8_16_5 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_6_LC_8_16_5 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_6_LC_8_16_5 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \uart_pc.data_Aux_RNO_0_6_LC_8_16_5  (
            .in0(N__43081),
            .in1(_gnd_net_),
            .in2(N__43044),
            .in3(N__42996),
            .lcout(\uart_pc.data_Auxce_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIEAGS_4_LC_8_16_6 .C_ON=1'b0;
    defparam \uart_pc.state_RNIEAGS_4_LC_8_16_6 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIEAGS_4_LC_8_16_6 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \uart_pc.state_RNIEAGS_4_LC_8_16_6  (
            .in0(N__45856),
            .in1(N__45789),
            .in2(_gnd_net_),
            .in3(N__70960),
            .lcout(\uart_pc.state_RNIEAGSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_6_LC_8_17_0 .C_ON=1'b0;
    defparam \uart_pc.data_6_LC_8_17_0 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_6_LC_8_17_0 .LUT_INIT=16'b0101110100001000;
    LogicCell40 \uart_pc.data_6_LC_8_17_0  (
            .in0(N__46265),
            .in1(N__45520),
            .in2(N__45918),
            .in3(N__92052),
            .lcout(uart_pc_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94291),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNILR1B2_2_LC_8_17_1 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNILR1B2_2_LC_8_17_1 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNILR1B2_2_LC_8_17_1 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \uart_pc.timer_Count_RNILR1B2_2_LC_8_17_1  (
            .in0(N__70981),
            .in1(N__52225),
            .in2(_gnd_net_),
            .in3(N__52124),
            .lcout(\uart_pc.timer_Count_RNILR1B2Z0Z_2 ),
            .ltout(\uart_pc.timer_Count_RNILR1B2Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_4_LC_8_17_2 .C_ON=1'b0;
    defparam \uart_pc.data_4_LC_8_17_2 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_4_LC_8_17_2 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \uart_pc.data_4_LC_8_17_2  (
            .in0(N__52125),
            .in1(N__45697),
            .in2(N__43165),
            .in3(N__88768),
            .lcout(uart_pc_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94291),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_ns_i_a2_2_1_0_LC_8_17_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_ns_i_a2_2_1_0_LC_8_17_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_ns_i_a2_2_1_0_LC_8_17_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_ns_i_a2_2_1_0_LC_8_17_3  (
            .in0(_gnd_net_),
            .in1(N__88392),
            .in2(_gnd_net_),
            .in3(N__92191),
            .lcout(),
            .ltout(\Commands_frame_decoder.state_ns_i_a2_2_1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_ns_i_a2_2_0_LC_8_17_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_ns_i_a2_2_0_LC_8_17_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_ns_i_a2_2_0_LC_8_17_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Commands_frame_decoder.state_ns_i_a2_2_0_LC_8_17_4  (
            .in0(N__55254),
            .in1(N__88767),
            .in2(N__43162),
            .in3(N__85414),
            .lcout(\Commands_frame_decoder.N_410 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_5_LC_8_17_5 .C_ON=1'b0;
    defparam \uart_pc.data_5_LC_8_17_5 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_5_LC_8_17_5 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \uart_pc.data_5_LC_8_17_5  (
            .in0(N__46033),
            .in1(N__46266),
            .in2(N__88457),
            .in3(N__45908),
            .lcout(uart_pc_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94291),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNIMQ8T1_2_LC_8_17_6 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNIMQ8T1_2_LC_8_17_6 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNIMQ8T1_2_LC_8_17_6 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \uart_pc.timer_Count_RNIMQ8T1_2_LC_8_17_6  (
            .in0(N__52123),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70980),
            .lcout(\uart_pc.timer_Count_RNIMQ8T1Z0Z_2 ),
            .ltout(\uart_pc.timer_Count_RNIMQ8T1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_3_LC_8_17_7 .C_ON=1'b0;
    defparam \uart_pc.data_3_LC_8_17_7 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_3_LC_8_17_7 .LUT_INIT=16'b0010111100100000;
    LogicCell40 \uart_pc.data_3_LC_8_17_7  (
            .in0(N__45714),
            .in1(N__45907),
            .in2(N__43141),
            .in3(N__92192),
            .lcout(uart_pc_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94291),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_0_LC_8_18_0 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_0_LC_8_18_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_0_LC_8_18_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_0_LC_8_18_0  (
            .in0(_gnd_net_),
            .in1(N__43138),
            .in2(N__43300),
            .in3(N__43299),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_0 ),
            .ltout(),
            .carryin(bfn_8_18_0_),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_0 ),
            .clk(N__94306),
            .ce(),
            .sr(N__43375));
    defparam \dron_frame_decoder_1.WDT_1_LC_8_18_1 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_1_LC_8_18_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_1_LC_8_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_1_LC_8_18_1  (
            .in0(_gnd_net_),
            .in1(N__43132),
            .in2(_gnd_net_),
            .in3(N__43126),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_1 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_0 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_1 ),
            .clk(N__94306),
            .ce(),
            .sr(N__43375));
    defparam \dron_frame_decoder_1.WDT_2_LC_8_18_2 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_2_LC_8_18_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_2_LC_8_18_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_2_LC_8_18_2  (
            .in0(_gnd_net_),
            .in1(N__43123),
            .in2(_gnd_net_),
            .in3(N__43117),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_2 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_1 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_2 ),
            .clk(N__94306),
            .ce(),
            .sr(N__43375));
    defparam \dron_frame_decoder_1.WDT_3_LC_8_18_3 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_3_LC_8_18_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_3_LC_8_18_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_3_LC_8_18_3  (
            .in0(_gnd_net_),
            .in1(N__43198),
            .in2(_gnd_net_),
            .in3(N__43192),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_3 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_2 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_3 ),
            .clk(N__94306),
            .ce(),
            .sr(N__43375));
    defparam \dron_frame_decoder_1.WDT_4_LC_8_18_4 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_4_LC_8_18_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_4_LC_8_18_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_4_LC_8_18_4  (
            .in0(_gnd_net_),
            .in1(N__43233),
            .in2(_gnd_net_),
            .in3(N__43189),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_4 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_3 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_4 ),
            .clk(N__94306),
            .ce(),
            .sr(N__43375));
    defparam \dron_frame_decoder_1.WDT_5_LC_8_18_5 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_5_LC_8_18_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_5_LC_8_18_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_5_LC_8_18_5  (
            .in0(_gnd_net_),
            .in1(N__43263),
            .in2(_gnd_net_),
            .in3(N__43186),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_5 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_4 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_5 ),
            .clk(N__94306),
            .ce(),
            .sr(N__43375));
    defparam \dron_frame_decoder_1.WDT_6_LC_8_18_6 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_6_LC_8_18_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_6_LC_8_18_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_6_LC_8_18_6  (
            .in0(_gnd_net_),
            .in1(N__43347),
            .in2(_gnd_net_),
            .in3(N__43183),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_6 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_5 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_6 ),
            .clk(N__94306),
            .ce(),
            .sr(N__43375));
    defparam \dron_frame_decoder_1.WDT_7_LC_8_18_7 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_7_LC_8_18_7 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_7_LC_8_18_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_7_LC_8_18_7  (
            .in0(_gnd_net_),
            .in1(N__43332),
            .in2(_gnd_net_),
            .in3(N__43180),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_7 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_6 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_7 ),
            .clk(N__94306),
            .ce(),
            .sr(N__43375));
    defparam \dron_frame_decoder_1.WDT_8_LC_8_19_0 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_8_LC_8_19_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_8_LC_8_19_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_8_LC_8_19_0  (
            .in0(_gnd_net_),
            .in1(N__43276),
            .in2(_gnd_net_),
            .in3(N__43177),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_8 ),
            .ltout(),
            .carryin(bfn_8_19_0_),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_8 ),
            .clk(N__94324),
            .ce(),
            .sr(N__43371));
    defparam \dron_frame_decoder_1.WDT_9_LC_8_19_1 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_9_LC_8_19_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_9_LC_8_19_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_9_LC_8_19_1  (
            .in0(_gnd_net_),
            .in1(N__43248),
            .in2(_gnd_net_),
            .in3(N__43174),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_9 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_8 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_9 ),
            .clk(N__94324),
            .ce(),
            .sr(N__43371));
    defparam \dron_frame_decoder_1.WDT_10_LC_8_19_2 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_10_LC_8_19_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_10_LC_8_19_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_10_LC_8_19_2  (
            .in0(_gnd_net_),
            .in1(N__43317),
            .in2(_gnd_net_),
            .in3(N__43171),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_10 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_9 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_10 ),
            .clk(N__94324),
            .ce(),
            .sr(N__43371));
    defparam \dron_frame_decoder_1.WDT_11_LC_8_19_3 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_11_LC_8_19_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_11_LC_8_19_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_11_LC_8_19_3  (
            .in0(_gnd_net_),
            .in1(N__43213),
            .in2(_gnd_net_),
            .in3(N__43168),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_11 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_10 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_11 ),
            .clk(N__94324),
            .ce(),
            .sr(N__43371));
    defparam \dron_frame_decoder_1.WDT_12_LC_8_19_4 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_12_LC_8_19_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_12_LC_8_19_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_12_LC_8_19_4  (
            .in0(_gnd_net_),
            .in1(N__43495),
            .in2(_gnd_net_),
            .in3(N__43387),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_12 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_11 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_12 ),
            .clk(N__94324),
            .ce(),
            .sr(N__43371));
    defparam \dron_frame_decoder_1.WDT_13_LC_8_19_5 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_13_LC_8_19_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_13_LC_8_19_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_13_LC_8_19_5  (
            .in0(_gnd_net_),
            .in1(N__43479),
            .in2(_gnd_net_),
            .in3(N__43384),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_13 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_12 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_13 ),
            .clk(N__94324),
            .ce(),
            .sr(N__43371));
    defparam \dron_frame_decoder_1.WDT_14_LC_8_19_6 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_14_LC_8_19_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_14_LC_8_19_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_14_LC_8_19_6  (
            .in0(_gnd_net_),
            .in1(N__43449),
            .in2(_gnd_net_),
            .in3(N__43381),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_14 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_13 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_14 ),
            .clk(N__94324),
            .ce(),
            .sr(N__43371));
    defparam \dron_frame_decoder_1.WDT_15_LC_8_19_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_15_LC_8_19_7 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_15_LC_8_19_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \dron_frame_decoder_1.WDT_15_LC_8_19_7  (
            .in0(_gnd_net_),
            .in1(N__43429),
            .in2(_gnd_net_),
            .in3(N__43378),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94324),
            .ce(),
            .sr(N__43371));
    defparam \dron_frame_decoder_1.WDT_RNI9TKF_6_LC_8_20_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNI9TKF_6_LC_8_20_0 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNI9TKF_6_LC_8_20_0 .LUT_INIT=16'b1110000011110000;
    LogicCell40 \dron_frame_decoder_1.WDT_RNI9TKF_6_LC_8_20_0  (
            .in0(N__43348),
            .in1(N__43333),
            .in2(N__43318),
            .in3(N__43219),
            .lcout(\dron_frame_decoder_1.WDT10lt12_0 ),
            .ltout(\dron_frame_decoder_1.WDT10lt12_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_RNIBUTU2_15_LC_8_20_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNIBUTU2_15_LC_8_20_1 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNIBUTU2_15_LC_8_20_1 .LUT_INIT=16'b0111111100110011;
    LogicCell40 \dron_frame_decoder_1.WDT_RNIBUTU2_15_LC_8_20_1  (
            .in0(N__43475),
            .in1(N__43427),
            .in2(N__43303),
            .in3(N__43282),
            .lcout(\dron_frame_decoder_1.WDT10_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_RNIA9RK1_11_LC_8_20_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNIA9RK1_11_LC_8_20_2 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNIA9RK1_11_LC_8_20_2 .LUT_INIT=16'b0000001100000111;
    LogicCell40 \dron_frame_decoder_1.WDT_RNIA9RK1_11_LC_8_20_2  (
            .in0(N__43211),
            .in1(N__43474),
            .in2(N__43450),
            .in3(N__43493),
            .lcout(\dron_frame_decoder_1.WDT10_0_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_RNIM3K1_4_LC_8_20_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNIM3K1_4_LC_8_20_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNIM3K1_4_LC_8_20_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \dron_frame_decoder_1.WDT_RNIM3K1_4_LC_8_20_3  (
            .in0(N__43275),
            .in1(N__43264),
            .in2(N__43249),
            .in3(N__43234),
            .lcout(\dron_frame_decoder_1.WDT10lto9_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_RNINA9N1_11_LC_8_20_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNINA9N1_11_LC_8_20_4 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNINA9N1_11_LC_8_20_4 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \dron_frame_decoder_1.WDT_RNINA9N1_11_LC_8_20_4  (
            .in0(N__43212),
            .in1(N__43494),
            .in2(N__43480),
            .in3(N__43456),
            .lcout(),
            .ltout(\dron_frame_decoder_1.WDT10lt14_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_RNIPI9R2_15_LC_8_20_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNIPI9R2_15_LC_8_20_5 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNIPI9R2_15_LC_8_20_5 .LUT_INIT=16'b0000000101010101;
    LogicCell40 \dron_frame_decoder_1.WDT_RNIPI9R2_15_LC_8_20_5  (
            .in0(N__48548),
            .in1(N__43448),
            .in2(N__43432),
            .in3(N__43428),
            .lcout(\dron_frame_decoder_1.N_218 ),
            .ltout(\dron_frame_decoder_1.N_218_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_2_LC_8_20_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_2_LC_8_20_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_2_LC_8_20_6 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \dron_frame_decoder_1.state_2_LC_8_20_6  (
            .in0(N__48550),
            .in1(N__46286),
            .in2(N__43414),
            .in3(N__43411),
            .lcout(\dron_frame_decoder_1.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94339),
            .ce(),
            .sr(N__86431));
    defparam \dron_frame_decoder_1.state_RNI7GSU_2_LC_8_20_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNI7GSU_2_LC_8_20_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNI7GSU_2_LC_8_20_7 .LUT_INIT=16'b1011101010101010;
    LogicCell40 \dron_frame_decoder_1.state_RNI7GSU_2_LC_8_20_7  (
            .in0(N__86602),
            .in1(N__43410),
            .in2(N__46288),
            .in3(N__48549),
            .lcout(\dron_frame_decoder_1.N_700_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_10_LC_8_21_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_10_LC_8_21_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_10_LC_8_21_5 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \Commands_frame_decoder.state_10_LC_8_21_5  (
            .in0(N__48254),
            .in1(N__45475),
            .in2(_gnd_net_),
            .in3(N__69417),
            .lcout(\Commands_frame_decoder.stateZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94354),
            .ce(),
            .sr(N__86422));
    defparam \Commands_frame_decoder.state_13_LC_8_21_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_13_LC_8_21_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_13_LC_8_21_7 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \Commands_frame_decoder.state_13_LC_8_21_7  (
            .in0(N__48617),
            .in1(N__48583),
            .in2(_gnd_net_),
            .in3(N__69418),
            .lcout(\Commands_frame_decoder.stateZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94354),
            .ce(),
            .sr(N__86422));
    defparam \ppm_encoder_1.init_pulses_RNIB3081_0_6_LC_9_1_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIB3081_0_6_LC_9_1_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIB3081_0_6_LC_9_1_0 .LUT_INIT=16'b0000111110000111;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIB3081_0_6_LC_9_1_0  (
            .in0(N__53693),
            .in1(N__43738),
            .in2(N__49137),
            .in3(N__52895),
            .lcout(),
            .ltout(\ppm_encoder_1.N_262_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNINSI75_6_LC_9_1_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNINSI75_6_LC_9_1_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNINSI75_6_LC_9_1_1 .LUT_INIT=16'b1111000011100001;
    LogicCell40 \ppm_encoder_1.init_pulses_RNINSI75_6_LC_9_1_1  (
            .in0(N__53550),
            .in1(N__49092),
            .in2(N__43393),
            .in3(N__44513),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_0_axb_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI20JF6_6_LC_9_1_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI20JF6_6_LC_9_1_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI20JF6_6_LC_9_1_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI20JF6_6_LC_9_1_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43390),
            .in3(N__43916),
            .lcout(\ppm_encoder_1.init_pulses_RNI20JF6Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIL06I1_6_LC_9_1_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIL06I1_6_LC_9_1_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIL06I1_6_LC_9_1_3 .LUT_INIT=16'b1100111000001010;
    LogicCell40 \ppm_encoder_1.elevator_RNIL06I1_6_LC_9_1_3  (
            .in0(N__43779),
            .in1(N__53692),
            .in2(N__47452),
            .in3(N__43746),
            .lcout(\ppm_encoder_1.N_306 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_6_LC_9_1_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_6_LC_9_1_4 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_6_LC_9_1_4 .LUT_INIT=16'b1010010111001100;
    LogicCell40 \ppm_encoder_1.elevator_6_LC_9_1_4  (
            .in0(N__47671),
            .in1(N__43780),
            .in2(N__54613),
            .in3(N__51378),
            .lcout(\ppm_encoder_1.elevatorZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94089),
            .ce(),
            .sr(N__86513));
    defparam \ppm_encoder_1.rudder_6_LC_9_1_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_6_LC_9_1_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.rudder_6_LC_9_1_5 .LUT_INIT=16'b0101111101010000;
    LogicCell40 \ppm_encoder_1.rudder_6_LC_9_1_5  (
            .in0(N__43771),
            .in1(_gnd_net_),
            .in2(N__51379),
            .in3(N__43747),
            .lcout(\ppm_encoder_1.rudderZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94089),
            .ce(),
            .sr(N__86513));
    defparam \ppm_encoder_1.init_pulses_RNIB3081_6_LC_9_1_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIB3081_6_LC_9_1_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIB3081_6_LC_9_1_6 .LUT_INIT=16'b1111000001111000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIB3081_6_LC_9_1_6  (
            .in0(N__53694),
            .in1(N__43737),
            .in2(N__49136),
            .in3(N__52894),
            .lcout(\ppm_encoder_1.N_262_i_i ),
            .ltout(\ppm_encoder_1.N_262_i_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIQOIP3_6_LC_9_1_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIQOIP3_6_LC_9_1_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIQOIP3_6_LC_9_1_7 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIQOIP3_6_LC_9_1_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43672),
            .in3(N__43669),
            .lcout(\ppm_encoder_1.init_pulses_RNIQOIP3Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIJ0D66_0_LC_9_2_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNIJ0D66_0_LC_9_2_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIJ0D66_0_LC_9_2_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIJ0D66_0_LC_9_2_0  (
            .in0(_gnd_net_),
            .in1(N__44233),
            .in2(N__44281),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_2_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_1_LC_9_2_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_1_LC_9_2_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_1_LC_9_2_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_1_LC_9_2_1  (
            .in0(_gnd_net_),
            .in1(N__43645),
            .in2(N__43633),
            .in3(N__43600),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_1 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_0 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_2_LC_9_2_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_2_LC_9_2_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_2_LC_9_2_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_2_LC_9_2_2  (
            .in0(_gnd_net_),
            .in1(N__43597),
            .in2(N__43585),
            .in3(N__43546),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_2 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_1 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_3_LC_9_2_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_3_LC_9_2_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_3_LC_9_2_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_3_LC_9_2_3  (
            .in0(_gnd_net_),
            .in1(N__43543),
            .in2(N__43531),
            .in3(N__43498),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_3 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_2 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_4_LC_9_2_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_4_LC_9_2_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_4_LC_9_2_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_4_LC_9_2_4  (
            .in0(_gnd_net_),
            .in1(N__44011),
            .in2(N__43996),
            .in3(N__43966),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_4 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_3 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_5_LC_9_2_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_5_LC_9_2_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_5_LC_9_2_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_5_LC_9_2_5  (
            .in0(_gnd_net_),
            .in1(N__43963),
            .in2(N__43954),
            .in3(N__43933),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_5 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_4 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_6_LC_9_2_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_6_LC_9_2_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_6_LC_9_2_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_6_LC_9_2_6  (
            .in0(_gnd_net_),
            .in1(N__43930),
            .in2(N__43923),
            .in3(N__43900),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_6 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_5 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_7_LC_9_2_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_7_LC_9_2_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_7_LC_9_2_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_7_LC_9_2_7  (
            .in0(_gnd_net_),
            .in1(N__44185),
            .in2(N__44149),
            .in3(N__43897),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_7 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_6 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_8_LC_9_3_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_8_LC_9_3_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_8_LC_9_3_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_8_LC_9_3_0  (
            .in0(_gnd_net_),
            .in1(N__43894),
            .in2(N__43882),
            .in3(N__43864),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_8 ),
            .ltout(),
            .carryin(bfn_9_3_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_9_LC_9_3_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_9_LC_9_3_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_9_LC_9_3_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_9_LC_9_3_1  (
            .in0(_gnd_net_),
            .in1(N__43861),
            .in2(N__43849),
            .in3(N__43825),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_9 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_8 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_10_LC_9_3_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_10_LC_9_3_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_10_LC_9_3_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_10_LC_9_3_2  (
            .in0(_gnd_net_),
            .in1(N__43822),
            .in2(N__43810),
            .in3(N__43786),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_10 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_9 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_11_LC_9_3_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_11_LC_9_3_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_11_LC_9_3_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_11_LC_9_3_3  (
            .in0(_gnd_net_),
            .in1(N__44197),
            .in2(N__44224),
            .in3(N__43783),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_11 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_10 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_12_LC_9_3_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_12_LC_9_3_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_12_LC_9_3_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_12_LC_9_3_4  (
            .in0(_gnd_net_),
            .in1(N__56083),
            .in2(N__56110),
            .in3(N__44131),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_12 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_11 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_13_LC_9_3_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_13_LC_9_3_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_13_LC_9_3_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_13_LC_9_3_5  (
            .in0(_gnd_net_),
            .in1(N__44128),
            .in2(N__44122),
            .in3(N__44086),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_13 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_12 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_14_LC_9_3_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_14_LC_9_3_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_14_LC_9_3_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_14_LC_9_3_6  (
            .in0(_gnd_net_),
            .in1(N__44410),
            .in2(N__44389),
            .in3(N__44077),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_14 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_13 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_15_LC_9_3_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_15_LC_9_3_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_15_LC_9_3_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_15_LC_9_3_7  (
            .in0(_gnd_net_),
            .in1(N__44074),
            .in2(N__44068),
            .in3(N__44053),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_15 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_14 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_16_LC_9_4_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_16_LC_9_4_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_16_LC_9_4_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_16_LC_9_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__46864),
            .in3(N__44044),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_16 ),
            .ltout(),
            .carryin(bfn_9_4_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_17_LC_9_4_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_17_LC_9_4_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_17_LC_9_4_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_17_LC_9_4_1  (
            .in0(_gnd_net_),
            .in1(N__44041),
            .in2(_gnd_net_),
            .in3(N__44023),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_17 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_16 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_18_LC_9_4_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNO_0_18_LC_9_4_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_18_LC_9_4_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_18_LC_9_4_2  (
            .in0(_gnd_net_),
            .in1(N__49004),
            .in2(_gnd_net_),
            .in3(N__44020),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIOLS41_11_LC_9_4_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIOLS41_11_LC_9_4_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIOLS41_11_LC_9_4_4 .LUT_INIT=16'b1111000001111000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIOLS41_11_LC_9_4_4  (
            .in0(N__53809),
            .in1(N__53679),
            .in2(N__46792),
            .in3(N__52890),
            .lcout(\ppm_encoder_1.N_266_i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_0_LC_9_4_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNO_1_0_LC_9_4_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_0_LC_9_4_5 .LUT_INIT=16'b1010101010011001;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_0_LC_9_4_5  (
            .in0(N__44256),
            .in1(N__44344),
            .in2(_gnd_net_),
            .in3(N__47521),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNI0EA05_0_LC_9_4_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNI0EA05_0_LC_9_4_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNI0EA05_0_LC_9_4_6 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \ppm_encoder_1.throttle_RNI0EA05_0_LC_9_4_6  (
            .in0(N__44304),
            .in1(N__44292),
            .in2(N__44279),
            .in3(N__44502),
            .lcout(\ppm_encoder_1.throttle_RNI0EA05Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIU1F76_11_LC_9_4_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIU1F76_11_LC_9_4_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIU1F76_11_LC_9_4_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIU1F76_11_LC_9_4_7  (
            .in0(_gnd_net_),
            .in1(N__44220),
            .in2(_gnd_net_),
            .in3(N__44209),
            .lcout(\ppm_encoder_1.init_pulses_RNIU1F76Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNID4081_0_7_LC_9_5_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNID4081_0_7_LC_9_5_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNID4081_0_7_LC_9_5_0 .LUT_INIT=16'b0000111110000111;
    LogicCell40 \ppm_encoder_1.init_pulses_RNID4081_0_7_LC_9_5_0  (
            .in0(N__53796),
            .in1(N__53639),
            .in2(N__49071),
            .in3(N__52886),
            .lcout(),
            .ltout(\ppm_encoder_1.N_263_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIF99E5_7_LC_9_5_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIF99E5_7_LC_9_5_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIF99E5_7_LC_9_5_1 .LUT_INIT=16'b0000111100011110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIF99E5_7_LC_9_5_1  (
            .in0(N__44176),
            .in1(N__49035),
            .in2(N__44191),
            .in3(N__44510),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_0_axb_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNISD9M6_7_LC_9_5_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNISD9M6_7_LC_9_5_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNISD9M6_7_LC_9_5_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNISD9M6_7_LC_9_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__44188),
            .in3(N__44142),
            .lcout(\ppm_encoder_1.init_pulses_RNISD9M6Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIPQ8E1_7_LC_9_5_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIPQ8E1_7_LC_9_5_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIPQ8E1_7_LC_9_5_3 .LUT_INIT=16'b0101110100001100;
    LogicCell40 \ppm_encoder_1.throttle_RNIPQ8E1_7_LC_9_5_3  (
            .in0(N__54287),
            .in1(N__44680),
            .in2(N__54319),
            .in3(N__44594),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_0_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIN26I1_7_LC_9_5_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIN26I1_7_LC_9_5_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIN26I1_7_LC_9_5_4 .LUT_INIT=16'b0000110001011101;
    LogicCell40 \ppm_encoder_1.elevator_RNIN26I1_7_LC_9_5_4  (
            .in0(N__50284),
            .in1(N__53638),
            .in2(N__44170),
            .in3(N__47438),
            .lcout(\ppm_encoder_1.N_310 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNID4081_7_LC_9_5_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNID4081_7_LC_9_5_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNID4081_7_LC_9_5_5 .LUT_INIT=16'b1001110011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNID4081_7_LC_9_5_5  (
            .in0(N__52885),
            .in1(N__49064),
            .in2(N__53680),
            .in3(N__53795),
            .lcout(\ppm_encoder_1.N_263_i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNI4FET_1_LC_9_5_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNI4FET_1_LC_9_5_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNI4FET_1_LC_9_5_6 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_RNI4FET_1_LC_9_5_6  (
            .in0(N__53797),
            .in1(N__54238),
            .in2(_gnd_net_),
            .in3(N__54078),
            .lcout(\ppm_encoder_1.N_293 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_esr_RNI7CAL1_14_LC_9_6_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_RNI7CAL1_14_LC_9_6_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.aileron_esr_RNI7CAL1_14_LC_9_6_0 .LUT_INIT=16'b0101110100001100;
    LogicCell40 \ppm_encoder_1.aileron_esr_RNI7CAL1_14_LC_9_6_0  (
            .in0(N__53907),
            .in1(N__44686),
            .in2(N__53886),
            .in3(N__44608),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_i_i_0_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNISK6K5_14_LC_9_6_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNISK6K5_14_LC_9_6_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNISK6K5_14_LC_9_6_1 .LUT_INIT=16'b0011001100110110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNISK6K5_14_LC_9_6_1  (
            .in0(N__48726),
            .in1(N__44350),
            .in2(N__44521),
            .in3(N__44511),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_0_axb_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIP98N6_14_LC_9_6_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIP98N6_14_LC_9_6_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIP98N6_14_LC_9_6_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIP98N6_14_LC_9_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__44413),
            .in3(N__44382),
            .lcout(\ppm_encoder_1.init_pulses_RNIP98N6Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_esr_RNI6C0M1_14_LC_9_6_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_esr_RNI6C0M1_14_LC_9_6_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_esr_RNI6C0M1_14_LC_9_6_3 .LUT_INIT=16'b0000010111001101;
    LogicCell40 \ppm_encoder_1.elevator_esr_RNI6C0M1_14_LC_9_6_3  (
            .in0(N__47566),
            .in1(N__56215),
            .in2(N__47451),
            .in3(N__44401),
            .lcout(\ppm_encoder_1.N_309 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNITK131_14_LC_9_6_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNITK131_14_LC_9_6_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNITK131_14_LC_9_6_4 .LUT_INIT=16'b1001110011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNITK131_14_LC_9_6_4  (
            .in0(N__52889),
            .in1(N__48763),
            .in2(N__56251),
            .in3(N__49658),
            .lcout(\ppm_encoder_1.N_269_i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_11_LC_9_6_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_11_LC_9_6_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_11_LC_9_6_5 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_11_LC_9_6_5  (
            .in0(N__46796),
            .in1(N__44371),
            .in2(N__44362),
            .in3(N__50920),
            .lcout(\ppm_encoder_1.pulses2count_9_0_3_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNITK131_1_14_LC_9_6_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNITK131_1_14_LC_9_6_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNITK131_1_14_LC_9_6_7 .LUT_INIT=16'b0010110100001111;
    LogicCell40 \ppm_encoder_1.init_pulses_RNITK131_1_14_LC_9_6_7  (
            .in0(N__49657),
            .in1(N__52888),
            .in2(N__48770),
            .in3(N__56216),
            .lcout(\ppm_encoder_1.N_269_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_LC_9_7_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_LC_9_7_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_LC_9_7_1 .LUT_INIT=16'b0000101100000001;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_2_LC_9_7_1  (
            .in0(N__52900),
            .in1(N__47129),
            .in2(N__71061),
            .in3(N__56242),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94134),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNI5HI71_6_LC_9_7_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNI5HI71_6_LC_9_7_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNI5HI71_6_LC_9_7_2 .LUT_INIT=16'b0011000010001000;
    LogicCell40 \ppm_encoder_1.throttle_RNI5HI71_6_LC_9_7_2  (
            .in0(N__44956),
            .in1(N__54047),
            .in2(N__44941),
            .in3(N__44921),
            .lcout(\ppm_encoder_1.un2_throttle_0_2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNI1I491_12_LC_9_7_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNI1I491_12_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNI1I491_12_LC_9_7_3 .LUT_INIT=16'b0001000100011111;
    LogicCell40 \ppm_encoder_1.throttle_RNI1I491_12_LC_9_7_3  (
            .in0(N__54048),
            .in1(N__47721),
            .in2(N__50696),
            .in3(N__54162),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_axb_12_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_LC_9_7_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_LC_9_7_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_LC_9_7_4 .LUT_INIT=16'b1110111011111100;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_0_LC_9_7_4  (
            .in0(N__54164),
            .in1(N__71040),
            .in2(N__47186),
            .in3(N__52901),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94134),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_3_LC_9_7_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_3_LC_9_7_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_3_LC_9_7_5 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_3_LC_9_7_5  (
            .in0(N__50934),
            .in1(N__47296),
            .in2(_gnd_net_),
            .in3(N__44866),
            .lcout(\ppm_encoder_1.pulses2count_9_0_0_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_LC_9_7_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_LC_9_7_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_LC_9_7_6 .LUT_INIT=16'b0000000011000110;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_1_LC_9_7_6  (
            .in0(N__54165),
            .in1(N__54050),
            .in2(N__52906),
            .in3(N__71044),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94134),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_9_LC_9_7_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_9_LC_9_7_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_9_LC_9_7_7 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_9_LC_9_7_7  (
            .in0(N__54049),
            .in1(N__54163),
            .in2(_gnd_net_),
            .in3(N__44982),
            .lcout(\ppm_encoder_1.N_425 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_8_LC_9_8_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_8_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_8_LC_9_8_0 .LUT_INIT=16'b0000110001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_8_LC_9_8_0  (
            .in0(N__44818),
            .in1(N__54076),
            .in2(N__44788),
            .in3(N__54193),
            .lcout(\ppm_encoder_1.pulses2count_9_i_1_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_9_LC_9_8_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_9_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_9_LC_9_8_3 .LUT_INIT=16'b0010000000101010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_9_LC_9_8_3  (
            .in0(N__54077),
            .in1(N__44708),
            .in2(N__54227),
            .in3(N__44753),
            .lcout(\ppm_encoder_1.pulses2count_9_i_1_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_9_LC_9_8_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_9_LC_9_8_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_9_LC_9_8_4 .LUT_INIT=16'b0010111011100010;
    LogicCell40 \ppm_encoder_1.elevator_9_LC_9_8_4  (
            .in0(N__44709),
            .in1(N__51267),
            .in2(N__54514),
            .in3(N__47635),
            .lcout(\ppm_encoder_1.elevatorZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94140),
            .ce(),
            .sr(N__86488));
    defparam \ppm_encoder_1.aileron_7_LC_9_8_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_7_LC_9_8_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_7_LC_9_8_6 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.aileron_7_LC_9_8_6  (
            .in0(N__47803),
            .in1(N__54415),
            .in2(N__54289),
            .in3(N__51271),
            .lcout(\ppm_encoder_1.aileronZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94140),
            .ce(),
            .sr(N__86488));
    defparam \ppm_encoder_1.throttle_7_LC_9_8_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_7_LC_9_8_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_7_LC_9_8_7 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.throttle_7_LC_9_8_7  (
            .in0(N__45151),
            .in1(N__45136),
            .in2(N__51350),
            .in3(N__54311),
            .lcout(\ppm_encoder_1.throttleZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94140),
            .ce(),
            .sr(N__86488));
    defparam \ppm_encoder_1.throttle_8_LC_9_9_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_8_LC_9_9_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_8_LC_9_9_0 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.throttle_8_LC_9_9_0  (
            .in0(N__45106),
            .in1(N__45076),
            .in2(N__45059),
            .in3(N__51278),
            .lcout(\ppm_encoder_1.throttleZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94153),
            .ce(),
            .sr(N__86481));
    defparam \ppm_encoder_1.throttle_9_LC_9_9_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_9_LC_9_9_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_9_LC_9_9_1 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.throttle_9_LC_9_9_1  (
            .in0(N__45028),
            .in1(N__45001),
            .in2(N__51352),
            .in3(N__44978),
            .lcout(\ppm_encoder_1.throttleZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94153),
            .ce(),
            .sr(N__86481));
    defparam \ppm_encoder_1.aileron_6_LC_9_9_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_6_LC_9_9_3 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_6_LC_9_9_3 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \ppm_encoder_1.aileron_6_LC_9_9_3  (
            .in0(N__47812),
            .in1(N__54447),
            .in2(N__51351),
            .in3(N__44955),
            .lcout(\ppm_encoder_1.aileronZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94153),
            .ce(),
            .sr(N__86481));
    defparam \uart_drone.bit_Count_0_LC_9_9_4 .C_ON=1'b0;
    defparam \uart_drone.bit_Count_0_LC_9_9_4 .SEQ_MODE=4'b1000;
    defparam \uart_drone.bit_Count_0_LC_9_9_4 .LUT_INIT=16'b0000001011001100;
    LogicCell40 \uart_drone.bit_Count_0_LC_9_9_4  (
            .in0(N__53986),
            .in1(N__56606),
            .in2(N__56770),
            .in3(N__51468),
            .lcout(\uart_drone.bit_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94153),
            .ce(),
            .sr(N__86481));
    defparam \uart_drone.bit_Count_1_LC_9_9_5 .C_ON=1'b0;
    defparam \uart_drone.bit_Count_1_LC_9_9_5 .SEQ_MODE=4'b1000;
    defparam \uart_drone.bit_Count_1_LC_9_9_5 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \uart_drone.bit_Count_1_LC_9_9_5  (
            .in0(N__51469),
            .in1(N__56539),
            .in2(N__56620),
            .in3(N__47739),
            .lcout(\uart_drone.bit_CountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94153),
            .ce(),
            .sr(N__86481));
    defparam \uart_drone.bit_Count_2_LC_9_9_6 .C_ON=1'b0;
    defparam \uart_drone.bit_Count_2_LC_9_9_6 .SEQ_MODE=4'b1000;
    defparam \uart_drone.bit_Count_2_LC_9_9_6 .LUT_INIT=16'b0001010001000100;
    LogicCell40 \uart_drone.bit_Count_2_LC_9_9_6  (
            .in0(N__47740),
            .in1(N__56478),
            .in2(N__56554),
            .in3(N__47731),
            .lcout(\uart_drone.bit_CountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94153),
            .ce(),
            .sr(N__86481));
    defparam \scaler_4.source_data_1_4_LC_9_10_0 .C_ON=1'b0;
    defparam \scaler_4.source_data_1_4_LC_9_10_0 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_4_LC_9_10_0 .LUT_INIT=16'b0111001011011000;
    LogicCell40 \scaler_4.source_data_1_4_LC_9_10_0  (
            .in0(N__48108),
            .in1(N__45182),
            .in2(N__47046),
            .in3(N__45237),
            .lcout(scaler_4_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94164),
            .ce(),
            .sr(N__86471));
    defparam \ppm_encoder_1.aileron_4_LC_9_10_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_4_LC_9_10_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_4_LC_9_10_6 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.aileron_4_LC_9_10_6  (
            .in0(N__47839),
            .in1(N__59332),
            .in2(N__46739),
            .in3(N__51259),
            .lcout(\ppm_encoder_1.aileronZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94164),
            .ce(),
            .sr(N__86471));
    defparam \uart_drone.timer_Count_RNI9E9J_2_LC_9_11_2 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNI9E9J_2_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNI9E9J_2_LC_9_11_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_drone.timer_Count_RNI9E9J_2_LC_9_11_2  (
            .in0(_gnd_net_),
            .in1(N__47885),
            .in2(_gnd_net_),
            .in3(N__51497),
            .lcout(\uart_drone.N_126_li ),
            .ltout(\uart_drone.N_126_li_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNIAT1D1_4_LC_9_11_3 .C_ON=1'b0;
    defparam \uart_drone.state_RNIAT1D1_4_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNIAT1D1_4_LC_9_11_3 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \uart_drone.state_RNIAT1D1_4_LC_9_11_3  (
            .in0(N__54823),
            .in1(N__54756),
            .in2(N__45274),
            .in3(N__70918),
            .lcout(\uart_drone.N_143 ),
            .ltout(\uart_drone.N_143_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_2_LC_9_11_4 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_2_LC_9_11_4 .SEQ_MODE=4'b1000;
    defparam \uart_drone.timer_Count_2_LC_9_11_4 .LUT_INIT=16'b0011001000000000;
    LogicCell40 \uart_drone.timer_Count_2_LC_9_11_4  (
            .in0(N__51563),
            .in1(N__70929),
            .in2(N__45271),
            .in3(N__47869),
            .lcout(\uart_drone.timer_CountZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94177),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNIDGR31_2_LC_9_11_5 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNIDGR31_2_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNIDGR31_2_LC_9_11_5 .LUT_INIT=16'b1100110010000000;
    LogicCell40 \uart_drone.timer_Count_RNIDGR31_2_LC_9_11_5  (
            .in0(N__51496),
            .in1(N__54822),
            .in2(N__47887),
            .in3(N__54755),
            .lcout(\uart_drone.data_rdyc_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un2_source_data_0_cry_1_c_RNO_LC_9_11_7 .C_ON=1'b0;
    defparam \scaler_4.un2_source_data_0_cry_1_c_RNO_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un2_source_data_0_cry_1_c_RNO_LC_9_11_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \scaler_4.un2_source_data_0_cry_1_c_RNO_LC_9_11_7  (
            .in0(N__45181),
            .in1(N__45266),
            .in2(_gnd_net_),
            .in3(N__45236),
            .lcout(\scaler_4.un2_source_data_0_cry_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_0_LC_9_12_1 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_0_LC_9_12_1 .SEQ_MODE=4'b1000;
    defparam \uart_drone.timer_Count_0_LC_9_12_1 .LUT_INIT=16'b0000000000110010;
    LogicCell40 \uart_drone.timer_Count_0_LC_9_12_1  (
            .in0(N__50778),
            .in1(N__47912),
            .in2(N__51568),
            .in3(N__70839),
            .lcout(\uart_drone.timer_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94191),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.state_RNICP2N1_0_LC_9_12_3 .C_ON=1'b0;
    defparam \pid_alt.state_RNICP2N1_0_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.state_RNICP2N1_0_LC_9_12_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pid_alt.state_RNICP2N1_0_LC_9_12_3  (
            .in0(_gnd_net_),
            .in1(N__46417),
            .in2(_gnd_net_),
            .in3(N__93122),
            .lcout(\pid_alt.N_933_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_offset4data_esr_0_LC_9_13_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_0_LC_9_13_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_0_LC_9_13_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_0_LC_9_13_0  (
            .in0(N__88260),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(frame_decoder_OFF4data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94206),
            .ce(N__45460),
            .sr(N__86455));
    defparam \Commands_frame_decoder.source_offset4data_esr_1_LC_9_13_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_1_LC_9_13_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_1_LC_9_13_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_1_LC_9_13_1  (
            .in0(N__85468),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(frame_decoder_OFF4data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94206),
            .ce(N__45460),
            .sr(N__86455));
    defparam \Commands_frame_decoder.source_offset4data_esr_2_LC_9_13_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_2_LC_9_13_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_2_LC_9_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_2_LC_9_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__92494),
            .lcout(frame_decoder_OFF4data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94206),
            .ce(N__45460),
            .sr(N__86455));
    defparam \Commands_frame_decoder.source_offset4data_esr_3_LC_9_13_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_3_LC_9_13_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_3_LC_9_13_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_3_LC_9_13_3  (
            .in0(N__92301),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(frame_decoder_OFF4data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94206),
            .ce(N__45460),
            .sr(N__86455));
    defparam \Commands_frame_decoder.source_offset4data_esr_4_LC_9_13_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_4_LC_9_13_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_4_LC_9_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_4_LC_9_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88847),
            .lcout(frame_decoder_OFF4data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94206),
            .ce(N__45460),
            .sr(N__86455));
    defparam \Commands_frame_decoder.source_offset4data_esr_5_LC_9_13_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_5_LC_9_13_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_5_LC_9_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_5_LC_9_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88663),
            .lcout(frame_decoder_OFF4data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94206),
            .ce(N__45460),
            .sr(N__86455));
    defparam \Commands_frame_decoder.source_offset4data_esr_6_LC_9_13_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_6_LC_9_13_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_6_LC_9_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_6_LC_9_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88505),
            .lcout(frame_decoder_OFF4data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94206),
            .ce(N__45460),
            .sr(N__86455));
    defparam \Commands_frame_decoder.source_offset4data_ess_7_LC_9_13_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_ess_7_LC_9_13_7 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_offset4data_ess_7_LC_9_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_ess_7_LC_9_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__92071),
            .lcout(frame_decoder_OFF4data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94206),
            .ce(N__45460),
            .sr(N__86455));
    defparam \Commands_frame_decoder.source_xy_kp_e_0_0_LC_9_14_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_0_LC_9_14_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_0_LC_9_14_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \Commands_frame_decoder.source_xy_kp_e_0_0_LC_9_14_0  (
            .in0(N__88254),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__93143),
            .lcout(xy_kp_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94223),
            .ce(N__48031),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kp_e_0_1_LC_9_14_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_1_LC_9_14_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_1_LC_9_14_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_kp_e_0_1_LC_9_14_1  (
            .in0(N__93144),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85464),
            .lcout(xy_kp_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94223),
            .ce(N__48031),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kp_e_0_2_LC_9_14_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_2_LC_9_14_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_2_LC_9_14_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_xy_kp_e_0_2_LC_9_14_2  (
            .in0(_gnd_net_),
            .in1(N__92465),
            .in2(_gnd_net_),
            .in3(N__93145),
            .lcout(xy_kp_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94223),
            .ce(N__48031),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kp_e_0_3_LC_9_14_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_3_LC_9_14_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_3_LC_9_14_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_kp_e_0_3_LC_9_14_3  (
            .in0(N__93146),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__92279),
            .lcout(xy_kp_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94223),
            .ce(N__48031),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kp_0_e_0_4_LC_9_14_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kp_0_e_0_4_LC_9_14_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kp_0_e_0_4_LC_9_14_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_xy_kp_0_e_0_4_LC_9_14_4  (
            .in0(_gnd_net_),
            .in1(N__88636),
            .in2(_gnd_net_),
            .in3(N__93142),
            .lcout(xy_kp_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94223),
            .ce(N__48031),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kp_e_0_5_LC_9_14_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_5_LC_9_14_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_5_LC_9_14_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_kp_e_0_5_LC_9_14_5  (
            .in0(N__93147),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88489),
            .lcout(xy_kp_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94223),
            .ce(N__48031),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kp_e_0_6_LC_9_14_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_6_LC_9_14_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_6_LC_9_14_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_xy_kp_e_0_6_LC_9_14_6  (
            .in0(_gnd_net_),
            .in1(N__92070),
            .in2(_gnd_net_),
            .in3(N__93148),
            .lcout(xy_kp_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94223),
            .ce(N__48031),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_7_LC_9_15_0 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_7_LC_9_15_0 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_7_LC_9_15_0 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \uart_pc.data_Aux_7_LC_9_15_0  (
            .in0(N__52237),
            .in1(N__45537),
            .in2(N__45516),
            .in3(N__46077),
            .lcout(\uart_pc.data_AuxZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94240),
            .ce(),
            .sr(N__46021));
    defparam \Commands_frame_decoder.state_RNIL23J_2_LC_9_15_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIL23J_2_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIL23J_2_LC_9_15_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Commands_frame_decoder.state_RNIL23J_2_LC_9_15_1  (
            .in0(_gnd_net_),
            .in1(N__52464),
            .in2(_gnd_net_),
            .in3(N__86589),
            .lcout(\Commands_frame_decoder.un1_sink_data_valid_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNILP1J_9_LC_9_15_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNILP1J_9_LC_9_15_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNILP1J_9_LC_9_15_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_RNILP1J_9_LC_9_15_2  (
            .in0(_gnd_net_),
            .in1(N__48216),
            .in2(_gnd_net_),
            .in3(N__55258),
            .lcout(\Commands_frame_decoder.source_offset4data_1_sqmuxa ),
            .ltout(\Commands_frame_decoder.source_offset4data_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIS93J_9_LC_9_15_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIS93J_9_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIS93J_9_LC_9_15_3 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \Commands_frame_decoder.state_RNIS93J_9_LC_9_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__45463),
            .in3(N__86593),
            .lcout(\Commands_frame_decoder.source_offset4data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIM33J_3_LC_9_15_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIM33J_3_LC_9_15_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIM33J_3_LC_9_15_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \Commands_frame_decoder.state_RNIM33J_3_LC_9_15_4  (
            .in0(N__86590),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52401),
            .lcout(\Commands_frame_decoder.source_CH2data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIN43J_4_LC_9_15_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIN43J_4_LC_9_15_5 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIN43J_4_LC_9_15_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Commands_frame_decoder.state_RNIN43J_4_LC_9_15_5  (
            .in0(_gnd_net_),
            .in1(N__69441),
            .in2(_gnd_net_),
            .in3(N__86591),
            .lcout(\Commands_frame_decoder.source_CH3data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIO53J_5_LC_9_15_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIO53J_5_LC_9_15_6 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIO53J_5_LC_9_15_6 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \Commands_frame_decoder.state_RNIO53J_5_LC_9_15_6  (
            .in0(N__86592),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51940),
            .lcout(\Commands_frame_decoder.source_CH4data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNID98K_4_LC_9_15_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNID98K_4_LC_9_15_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNID98K_4_LC_9_15_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \dron_frame_decoder_1.state_RNID98K_4_LC_9_15_7  (
            .in0(_gnd_net_),
            .in1(N__69315),
            .in2(_gnd_net_),
            .in3(N__86594),
            .lcout(\dron_frame_decoder_1.N_724_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIBLRB2_4_LC_9_16_0 .C_ON=1'b0;
    defparam \uart_pc.state_RNIBLRB2_4_LC_9_16_0 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIBLRB2_4_LC_9_16_0 .LUT_INIT=16'b1101111111001100;
    LogicCell40 \uart_pc.state_RNIBLRB2_4_LC_9_16_0  (
            .in0(N__45874),
            .in1(N__45855),
            .in2(N__45811),
            .in3(N__45795),
            .lcout(\uart_pc.un1_state_2_0 ),
            .ltout(\uart_pc.un1_state_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_0_LC_9_16_1 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_0_LC_9_16_1 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_0_LC_9_16_1 .LUT_INIT=16'b1100101011001100;
    LogicCell40 \uart_pc.data_Aux_0_LC_9_16_1  (
            .in0(N__52206),
            .in1(N__45945),
            .in2(N__45748),
            .in3(N__45745),
            .lcout(\uart_pc.data_AuxZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94257),
            .ce(),
            .sr(N__46017));
    defparam \uart_pc.data_Aux_1_LC_9_16_2 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_1_LC_9_16_2 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_1_LC_9_16_2 .LUT_INIT=16'b1010110010101010;
    LogicCell40 \uart_pc.data_Aux_1_LC_9_16_2  (
            .in0(N__46242),
            .in1(N__52207),
            .in2(N__46078),
            .in3(N__45739),
            .lcout(\uart_pc.data_AuxZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94257),
            .ce(),
            .sr(N__46017));
    defparam \uart_pc.data_Aux_2_LC_9_16_3 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_2_LC_9_16_3 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_2_LC_9_16_3 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \uart_pc.data_Aux_2_LC_9_16_3  (
            .in0(N__45733),
            .in1(N__46069),
            .in2(N__52234),
            .in3(N__45999),
            .lcout(\uart_pc.data_AuxZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94257),
            .ce(),
            .sr(N__46017));
    defparam \uart_pc.data_Aux_3_LC_9_16_4 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_3_LC_9_16_4 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_3_LC_9_16_4 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_pc.data_Aux_3_LC_9_16_4  (
            .in0(N__45727),
            .in1(N__52208),
            .in2(N__45721),
            .in3(N__46075),
            .lcout(\uart_pc.data_AuxZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94257),
            .ce(),
            .sr(N__46017));
    defparam \uart_pc.data_Aux_4_LC_9_16_5 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_4_LC_9_16_5 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_4_LC_9_16_5 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \uart_pc.data_Aux_4_LC_9_16_5  (
            .in0(N__46073),
            .in1(N__45696),
            .in2(N__52235),
            .in3(N__45703),
            .lcout(\uart_pc.data_AuxZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94257),
            .ce(),
            .sr(N__46017));
    defparam \uart_pc.data_Aux_5_LC_9_16_6 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_5_LC_9_16_6 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_5_LC_9_16_6 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_pc.data_Aux_5_LC_9_16_6  (
            .in0(N__46084),
            .in1(N__52209),
            .in2(N__45934),
            .in3(N__46076),
            .lcout(\uart_pc.data_AuxZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94257),
            .ce(),
            .sr(N__46017));
    defparam \uart_pc.data_Aux_6_LC_9_16_7 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_6_LC_9_16_7 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_6_LC_9_16_7 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \uart_pc.data_Aux_6_LC_9_16_7  (
            .in0(N__46074),
            .in1(N__46032),
            .in2(N__52236),
            .in3(N__46045),
            .lcout(\uart_pc.data_AuxZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94257),
            .ce(),
            .sr(N__46017));
    defparam \uart_pc.data_2_LC_9_17_0 .C_ON=1'b0;
    defparam \uart_pc.data_2_LC_9_17_0 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_2_LC_9_17_0 .LUT_INIT=16'b0000110010101010;
    LogicCell40 \uart_pc.data_2_LC_9_17_0  (
            .in0(N__92392),
            .in1(N__46000),
            .in2(N__45919),
            .in3(N__46270),
            .lcout(uart_pc_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94276),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_ns_0_a3_0_1_2_LC_9_17_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_ns_0_a3_0_1_2_LC_9_17_1 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_ns_0_a3_0_1_2_LC_9_17_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Commands_frame_decoder.state_ns_0_a3_0_1_2_LC_9_17_1  (
            .in0(_gnd_net_),
            .in1(N__92391),
            .in2(_gnd_net_),
            .in3(N__88574),
            .lcout(),
            .ltout(\Commands_frame_decoder.state_ns_0_a3_0_1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNITVPE1_1_LC_9_17_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNITVPE1_1_LC_9_17_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNITVPE1_1_LC_9_17_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Commands_frame_decoder.state_RNITVPE1_1_LC_9_17_2  (
            .in0(N__92041),
            .in1(N__88194),
            .in2(N__45988),
            .in3(N__45985),
            .lcout(\Commands_frame_decoder.N_406 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNO_0_1_LC_9_17_3 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNO_0_1_LC_9_17_3 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNO_0_1_LC_9_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_drone.timer_Count_RNO_0_1_LC_9_17_3  (
            .in0(_gnd_net_),
            .in1(N__47914),
            .in2(_gnd_net_),
            .in3(N__51025),
            .lcout(\uart_drone.timer_Count_RNO_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_0_LC_9_17_4 .C_ON=1'b0;
    defparam \uart_pc.data_0_LC_9_17_4 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_0_LC_9_17_4 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \uart_pc.data_0_LC_9_17_4  (
            .in0(N__45912),
            .in1(N__45946),
            .in2(N__88255),
            .in3(N__46268),
            .lcout(uart_pc_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94276),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_1_4_LC_9_17_5 .C_ON=1'b0;
    defparam \uart_pc.data_1_4_LC_9_17_5 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_1_4_LC_9_17_5 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \uart_pc.data_1_4_LC_9_17_5  (
            .in0(N__46267),
            .in1(N__45913),
            .in2(N__88640),
            .in3(N__45933),
            .lcout(uart_pc_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94276),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_1_LC_9_17_6 .C_ON=1'b0;
    defparam \uart_pc.data_1_LC_9_17_6 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_1_LC_9_17_6 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \uart_pc.data_1_LC_9_17_6  (
            .in0(N__45914),
            .in1(N__46269),
            .in2(N__46246),
            .in3(N__85445),
            .lcout(uart_pc_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94276),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_0_c_inv_LC_9_17_7 .C_ON=1'b0;
    defparam \pid_alt.error_cry_0_c_inv_LC_9_17_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_0_c_inv_LC_9_17_7 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pid_alt.error_cry_0_c_inv_LC_9_17_7  (
            .in0(N__65784),
            .in1(N__48371),
            .in2(_gnd_net_),
            .in3(N__46224),
            .lcout(\pid_alt.drone_altitude_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_13_LC_9_18_0 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_13_LC_9_18_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_13_LC_9_18_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \pid_side.error_i_acumm_13_LC_9_18_0  (
            .in0(_gnd_net_),
            .in1(N__62797),
            .in2(_gnd_net_),
            .in3(N__60454),
            .lcout(\pid_side.error_i_acummZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94292),
            .ce(N__60548),
            .sr(_gnd_net_));
    defparam \scaler_4.N_2928_i_l_ofx_LC_9_18_2 .C_ON=1'b0;
    defparam \scaler_4.N_2928_i_l_ofx_LC_9_18_2 .SEQ_MODE=4'b0000;
    defparam \scaler_4.N_2928_i_l_ofx_LC_9_18_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \scaler_4.N_2928_i_l_ofx_LC_9_18_2  (
            .in0(_gnd_net_),
            .in1(N__46210),
            .in2(_gnd_net_),
            .in3(N__46195),
            .lcout(\scaler_4.N_2928_i_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIHIDC_4_LC_9_18_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIHIDC_4_LC_9_18_4 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIHIDC_4_LC_9_18_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNIHIDC_4_LC_9_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48352),
            .lcout(drone_altitude_i_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIIJDC_5_LC_9_18_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIIJDC_5_LC_9_18_5 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIIJDC_5_LC_9_18_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNIIJDC_5_LC_9_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48490),
            .lcout(drone_altitude_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIJKDC_6_LC_9_18_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIJKDC_6_LC_9_18_6 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIJKDC_6_LC_9_18_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNIJKDC_6_LC_9_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48484),
            .lcout(drone_altitude_i_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIKLDC_7_LC_9_18_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIKLDC_7_LC_9_18_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIKLDC_7_LC_9_18_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNIKLDC_7_LC_9_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48478),
            .lcout(drone_altitude_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kd_1_LC_9_19_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kd_1_LC_9_19_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kd_1_LC_9_19_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_xy_kd_1_LC_9_19_1  (
            .in0(_gnd_net_),
            .in1(N__85457),
            .in2(_gnd_net_),
            .in3(N__93150),
            .lcout(xy_kd_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94307),
            .ce(N__91928),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIMNDC_9_LC_9_19_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIMNDC_9_LC_9_19_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIMNDC_9_LC_9_19_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNIMNDC_9_LC_9_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48715),
            .lcout(drone_altitude_i_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNI3T3K1_7_LC_9_20_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNI3T3K1_7_LC_9_20_0 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNI3T3K1_7_LC_9_20_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \dron_frame_decoder_1.state_RNI3T3K1_7_LC_9_20_0  (
            .in0(N__46329),
            .in1(N__46440),
            .in2(N__69246),
            .in3(N__46348),
            .lcout(\dron_frame_decoder_1.state_RNI3T3K1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_4_LC_9_20_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_4_LC_9_20_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_4_LC_9_20_2 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \dron_frame_decoder_1.state_4_LC_9_20_2  (
            .in0(N__46305),
            .in1(N__46334),
            .in2(N__48559),
            .in3(N__69272),
            .lcout(\dron_frame_decoder_1.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94325),
            .ce(),
            .sr(N__86423));
    defparam \dron_frame_decoder_1.state_5_LC_9_20_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_5_LC_9_20_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_5_LC_9_20_3 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \dron_frame_decoder_1.state_5_LC_9_20_3  (
            .in0(N__69273),
            .in1(N__46366),
            .in2(_gnd_net_),
            .in3(N__46306),
            .lcout(\dron_frame_decoder_1.stateZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94325),
            .ce(),
            .sr(N__86423));
    defparam \uart_drone.data_rdy_LC_9_20_4 .C_ON=1'b0;
    defparam \uart_drone.data_rdy_LC_9_20_4 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_rdy_LC_9_20_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_drone.data_rdy_LC_9_20_4  (
            .in0(_gnd_net_),
            .in1(N__56877),
            .in2(_gnd_net_),
            .in3(N__48205),
            .lcout(uart_drone_data_rdy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94325),
            .ce(),
            .sr(N__86423));
    defparam \dron_frame_decoder_1.state_RNI7Q6K_5_LC_9_20_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNI7Q6K_5_LC_9_20_5 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNI7Q6K_5_LC_9_20_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \dron_frame_decoder_1.state_RNI7Q6K_5_LC_9_20_5  (
            .in0(_gnd_net_),
            .in1(N__48543),
            .in2(_gnd_net_),
            .in3(N__46303),
            .lcout(\dron_frame_decoder_1.un1_sink_data_valid_5_i_0 ),
            .ltout(\dron_frame_decoder_1.un1_sink_data_valid_5_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNIA0H91_4_LC_9_20_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNIA0H91_4_LC_9_20_6 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNIA0H91_4_LC_9_20_6 .LUT_INIT=16'b1111111100000100;
    LogicCell40 \dron_frame_decoder_1.state_RNIA0H91_4_LC_9_20_6  (
            .in0(N__46330),
            .in1(N__46441),
            .in2(N__46342),
            .in3(N__86600),
            .lcout(\dron_frame_decoder_1.N_740_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNIBKSU_5_LC_9_20_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNIBKSU_5_LC_9_20_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNIBKSU_5_LC_9_20_7 .LUT_INIT=16'b1010111010101010;
    LogicCell40 \dron_frame_decoder_1.state_RNIBKSU_5_LC_9_20_7  (
            .in0(N__86601),
            .in1(N__48544),
            .in2(N__46338),
            .in3(N__46304),
            .lcout(\dron_frame_decoder_1.N_716_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNO_0_3_LC_9_21_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNO_0_3_LC_9_21_0 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNO_0_3_LC_9_21_0 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \dron_frame_decoder_1.state_RNO_0_3_LC_9_21_0  (
            .in0(N__48553),
            .in1(N__58035),
            .in2(N__57160),
            .in3(N__57328),
            .lcout(),
            .ltout(\dron_frame_decoder_1.state_ns_0_i_a2_0_2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_3_LC_9_21_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_3_LC_9_21_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_3_LC_9_21_1 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \dron_frame_decoder_1.state_3_LC_9_21_1  (
            .in0(N__46287),
            .in1(N__46450),
            .in2(N__46291),
            .in3(N__69274),
            .lcout(\dron_frame_decoder_1.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94340),
            .ce(),
            .sr(N__86412));
    defparam \dron_frame_decoder_1.state_RNO_1_3_LC_9_21_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNO_1_3_LC_9_21_2 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNO_1_3_LC_9_21_2 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \dron_frame_decoder_1.state_RNO_1_3_LC_9_21_2  (
            .in0(N__57952),
            .in1(N__48568),
            .in2(_gnd_net_),
            .in3(N__48870),
            .lcout(\dron_frame_decoder_1.state_ns_0_i_a2_0_3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_6_LC_9_21_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_6_LC_9_21_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_6_LC_9_21_3 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \dron_frame_decoder_1.state_6_LC_9_21_3  (
            .in0(N__46444),
            .in1(N__48555),
            .in2(N__69247),
            .in3(N__69275),
            .lcout(\dron_frame_decoder_1.stateZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94340),
            .ce(),
            .sr(N__86412));
    defparam \dron_frame_decoder_1.state_RNO_1_0_LC_9_21_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNO_1_0_LC_9_21_4 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNO_1_0_LC_9_21_4 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \dron_frame_decoder_1.state_RNO_1_0_LC_9_21_4  (
            .in0(N__48552),
            .in1(N__48869),
            .in2(N__48841),
            .in3(N__46442),
            .lcout(\dron_frame_decoder_1.N_200 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNO_2_0_LC_9_21_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNO_2_0_LC_9_21_5 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNO_2_0_LC_9_21_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \dron_frame_decoder_1.state_RNO_2_0_LC_9_21_5  (
            .in0(_gnd_net_),
            .in1(N__46439),
            .in2(_gnd_net_),
            .in3(N__48837),
            .lcout(\dron_frame_decoder_1.state_ns_i_a2_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_data_valid_LC_9_21_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_data_valid_LC_9_21_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_data_valid_LC_9_21_6 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \dron_frame_decoder_1.source_data_valid_LC_9_21_6  (
            .in0(N__48554),
            .in1(N__46443),
            .in2(_gnd_net_),
            .in3(N__69105),
            .lcout(debug_CH1_0A_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94340),
            .ce(),
            .sr(N__86412));
    defparam \pid_alt.state_RNIFCSD1_0_LC_9_21_7 .C_ON=1'b0;
    defparam \pid_alt.state_RNIFCSD1_0_LC_9_21_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.state_RNIFCSD1_0_LC_9_21_7 .LUT_INIT=16'b1100110011001110;
    LogicCell40 \pid_alt.state_RNIFCSD1_0_LC_9_21_7  (
            .in0(N__69104),
            .in1(N__71022),
            .in2(N__69079),
            .in3(N__68979),
            .lcout(\pid_alt.state_RNIFCSD1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNO_1_1_LC_9_22_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_1_1_LC_9_22_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_1_1_LC_9_22_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_RNO_1_1_LC_9_22_4  (
            .in0(_gnd_net_),
            .in1(N__92066),
            .in2(_gnd_net_),
            .in3(N__88256),
            .lcout(\Commands_frame_decoder.state_ns_0_a3_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_2_LC_9_23_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_2_LC_9_23_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_2_LC_9_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_2_LC_9_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46390),
            .lcout(\pid_front.error_p_regZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94364),
            .ce(N__93356),
            .sr(N__92990));
    defparam \ppm_encoder_1.counter24_0_I_1_c_LC_10_1_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_1_c_LC_10_1_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_1_c_LC_10_1_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_1_c_LC_10_1_0  (
            .in0(_gnd_net_),
            .in1(N__50266),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_1_0_),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_9_c_LC_10_1_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_9_c_LC_10_1_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_9_c_LC_10_1_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_9_c_LC_10_1_1  (
            .in0(_gnd_net_),
            .in1(N__50302),
            .in2(N__65865),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_0 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_15_c_LC_10_1_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_15_c_LC_10_1_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_15_c_LC_10_1_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_15_c_LC_10_1_2  (
            .in0(_gnd_net_),
            .in1(N__48811),
            .in2(N__65859),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_1 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_21_c_LC_10_1_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_21_c_LC_10_1_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_21_c_LC_10_1_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_21_c_LC_10_1_3  (
            .in0(_gnd_net_),
            .in1(N__49147),
            .in2(N__65862),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_2 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_27_c_LC_10_1_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_27_c_LC_10_1_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_27_c_LC_10_1_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_27_c_LC_10_1_4  (
            .in0(_gnd_net_),
            .in1(N__49861),
            .in2(N__65860),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_3 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_33_c_LC_10_1_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_33_c_LC_10_1_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_33_c_LC_10_1_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_33_c_LC_10_1_5  (
            .in0(_gnd_net_),
            .in1(N__50143),
            .in2(N__65863),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_4 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_39_c_LC_10_1_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_39_c_LC_10_1_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_39_c_LC_10_1_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_39_c_LC_10_1_6  (
            .in0(_gnd_net_),
            .in1(N__46669),
            .in2(N__65861),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_5 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_45_c_LC_10_1_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_45_c_LC_10_1_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_45_c_LC_10_1_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_45_c_LC_10_1_7  (
            .in0(_gnd_net_),
            .in1(N__52951),
            .in2(N__65864),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_6 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_51_c_LC_10_2_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_51_c_LC_10_2_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_51_c_LC_10_2_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_51_c_LC_10_2_0  (
            .in0(_gnd_net_),
            .in1(N__46675),
            .in2(N__65793),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_2_0_),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_57_c_LC_10_2_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_57_c_LC_10_2_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_57_c_LC_10_2_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_57_c_LC_10_2_1  (
            .in0(_gnd_net_),
            .in1(N__48982),
            .in2(N__65794),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_8 ),
            .carryout(\ppm_encoder_1.counter24_0_N_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_N_2_THRU_LUT4_0_LC_10_2_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_N_2_THRU_LUT4_0_LC_10_2_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_N_2_THRU_LUT4_0_LC_10_2_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.counter24_0_N_2_THRU_LUT4_0_LC_10_2_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46678),
            .lcout(\ppm_encoder_1.counter24_0_N_2_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_51_c_RNO_LC_10_2_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_51_c_RNO_LC_10_2_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_51_c_RNO_LC_10_2_5 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_51_c_RNO_LC_10_2_5  (
            .in0(N__49189),
            .in1(N__53262),
            .in2(N__49156),
            .in3(N__53292),
            .lcout(\ppm_encoder_1.counter24_0_I_51_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_39_c_RNO_LC_10_2_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_39_c_RNO_LC_10_2_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_39_c_RNO_LC_10_2_7 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_39_c_RNO_LC_10_2_7  (
            .in0(N__50671),
            .in1(N__53365),
            .in2(N__50716),
            .in3(N__53397),
            .lcout(\ppm_encoder_1.counter24_0_I_39_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_2_LC_10_3_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_2_LC_10_3_0 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_2_LC_10_3_0 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \ppm_encoder_1.init_pulses_2_LC_10_3_0  (
            .in0(N__49451),
            .in1(N__46663),
            .in2(N__49384),
            .in3(N__46651),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94090),
            .ce(),
            .sr(N__86504));
    defparam \ppm_encoder_1.init_pulses_5_LC_10_3_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_5_LC_10_3_1 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_5_LC_10_3_1 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \ppm_encoder_1.init_pulses_5_LC_10_3_1  (
            .in0(N__49369),
            .in1(N__49454),
            .in2(N__46609),
            .in3(N__46594),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94090),
            .ce(),
            .sr(N__86504));
    defparam \ppm_encoder_1.init_pulses_6_LC_10_3_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_6_LC_10_3_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_6_LC_10_3_2 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \ppm_encoder_1.init_pulses_6_LC_10_3_2  (
            .in0(N__49452),
            .in1(N__46588),
            .in2(N__49385),
            .in3(N__46576),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94090),
            .ce(),
            .sr(N__86504));
    defparam \ppm_encoder_1.init_pulses_7_LC_10_3_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_7_LC_10_3_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_7_LC_10_3_3 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \ppm_encoder_1.init_pulses_7_LC_10_3_3  (
            .in0(N__49370),
            .in1(N__49455),
            .in2(N__46570),
            .in3(N__46555),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94090),
            .ce(),
            .sr(N__86504));
    defparam \ppm_encoder_1.init_pulses_9_LC_10_3_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_9_LC_10_3_4 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_9_LC_10_3_4 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_9_LC_10_3_4  (
            .in0(N__49453),
            .in1(N__46549),
            .in2(N__49386),
            .in3(N__46543),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94090),
            .ce(),
            .sr(N__86504));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_10_LC_10_3_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_10_LC_10_3_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_10_LC_10_3_7 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_10_LC_10_3_7  (
            .in0(N__54255),
            .in1(N__46483),
            .in2(_gnd_net_),
            .in3(N__54110),
            .lcout(\ppm_encoder_1.N_378 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIVM131_0_16_LC_10_4_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIVM131_0_16_LC_10_4_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIVM131_0_16_LC_10_4_3 .LUT_INIT=16'b1111000001111000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIVM131_0_16_LC_10_4_3  (
            .in0(N__56270),
            .in1(N__49690),
            .in2(N__49219),
            .in3(N__52881),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIVM131_16_LC_10_4_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIVM131_16_LC_10_4_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIVM131_16_LC_10_4_4 .LUT_INIT=16'b1001110011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIVM131_16_LC_10_4_4  (
            .in0(N__52880),
            .in1(N__49217),
            .in2(N__49701),
            .in3(N__56269),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_8_LC_10_4_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_8_LC_10_4_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_8_LC_10_4_5 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \ppm_encoder_1.init_pulses_8_LC_10_4_5  (
            .in0(N__49444),
            .in1(N__46843),
            .in2(N__49383),
            .in3(N__46831),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94096),
            .ce(),
            .sr(N__86499));
    defparam \ppm_encoder_1.init_pulses_11_LC_10_4_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_11_LC_10_4_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_11_LC_10_4_6 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \ppm_encoder_1.init_pulses_11_LC_10_4_6  (
            .in0(N__49442),
            .in1(N__46825),
            .in2(N__49381),
            .in3(N__46813),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94096),
            .ce(),
            .sr(N__86499));
    defparam \ppm_encoder_1.init_pulses_12_LC_10_4_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_12_LC_10_4_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_12_LC_10_4_7 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \ppm_encoder_1.init_pulses_12_LC_10_4_7  (
            .in0(N__49443),
            .in1(N__46759),
            .in2(N__49382),
            .in3(N__46747),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94096),
            .ce(),
            .sr(N__86499));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_4_LC_10_5_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_4_LC_10_5_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_4_LC_10_5_0 .LUT_INIT=16'b0000101000100010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_4_LC_10_5_0  (
            .in0(N__54108),
            .in1(N__46740),
            .in2(N__46704),
            .in3(N__54250),
            .lcout(\ppm_encoder_1.pulses2count_9_i_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_4_LC_10_5_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_4_LC_10_5_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_4_LC_10_5_2 .LUT_INIT=16'b0111110100101000;
    LogicCell40 \ppm_encoder_1.elevator_4_LC_10_5_2  (
            .in0(N__51359),
            .in1(N__54979),
            .in2(N__47248),
            .in3(N__46700),
            .lcout(\ppm_encoder_1.elevatorZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94103),
            .ce(),
            .sr(N__86599));
    defparam \ppm_encoder_1.rudder_esr_ctle_14_LC_10_5_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_ctle_14_LC_10_5_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.rudder_esr_ctle_14_LC_10_5_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \ppm_encoder_1.rudder_esr_ctle_14_LC_10_5_3  (
            .in0(_gnd_net_),
            .in1(N__51357),
            .in2(_gnd_net_),
            .in3(N__86598),
            .lcout(\ppm_encoder_1.pid_altitude_dv_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_0_LC_10_5_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_0_LC_10_5_4 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_0_LC_10_5_4 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \ppm_encoder_1.elevator_0_LC_10_5_4  (
            .in0(N__51358),
            .in1(N__60271),
            .in2(_gnd_net_),
            .in3(N__47229),
            .lcout(\ppm_encoder_1.elevatorZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94103),
            .ce(),
            .sr(N__86599));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_0_LC_10_5_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_0_LC_10_5_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_0_LC_10_5_5 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_0_LC_10_5_5  (
            .in0(N__47228),
            .in1(N__56300),
            .in2(N__47212),
            .in3(N__47436),
            .lcout(\ppm_encoder_1.pulses2count_9_0_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m2_0_a2_0_a2_LC_10_5_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m2_0_a2_0_a2_LC_10_5_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m2_0_a2_0_a2_LC_10_5_6 .LUT_INIT=16'b0000000001110111;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m2_0_a2_0_a2_LC_10_5_6  (
            .in0(N__56299),
            .in1(N__49692),
            .in2(_gnd_net_),
            .in3(N__54249),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_ns_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m6_i_0_LC_10_5_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m6_i_0_LC_10_5_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m6_i_0_LC_10_5_7 .LUT_INIT=16'b1011101111001100;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m6_i_0_LC_10_5_7  (
            .in0(N__49691),
            .in1(N__56298),
            .in2(_gnd_net_),
            .in3(N__47435),
            .lcout(\ppm_encoder_1.N_56 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_10_LC_10_6_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_10_LC_10_6_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_10_LC_10_6_0 .LUT_INIT=16'b1111101011111110;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_10_LC_10_6_0  (
            .in0(N__53519),
            .in1(N__56239),
            .in2(N__47101),
            .in3(N__47089),
            .lcout(\ppm_encoder_1.pulses2count_9_i_0_2_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_4_LC_10_6_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_4_LC_10_6_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_4_LC_10_6_1 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_4_LC_10_6_1  (
            .in0(N__56241),
            .in1(N__53521),
            .in2(N__47062),
            .in3(N__47025),
            .lcout(\ppm_encoder_1.pulses2count_9_i_2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_esr_4_LC_10_6_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_4_LC_10_6_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_esr_4_LC_10_6_2 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \ppm_encoder_1.rudder_esr_4_LC_10_6_2  (
            .in0(_gnd_net_),
            .in1(N__47050),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\ppm_encoder_1.rudderZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94109),
            .ce(N__47954),
            .sr(N__86489));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_8_LC_10_6_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_8_LC_10_6_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_8_LC_10_6_3 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_8_LC_10_6_3  (
            .in0(N__56240),
            .in1(N__53520),
            .in2(N__47011),
            .in3(N__46996),
            .lcout(\ppm_encoder_1.pulses2count_9_i_2_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_9_LC_10_6_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_9_LC_10_6_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_9_LC_10_6_4 .LUT_INIT=16'b1111111110101110;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_9_LC_10_6_4  (
            .in0(N__53518),
            .in1(N__56236),
            .in2(N__46966),
            .in3(N__46933),
            .lcout(\ppm_encoder_1.pulses2count_9_i_2_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_0_i_LC_10_6_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_0_i_LC_10_6_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_0_i_LC_10_6_5 .LUT_INIT=16'b1011101110011001;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_0_i_LC_10_6_5  (
            .in0(N__56237),
            .in1(N__49672),
            .in2(_gnd_net_),
            .in3(N__47446),
            .lcout(\ppm_encoder_1.N_275 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIC2521_3_LC_10_6_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIC2521_3_LC_10_6_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIC2521_3_LC_10_6_6 .LUT_INIT=16'b1111010111110000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_RNIC2521_3_LC_10_6_6  (
            .in0(N__47447),
            .in1(_gnd_net_),
            .in2(N__49696),
            .in3(N__56238),
            .lcout(\ppm_encoder_1.N_304 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_3_LC_10_6_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_3_LC_10_6_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_3_LC_10_6_7 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_3_LC_10_6_7  (
            .in0(N__47553),
            .in1(N__47520),
            .in2(_gnd_net_),
            .in3(N__47445),
            .lcout(\ppm_encoder_1.pulses2count_9_0_0_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_0_c_LC_10_7_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_0_c_LC_10_7_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_0_c_LC_10_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_0_c_LC_10_7_0  (
            .in0(_gnd_net_),
            .in1(N__60267),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_7_0_),
            .carryout(\ppm_encoder_1.un1_elevator_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_0_THRU_LUT4_0_LC_10_7_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_0_THRU_LUT4_0_LC_10_7_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_0_THRU_LUT4_0_LC_10_7_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_0_THRU_LUT4_0_LC_10_7_1  (
            .in0(_gnd_net_),
            .in1(N__54996),
            .in2(N__65699),
            .in3(N__47278),
            .lcout(\ppm_encoder_1.un1_elevator_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_0 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_1_THRU_LUT4_0_LC_10_7_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_1_THRU_LUT4_0_LC_10_7_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_1_THRU_LUT4_0_LC_10_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_1_THRU_LUT4_0_LC_10_7_2  (
            .in0(_gnd_net_),
            .in1(N__60219),
            .in2(_gnd_net_),
            .in3(N__47263),
            .lcout(\ppm_encoder_1.un1_elevator_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_1 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_2_THRU_LUT4_0_LC_10_7_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_2_THRU_LUT4_0_LC_10_7_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_2_THRU_LUT4_0_LC_10_7_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_2_THRU_LUT4_0_LC_10_7_3  (
            .in0(_gnd_net_),
            .in1(N__60057),
            .in2(N__65700),
            .in3(N__47251),
            .lcout(\ppm_encoder_1.un1_elevator_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_2 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_3_THRU_LUT4_0_LC_10_7_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_3_THRU_LUT4_0_LC_10_7_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_3_THRU_LUT4_0_LC_10_7_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_3_THRU_LUT4_0_LC_10_7_4  (
            .in0(_gnd_net_),
            .in1(N__54975),
            .in2(_gnd_net_),
            .in3(N__47236),
            .lcout(\ppm_encoder_1.un1_elevator_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_3 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_4_THRU_LUT4_0_LC_10_7_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_4_THRU_LUT4_0_LC_10_7_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_4_THRU_LUT4_0_LC_10_7_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_4_THRU_LUT4_0_LC_10_7_5  (
            .in0(_gnd_net_),
            .in1(N__52533),
            .in2(_gnd_net_),
            .in3(N__47233),
            .lcout(\ppm_encoder_1.un1_elevator_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_4 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_5_THRU_LUT4_0_LC_10_7_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_5_THRU_LUT4_0_LC_10_7_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_5_THRU_LUT4_0_LC_10_7_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_5_THRU_LUT4_0_LC_10_7_6  (
            .in0(_gnd_net_),
            .in1(N__54603),
            .in2(N__65638),
            .in3(N__47659),
            .lcout(\ppm_encoder_1.un1_elevator_cry_5_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_5 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_6_THRU_LUT4_0_LC_10_7_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_6_THRU_LUT4_0_LC_10_7_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_6_THRU_LUT4_0_LC_10_7_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_6_THRU_LUT4_0_LC_10_7_7  (
            .in0(_gnd_net_),
            .in1(N__54570),
            .in2(_gnd_net_),
            .in3(N__47656),
            .lcout(\ppm_encoder_1.un1_elevator_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_6 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_7_THRU_LUT4_0_LC_10_8_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_7_THRU_LUT4_0_LC_10_8_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_7_THRU_LUT4_0_LC_10_8_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_7_THRU_LUT4_0_LC_10_8_0  (
            .in0(_gnd_net_),
            .in1(N__54543),
            .in2(_gnd_net_),
            .in3(N__47638),
            .lcout(\ppm_encoder_1.un1_elevator_cry_7_THRU_CO ),
            .ltout(),
            .carryin(bfn_10_8_0_),
            .carryout(\ppm_encoder_1.un1_elevator_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_8_THRU_LUT4_0_LC_10_8_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_8_THRU_LUT4_0_LC_10_8_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_8_THRU_LUT4_0_LC_10_8_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_8_THRU_LUT4_0_LC_10_8_1  (
            .in0(_gnd_net_),
            .in1(N__54510),
            .in2(_gnd_net_),
            .in3(N__47629),
            .lcout(\ppm_encoder_1.un1_elevator_cry_8_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_8 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_9_THRU_LUT4_0_LC_10_8_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_9_THRU_LUT4_0_LC_10_8_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_9_THRU_LUT4_0_LC_10_8_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_9_THRU_LUT4_0_LC_10_8_2  (
            .in0(_gnd_net_),
            .in1(N__54672),
            .in2(_gnd_net_),
            .in3(N__47617),
            .lcout(\ppm_encoder_1.un1_elevator_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_9 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_10_THRU_LUT4_0_LC_10_8_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_10_THRU_LUT4_0_LC_10_8_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_10_THRU_LUT4_0_LC_10_8_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_10_THRU_LUT4_0_LC_10_8_3  (
            .in0(_gnd_net_),
            .in1(N__54642),
            .in2(_gnd_net_),
            .in3(N__47605),
            .lcout(\ppm_encoder_1.un1_elevator_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_10 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_11_THRU_LUT4_0_LC_10_8_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_11_THRU_LUT4_0_LC_10_8_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_11_THRU_LUT4_0_LC_10_8_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_11_THRU_LUT4_0_LC_10_8_4  (
            .in0(_gnd_net_),
            .in1(N__55701),
            .in2(_gnd_net_),
            .in3(N__47587),
            .lcout(\ppm_encoder_1.un1_elevator_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_11 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_12_THRU_LUT4_0_LC_10_8_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_12_THRU_LUT4_0_LC_10_8_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_12_THRU_LUT4_0_LC_10_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_12_THRU_LUT4_0_LC_10_8_5  (
            .in0(_gnd_net_),
            .in1(N__55743),
            .in2(N__65628),
            .in3(N__47572),
            .lcout(\ppm_encoder_1.un1_elevator_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_12 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_esr_14_LC_10_8_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_esr_14_LC_10_8_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_esr_14_LC_10_8_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.elevator_esr_14_LC_10_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47569),
            .lcout(\ppm_encoder_1.elevatorZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94126),
            .ce(N__47980),
            .sr(N__86472));
    defparam CONSTANT_ONE_LUT4_LC_10_8_7.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_10_8_7.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_10_8_7.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_10_8_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.bit_Count_RNIJOJC1_2_LC_10_9_2 .C_ON=1'b0;
    defparam \uart_drone.bit_Count_RNIJOJC1_2_LC_10_9_2 .SEQ_MODE=4'b0000;
    defparam \uart_drone.bit_Count_RNIJOJC1_2_LC_10_9_2 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \uart_drone.bit_Count_RNIJOJC1_2_LC_10_9_2  (
            .in0(N__56594),
            .in1(_gnd_net_),
            .in2(N__56543),
            .in3(N__56467),
            .lcout(\uart_drone.N_152 ),
            .ltout(\uart_drone.N_152_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNI63LK2_3_LC_10_9_3 .C_ON=1'b0;
    defparam \uart_drone.state_RNI63LK2_3_LC_10_9_3 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNI63LK2_3_LC_10_9_3 .LUT_INIT=16'b1010000010101010;
    LogicCell40 \uart_drone.state_RNI63LK2_3_LC_10_9_3  (
            .in0(N__51459),
            .in1(_gnd_net_),
            .in2(N__47743),
            .in3(N__53974),
            .lcout(\uart_drone.un1_state_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.bit_Count_RNO_0_2_LC_10_9_4 .C_ON=1'b0;
    defparam \uart_drone.bit_Count_RNO_0_2_LC_10_9_4 .SEQ_MODE=4'b0000;
    defparam \uart_drone.bit_Count_RNO_0_2_LC_10_9_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uart_drone.bit_Count_RNO_0_2_LC_10_9_4  (
            .in0(N__56595),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51458),
            .lcout(\uart_drone.CO0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_12_LC_10_9_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_12_LC_10_9_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_12_LC_10_9_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_12_LC_10_9_6  (
            .in0(_gnd_net_),
            .in1(N__50583),
            .in2(_gnd_net_),
            .in3(N__47725),
            .lcout(\ppm_encoder_1.N_436 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNO_0_3_LC_10_9_7 .C_ON=1'b0;
    defparam \uart_drone.state_RNO_0_3_LC_10_9_7 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNO_0_3_LC_10_9_7 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \uart_drone.state_RNO_0_3_LC_10_9_7  (
            .in0(N__53975),
            .in1(N__51519),
            .in2(N__51592),
            .in3(N__54782),
            .lcout(\uart_drone.N_145 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_0_c_LC_10_10_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_0_c_LC_10_10_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_0_c_LC_10_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_0_c_LC_10_10_0  (
            .in0(_gnd_net_),
            .in1(N__59176),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_10_0_),
            .carryout(\ppm_encoder_1.un1_aileron_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_0_THRU_LUT4_0_LC_10_10_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_0_THRU_LUT4_0_LC_10_10_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_0_THRU_LUT4_0_LC_10_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_0_THRU_LUT4_0_LC_10_10_1  (
            .in0(_gnd_net_),
            .in1(N__56055),
            .in2(N__65704),
            .in3(N__47689),
            .lcout(\ppm_encoder_1.un1_aileron_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_0 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_1_THRU_LUT4_0_LC_10_10_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_1_THRU_LUT4_0_LC_10_10_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_1_THRU_LUT4_0_LC_10_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_1_THRU_LUT4_0_LC_10_10_2  (
            .in0(_gnd_net_),
            .in1(N__56031),
            .in2(_gnd_net_),
            .in3(N__47674),
            .lcout(\ppm_encoder_1.un1_aileron_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_1 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_2_THRU_LUT4_0_LC_10_10_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_2_THRU_LUT4_0_LC_10_10_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_2_THRU_LUT4_0_LC_10_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_2_THRU_LUT4_0_LC_10_10_3  (
            .in0(_gnd_net_),
            .in1(N__56004),
            .in2(N__65705),
            .in3(N__47842),
            .lcout(\ppm_encoder_1.un1_aileron_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_2 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_3_THRU_LUT4_0_LC_10_10_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_3_THRU_LUT4_0_LC_10_10_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_3_THRU_LUT4_0_LC_10_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_3_THRU_LUT4_0_LC_10_10_4  (
            .in0(_gnd_net_),
            .in1(N__59331),
            .in2(_gnd_net_),
            .in3(N__47833),
            .lcout(\ppm_encoder_1.un1_aileron_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_3 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_4_THRU_LUT4_0_LC_10_10_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_4_THRU_LUT4_0_LC_10_10_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_4_THRU_LUT4_0_LC_10_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_4_THRU_LUT4_0_LC_10_10_5  (
            .in0(_gnd_net_),
            .in1(N__59283),
            .in2(_gnd_net_),
            .in3(N__47815),
            .lcout(\ppm_encoder_1.un1_aileron_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_4 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_5_THRU_LUT4_0_LC_10_10_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_5_THRU_LUT4_0_LC_10_10_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_5_THRU_LUT4_0_LC_10_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_5_THRU_LUT4_0_LC_10_10_6  (
            .in0(_gnd_net_),
            .in1(N__65645),
            .in2(N__54451),
            .in3(N__47806),
            .lcout(\ppm_encoder_1.un1_aileron_cry_5_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_5 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_6_THRU_LUT4_0_LC_10_10_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_6_THRU_LUT4_0_LC_10_10_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_6_THRU_LUT4_0_LC_10_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_6_THRU_LUT4_0_LC_10_10_7  (
            .in0(_gnd_net_),
            .in1(N__54414),
            .in2(_gnd_net_),
            .in3(N__47791),
            .lcout(\ppm_encoder_1.un1_aileron_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_6 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_7_THRU_LUT4_0_LC_10_11_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_7_THRU_LUT4_0_LC_10_11_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_7_THRU_LUT4_0_LC_10_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_7_THRU_LUT4_0_LC_10_11_0  (
            .in0(_gnd_net_),
            .in1(N__54384),
            .in2(_gnd_net_),
            .in3(N__47776),
            .lcout(\ppm_encoder_1.un1_aileron_cry_7_THRU_CO ),
            .ltout(),
            .carryin(bfn_10_11_0_),
            .carryout(\ppm_encoder_1.un1_aileron_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_8_THRU_LUT4_0_LC_10_11_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_8_THRU_LUT4_0_LC_10_11_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_8_THRU_LUT4_0_LC_10_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_8_THRU_LUT4_0_LC_10_11_1  (
            .in0(_gnd_net_),
            .in1(N__54348),
            .in2(_gnd_net_),
            .in3(N__47761),
            .lcout(\ppm_encoder_1.un1_aileron_cry_8_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_8 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_9_THRU_LUT4_0_LC_10_11_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_9_THRU_LUT4_0_LC_10_11_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_9_THRU_LUT4_0_LC_10_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_9_THRU_LUT4_0_LC_10_11_2  (
            .in0(_gnd_net_),
            .in1(N__53454),
            .in2(_gnd_net_),
            .in3(N__47746),
            .lcout(\ppm_encoder_1.un1_aileron_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_9 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_10_THRU_LUT4_0_LC_10_11_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_10_THRU_LUT4_0_LC_10_11_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_10_THRU_LUT4_0_LC_10_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_10_THRU_LUT4_0_LC_10_11_3  (
            .in0(_gnd_net_),
            .in1(N__54484),
            .in2(_gnd_net_),
            .in3(N__48010),
            .lcout(\ppm_encoder_1.un1_aileron_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_10 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_11_THRU_LUT4_0_LC_10_11_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_11_THRU_LUT4_0_LC_10_11_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_11_THRU_LUT4_0_LC_10_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_11_THRU_LUT4_0_LC_10_11_4  (
            .in0(_gnd_net_),
            .in1(N__53185),
            .in2(_gnd_net_),
            .in3(N__47995),
            .lcout(\ppm_encoder_1.un1_aileron_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_11 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_12_THRU_LUT4_0_LC_10_11_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_12_THRU_LUT4_0_LC_10_11_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_12_THRU_LUT4_0_LC_10_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_12_THRU_LUT4_0_LC_10_11_5  (
            .in0(_gnd_net_),
            .in1(N__53932),
            .in2(N__65706),
            .in3(N__47992),
            .lcout(\ppm_encoder_1.un1_aileron_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_12 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_esr_14_LC_10_11_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_14_LC_10_11_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_esr_14_LC_10_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.aileron_esr_14_LC_10_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47989),
            .lcout(\ppm_encoder_1.aileronZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94154),
            .ce(N__47973),
            .sr(N__86456));
    defparam \uart_drone.timer_Count_RNI5A9J_1_LC_10_12_0 .C_ON=1'b1;
    defparam \uart_drone.timer_Count_RNI5A9J_1_LC_10_12_0 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNI5A9J_1_LC_10_12_0 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \uart_drone.timer_Count_RNI5A9J_1_LC_10_12_0  (
            .in0(N__47908),
            .in1(N__51018),
            .in2(N__47913),
            .in3(_gnd_net_),
            .lcout(\uart_drone.un1_state_2_0_a3_0 ),
            .ltout(),
            .carryin(bfn_10_12_0_),
            .carryout(\uart_drone.un4_timer_Count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNO_0_2_LC_10_12_1 .C_ON=1'b1;
    defparam \uart_drone.timer_Count_RNO_0_2_LC_10_12_1 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNO_0_2_LC_10_12_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_drone.timer_Count_RNO_0_2_LC_10_12_1  (
            .in0(_gnd_net_),
            .in1(N__47886),
            .in2(_gnd_net_),
            .in3(N__47863),
            .lcout(\uart_drone.timer_Count_RNO_0_0_2 ),
            .ltout(),
            .carryin(\uart_drone.un4_timer_Count_1_cry_1 ),
            .carryout(\uart_drone.un4_timer_Count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNO_0_3_LC_10_12_2 .C_ON=1'b1;
    defparam \uart_drone.timer_Count_RNO_0_3_LC_10_12_2 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNO_0_3_LC_10_12_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_drone.timer_Count_RNO_0_3_LC_10_12_2  (
            .in0(_gnd_net_),
            .in1(N__51509),
            .in2(_gnd_net_),
            .in3(N__47860),
            .lcout(\uart_drone.timer_Count_RNO_0_0_3 ),
            .ltout(),
            .carryin(\uart_drone.un4_timer_Count_1_cry_2 ),
            .carryout(\uart_drone.un4_timer_Count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNO_0_4_LC_10_12_3 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNO_0_4_LC_10_12_3 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNO_0_4_LC_10_12_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uart_drone.timer_Count_RNO_0_4_LC_10_12_3  (
            .in0(_gnd_net_),
            .in1(N__54772),
            .in2(_gnd_net_),
            .in3(N__47857),
            .lcout(\uart_drone.timer_Count_RNO_0_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNIES9Q1_2_LC_10_12_4 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNIES9Q1_2_LC_10_12_4 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNIES9Q1_2_LC_10_12_4 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \uart_drone.timer_Count_RNIES9Q1_2_LC_10_12_4  (
            .in0(N__56798),
            .in1(N__48194),
            .in2(_gnd_net_),
            .in3(N__70794),
            .lcout(\uart_drone.timer_Count_RNIES9Q1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNIRC5U2_2_LC_10_12_5 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNIRC5U2_2_LC_10_12_5 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNIRC5U2_2_LC_10_12_5 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \uart_drone.timer_Count_RNIRC5U2_2_LC_10_12_5  (
            .in0(N__48195),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56949),
            .lcout(\uart_drone.data_rdyc_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_4_LC_10_12_6 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_4_LC_10_12_6 .SEQ_MODE=4'b1000;
    defparam \uart_drone.timer_Count_4_LC_10_12_6 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \uart_drone.timer_Count_4_LC_10_12_6  (
            .in0(N__50783),
            .in1(N__70796),
            .in2(N__48181),
            .in3(N__51561),
            .lcout(\uart_drone.timer_CountZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94166),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_3_LC_10_12_7 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_3_LC_10_12_7 .SEQ_MODE=4'b1000;
    defparam \uart_drone.timer_Count_3_LC_10_12_7 .LUT_INIT=16'b0100010001000000;
    LogicCell40 \uart_drone.timer_Count_3_LC_10_12_7  (
            .in0(N__70795),
            .in1(N__48169),
            .in2(N__51567),
            .in3(N__50782),
            .lcout(\uart_drone.timer_CountZ1Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94166),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone_sync.aux_2__0__0_LC_10_13_1 .C_ON=1'b0;
    defparam \uart_drone_sync.aux_2__0__0_LC_10_13_1 .SEQ_MODE=4'b1000;
    defparam \uart_drone_sync.aux_2__0__0_LC_10_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone_sync.aux_2__0__0_LC_10_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48163),
            .lcout(\uart_drone_sync.aux_2__0__0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94179),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc_sync.aux_2__0__0_LC_10_13_2 .C_ON=1'b0;
    defparam \uart_pc_sync.aux_2__0__0_LC_10_13_2 .SEQ_MODE=4'b1000;
    defparam \uart_pc_sync.aux_2__0__0_LC_10_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_pc_sync.aux_2__0__0_LC_10_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48145),
            .lcout(\uart_pc_sync.aux_2__0_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94179),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc_sync.aux_3__0__0_LC_10_13_3 .C_ON=1'b0;
    defparam \uart_pc_sync.aux_3__0__0_LC_10_13_3 .SEQ_MODE=4'b1000;
    defparam \uart_pc_sync.aux_3__0__0_LC_10_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_pc_sync.aux_3__0__0_LC_10_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48130),
            .lcout(\uart_pc_sync.aux_3__0_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94179),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc_sync.Q_0__0_LC_10_13_7 .C_ON=1'b0;
    defparam \uart_pc_sync.Q_0__0_LC_10_13_7 .SEQ_MODE=4'b1000;
    defparam \uart_pc_sync.Q_0__0_LC_10_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_pc_sync.Q_0__0_LC_10_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48124),
            .lcout(debug_CH2_18A_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94179),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.source_data_1_esr_ctle_14_LC_10_14_3 .C_ON=1'b0;
    defparam \scaler_4.source_data_1_esr_ctle_14_LC_10_14_3 .SEQ_MODE=4'b0000;
    defparam \scaler_4.source_data_1_esr_ctle_14_LC_10_14_3 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \scaler_4.source_data_1_esr_ctle_14_LC_10_14_3  (
            .in0(N__48107),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86595),
            .lcout(\scaler_4.debug_CH3_20A_c_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIG48S_7_LC_10_14_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIG48S_7_LC_10_14_5 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIG48S_7_LC_10_14_5 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \Commands_frame_decoder.state_RNIG48S_7_LC_10_14_5  (
            .in0(N__52045),
            .in1(N__55262),
            .in2(_gnd_net_),
            .in3(N__70880),
            .lcout(\Commands_frame_decoder.state_RNIG48SZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_12_LC_10_15_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_12_LC_10_15_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_12_LC_10_15_0 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \Commands_frame_decoder.state_12_LC_10_15_0  (
            .in0(N__48597),
            .in1(N__55241),
            .in2(N__51630),
            .in3(N__69371),
            .lcout(\Commands_frame_decoder.stateZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94208),
            .ce(),
            .sr(N__86442));
    defparam \Commands_frame_decoder.WDT_RNIPRJG5_0_14_LC_10_15_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNIPRJG5_0_14_LC_10_15_1 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNIPRJG5_0_14_LC_10_15_1 .LUT_INIT=16'b0000010100010101;
    LogicCell40 \Commands_frame_decoder.WDT_RNIPRJG5_0_14_LC_10_15_1  (
            .in0(N__55240),
            .in1(N__48346),
            .in2(N__48334),
            .in3(N__48295),
            .lcout(\Commands_frame_decoder.N_403 ),
            .ltout(\Commands_frame_decoder.N_403_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_11_LC_10_15_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_11_LC_10_15_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_11_LC_10_15_2 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \Commands_frame_decoder.state_11_LC_10_15_2  (
            .in0(N__51626),
            .in1(N__48265),
            .in2(N__48232),
            .in3(N__55247),
            .lcout(\Commands_frame_decoder.stateZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94208),
            .ce(),
            .sr(N__86442));
    defparam \Commands_frame_decoder.state_8_LC_10_15_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_8_LC_10_15_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_8_LC_10_15_4 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \Commands_frame_decoder.state_8_LC_10_15_4  (
            .in0(N__52049),
            .in1(N__55243),
            .in2(N__48229),
            .in3(N__69374),
            .lcout(\Commands_frame_decoder.stateZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94208),
            .ce(),
            .sr(N__86442));
    defparam \Commands_frame_decoder.state_9_LC_10_15_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_9_LC_10_15_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_9_LC_10_15_5 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \Commands_frame_decoder.state_9_LC_10_15_5  (
            .in0(N__69375),
            .in1(N__48225),
            .in2(N__55269),
            .in3(N__48217),
            .lcout(\Commands_frame_decoder.stateZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94208),
            .ce(),
            .sr(N__86442));
    defparam \Commands_frame_decoder.state_7_LC_10_15_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_7_LC_10_15_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_7_LC_10_15_6 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \Commands_frame_decoder.state_7_LC_10_15_6  (
            .in0(N__52105),
            .in1(N__55242),
            .in2(N__52056),
            .in3(N__69373),
            .lcout(\Commands_frame_decoder.stateZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94208),
            .ce(),
            .sr(N__86442));
    defparam \Commands_frame_decoder.state_6_LC_10_15_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_6_LC_10_15_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_6_LC_10_15_7 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \Commands_frame_decoder.state_6_LC_10_15_7  (
            .in0(N__69372),
            .in1(N__52106),
            .in2(_gnd_net_),
            .in3(N__51939),
            .lcout(\Commands_frame_decoder.stateZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94208),
            .ce(),
            .sr(N__86442));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_7_LC_10_16_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_7_LC_10_16_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_7_LC_10_16_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_7_LC_10_16_1  (
            .in0(N__57789),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\dron_frame_decoder_1.drone_H_disp_side_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94225),
            .ce(N__57072),
            .sr(N__86438));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIKAP4_8_LC_10_16_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIKAP4_8_LC_10_16_2 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIKAP4_8_LC_10_16_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_RNIKAP4_8_LC_10_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52276),
            .lcout(drone_H_disp_side_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNILBP4_9_LC_10_16_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNILBP4_9_LC_10_16_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNILBP4_9_LC_10_16_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_RNILBP4_9_LC_10_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52270),
            .lcout(drone_H_disp_side_i_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIT4RD_10_LC_10_16_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIT4RD_10_LC_10_16_4 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIT4RD_10_LC_10_16_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_RNIT4RD_10_LC_10_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51925),
            .lcout(drone_H_disp_side_i_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIV6RD_12_LC_10_16_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIV6RD_12_LC_10_16_5 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIV6RD_12_LC_10_16_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_RNIV6RD_12_LC_10_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77465),
            .lcout(drone_H_disp_side_i_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_axb_1_LC_10_16_6 .C_ON=1'b0;
    defparam \pid_alt.error_axb_1_LC_10_16_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_axb_1_LC_10_16_6 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pid_alt.error_axb_1_LC_10_16_6  (
            .in0(_gnd_net_),
            .in1(N__48358),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_axbZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_axb_12_LC_10_16_7 .C_ON=1'b0;
    defparam \pid_alt.error_axb_12_LC_10_16_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_axb_12_LC_10_16_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_axb_12_LC_10_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48460),
            .lcout(\pid_alt.error_axbZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_0_LC_10_17_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_0_LC_10_17_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_0_LC_10_17_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_0_LC_10_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57723),
            .lcout(drone_altitude_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94242),
            .ce(N__48472),
            .sr(N__86432));
    defparam \dron_frame_decoder_1.source_Altitude_esr_1_LC_10_17_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_1_LC_10_17_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_1_LC_10_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_1_LC_10_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57318),
            .lcout(drone_altitude_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94242),
            .ce(N__48472),
            .sr(N__86432));
    defparam \dron_frame_decoder_1.source_Altitude_esr_2_LC_10_17_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_2_LC_10_17_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_2_LC_10_17_2 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_2_LC_10_17_2  (
            .in0(_gnd_net_),
            .in1(N__57242),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(drone_altitude_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94242),
            .ce(N__48472),
            .sr(N__86432));
    defparam \dron_frame_decoder_1.source_Altitude_esr_3_LC_10_17_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_3_LC_10_17_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_3_LC_10_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_3_LC_10_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58029),
            .lcout(drone_altitude_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94242),
            .ce(N__48472),
            .sr(N__86432));
    defparam \dron_frame_decoder_1.source_Altitude_esr_4_LC_10_17_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_4_LC_10_17_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_4_LC_10_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_4_LC_10_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57939),
            .lcout(\dron_frame_decoder_1.drone_altitude_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94242),
            .ce(N__48472),
            .sr(N__86432));
    defparam \dron_frame_decoder_1.source_Altitude_esr_5_LC_10_17_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_5_LC_10_17_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_5_LC_10_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_5_LC_10_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57869),
            .lcout(\dron_frame_decoder_1.drone_altitude_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94242),
            .ce(N__48472),
            .sr(N__86432));
    defparam \dron_frame_decoder_1.source_Altitude_esr_6_LC_10_17_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_6_LC_10_17_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_6_LC_10_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_6_LC_10_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57151),
            .lcout(\dron_frame_decoder_1.drone_altitude_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94242),
            .ce(N__48472),
            .sr(N__86432));
    defparam \dron_frame_decoder_1.source_Altitude_esr_7_LC_10_17_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_7_LC_10_17_7 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_7_LC_10_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_7_LC_10_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57790),
            .lcout(\dron_frame_decoder_1.drone_altitude_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94242),
            .ce(N__48472),
            .sr(N__86432));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_1_LC_10_18_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_1_LC_10_18_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_1_LC_10_18_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_1_LC_10_18_0  (
            .in0(N__57325),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(drone_H_disp_front_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94259),
            .ce(N__57413),
            .sr(N__86424));
    defparam \dron_frame_decoder_1.source_Altitude_esr_10_LC_10_19_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_10_LC_10_19_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_10_LC_10_19_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_10_LC_10_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57249),
            .lcout(\dron_frame_decoder_1.drone_altitude_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94278),
            .ce(N__52329),
            .sr(N__86413));
    defparam \dron_frame_decoder_1.source_Altitude_esr_11_LC_10_19_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_11_LC_10_19_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_11_LC_10_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_11_LC_10_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58036),
            .lcout(\dron_frame_decoder_1.drone_altitude_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94278),
            .ce(N__52329),
            .sr(N__86413));
    defparam \dron_frame_decoder_1.source_Altitude_esr_12_LC_10_19_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_12_LC_10_19_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_12_LC_10_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_12_LC_10_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57946),
            .lcout(drone_altitude_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94278),
            .ce(N__52329),
            .sr(N__86413));
    defparam \dron_frame_decoder_1.source_Altitude_esr_15_LC_10_19_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_15_LC_10_19_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_15_LC_10_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_15_LC_10_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57791),
            .lcout(drone_altitude_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94278),
            .ce(N__52329),
            .sr(N__86413));
    defparam \dron_frame_decoder_1.source_Altitude_esr_8_LC_10_19_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_8_LC_10_19_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_8_LC_10_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_8_LC_10_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57727),
            .lcout(\dron_frame_decoder_1.drone_altitude_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94278),
            .ce(N__52329),
            .sr(N__86413));
    defparam \dron_frame_decoder_1.source_Altitude_esr_9_LC_10_19_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_9_LC_10_19_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_9_LC_10_19_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_9_LC_10_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57326),
            .lcout(\dron_frame_decoder_1.drone_altitude_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94278),
            .ce(N__52329),
            .sr(N__86413));
    defparam \Commands_frame_decoder.state_RNIF38S_6_LC_10_20_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIF38S_6_LC_10_20_0 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIF38S_6_LC_10_20_0 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \Commands_frame_decoder.state_RNIF38S_6_LC_10_20_0  (
            .in0(N__52107),
            .in1(N__55257),
            .in2(_gnd_net_),
            .in3(N__70964),
            .lcout(\Commands_frame_decoder.state_RNIF38SZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNIAD5K1_7_LC_10_20_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNIAD5K1_7_LC_10_20_1 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNIAD5K1_7_LC_10_20_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \dron_frame_decoder_1.state_RNIAD5K1_7_LC_10_20_1  (
            .in0(_gnd_net_),
            .in1(N__48652),
            .in2(_gnd_net_),
            .in3(N__86586),
            .lcout(\dron_frame_decoder_1.N_732_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIUHR9_10_LC_10_20_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIUHR9_10_LC_10_20_2 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIUHR9_10_LC_10_20_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNIUHR9_10_LC_10_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48646),
            .lcout(drone_altitude_i_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNITUI31_13_LC_10_20_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNITUI31_13_LC_10_20_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNITUI31_13_LC_10_20_4 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \Commands_frame_decoder.state_RNITUI31_13_LC_10_20_4  (
            .in0(N__48624),
            .in1(N__55256),
            .in2(_gnd_net_),
            .in3(N__70963),
            .lcout(\Commands_frame_decoder.state_RNITUI31Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIVGCQ_12_LC_10_20_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIVGCQ_12_LC_10_20_6 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIVGCQ_12_LC_10_20_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_RNIVGCQ_12_LC_10_20_6  (
            .in0(_gnd_net_),
            .in1(N__48598),
            .in2(_gnd_net_),
            .in3(N__55255),
            .lcout(\Commands_frame_decoder.source_xy_ki_1_sqmuxa ),
            .ltout(\Commands_frame_decoder.source_xy_ki_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNI61EQ_12_LC_10_20_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNI61EQ_12_LC_10_20_7 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNI61EQ_12_LC_10_20_7 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \Commands_frame_decoder.state_RNI61EQ_12_LC_10_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__48571),
            .in3(N__86585),
            .lcout(\Commands_frame_decoder.source_xy_ki_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_ns_0_i_a2_0_5_3_LC_10_21_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_ns_0_i_a2_0_5_3_LC_10_21_0 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_ns_0_i_a2_0_5_3_LC_10_21_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \dron_frame_decoder_1.state_ns_0_i_a2_0_5_3_LC_10_21_0  (
            .in0(N__57871),
            .in1(N__57248),
            .in2(N__57793),
            .in3(N__57721),
            .lcout(\dron_frame_decoder_1.N_230_5 ),
            .ltout(\dron_frame_decoder_1.N_230_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_ns_i_a2_2_0_a2_0_LC_10_21_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_ns_i_a2_2_0_a2_0_LC_10_21_1 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_ns_i_a2_2_0_a2_0_LC_10_21_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \dron_frame_decoder_1.state_ns_i_a2_2_0_a2_0_LC_10_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__48562),
            .in3(N__48551),
            .lcout(\dron_frame_decoder_1.N_224 ),
            .ltout(\dron_frame_decoder_1.N_224_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNO_0_0_LC_10_21_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNO_0_0_LC_10_21_2 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNO_0_0_LC_10_21_2 .LUT_INIT=16'b1111000010000000;
    LogicCell40 \dron_frame_decoder_1.state_RNO_0_0_LC_10_21_2  (
            .in0(N__48820),
            .in1(N__48901),
            .in2(N__48895),
            .in3(N__48889),
            .lcout(\dron_frame_decoder_1.N_198 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_ns_i_a2_1_1_0_LC_10_21_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_ns_i_a2_1_1_0_LC_10_21_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_ns_i_a2_1_1_0_LC_10_21_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \dron_frame_decoder_1.state_ns_i_a2_1_1_0_LC_10_21_3  (
            .in0(_gnd_net_),
            .in1(N__58033),
            .in2(_gnd_net_),
            .in3(N__57320),
            .lcout(),
            .ltout(\dron_frame_decoder_1.state_ns_i_a2_1_1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNIN9KQ1_0_LC_10_21_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNIN9KQ1_0_LC_10_21_4 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNIN9KQ1_0_LC_10_21_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \dron_frame_decoder_1.state_RNIN9KQ1_0_LC_10_21_4  (
            .in0(N__57155),
            .in1(N__57942),
            .in2(N__48892),
            .in3(N__48835),
            .lcout(\dron_frame_decoder_1.N_220 ),
            .ltout(\dron_frame_decoder_1.N_220_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_1_LC_10_21_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_1_LC_10_21_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_1_LC_10_21_5 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \dron_frame_decoder_1.state_1_LC_10_21_5  (
            .in0(N__48871),
            .in1(N__48883),
            .in2(N__48874),
            .in3(N__69290),
            .lcout(\dron_frame_decoder_1.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94309),
            .ce(),
            .sr(N__86393));
    defparam \dron_frame_decoder_1.state_0_LC_10_21_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_0_LC_10_21_6 .SEQ_MODE=4'b1001;
    defparam \dron_frame_decoder_1.state_0_LC_10_21_6 .LUT_INIT=16'b0000000000001101;
    LogicCell40 \dron_frame_decoder_1.state_0_LC_10_21_6  (
            .in0(N__69291),
            .in1(N__48836),
            .in2(N__48856),
            .in3(N__48847),
            .lcout(\dron_frame_decoder_1.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94309),
            .ce(),
            .sr(N__86393));
    defparam \dron_frame_decoder_1.state_RNO_3_0_LC_10_21_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNO_3_0_LC_10_21_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNO_3_0_LC_10_21_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \dron_frame_decoder_1.state_RNO_3_0_LC_10_21_7  (
            .in0(N__57941),
            .in1(N__58034),
            .in2(N__57159),
            .in3(N__57321),
            .lcout(\dron_frame_decoder_1.state_ns_i_a2_0_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_15_c_RNO_LC_11_1_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_15_c_RNO_LC_11_1_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_15_c_RNO_LC_11_1_0 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_15_c_RNO_LC_11_1_0  (
            .in0(N__53108),
            .in1(N__49981),
            .in2(N__49900),
            .in3(N__53129),
            .lcout(\ppm_encoder_1.counter24_0_I_15_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_15_LC_11_1_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_15_LC_11_1_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_15_LC_11_1_3 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_15_LC_11_1_3  (
            .in0(N__50983),
            .in1(N__48805),
            .in2(_gnd_net_),
            .in3(N__49699),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94080),
            .ce(N__50349),
            .sr(N__86507));
    defparam \ppm_encoder_1.pulses2count_esr_14_LC_11_1_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_14_LC_11_1_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_14_LC_11_1_5 .LUT_INIT=16'b0000000000001101;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_14_LC_11_1_5  (
            .in0(N__50986),
            .in1(N__48772),
            .in2(N__53848),
            .in3(N__48736),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94080),
            .ce(N__50349),
            .sr(N__86507));
    defparam \ppm_encoder_1.pulses2count_esr_16_LC_11_1_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_16_LC_11_1_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_16_LC_11_1_6 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_16_LC_11_1_6  (
            .in0(N__49698),
            .in1(N__49218),
            .in2(_gnd_net_),
            .in3(N__50984),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94080),
            .ce(N__50349),
            .sr(N__86507));
    defparam \ppm_encoder_1.pulses2count_esr_17_LC_11_1_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_17_LC_11_1_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_17_LC_11_1_7 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_17_LC_11_1_7  (
            .in0(N__50985),
            .in1(N__49183),
            .in2(_gnd_net_),
            .in3(N__49700),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94080),
            .ce(N__50349),
            .sr(N__86507));
    defparam \ppm_encoder_1.counter24_0_I_21_c_RNO_LC_11_2_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_21_c_RNO_LC_11_2_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_21_c_RNO_LC_11_2_0 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_21_c_RNO_LC_11_2_0  (
            .in0(N__53067),
            .in1(N__49081),
            .in2(N__49024),
            .in3(N__53087),
            .lcout(\ppm_encoder_1.counter24_0_I_21_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_6_LC_11_2_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_6_LC_11_2_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_6_LC_11_2_1 .LUT_INIT=16'b1111111111101010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_6_LC_11_2_1  (
            .in0(N__53533),
            .in1(N__50981),
            .in2(N__49141),
            .in3(N__49099),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94083),
            .ce(N__50379),
            .sr(N__86505));
    defparam \ppm_encoder_1.pulses2count_esr_7_LC_11_2_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_7_LC_11_2_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_7_LC_11_2_2 .LUT_INIT=16'b0000000000001101;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_7_LC_11_2_2  (
            .in0(N__50982),
            .in1(N__49063),
            .in2(N__53473),
            .in3(N__49042),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94083),
            .ce(N__50379),
            .sr(N__86505));
    defparam \ppm_encoder_1.pulses2count_esr_18_LC_11_2_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_18_LC_11_2_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_18_LC_11_2_3 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_18_LC_11_2_3  (
            .in0(N__49015),
            .in1(N__50979),
            .in2(_gnd_net_),
            .in3(N__49702),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94083),
            .ce(N__50379),
            .sr(N__86505));
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNO_LC_11_2_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNO_LC_11_2_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNO_LC_11_2_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.counter24_0_I_57_c_RNO_LC_11_2_4  (
            .in0(_gnd_net_),
            .in1(N__48988),
            .in2(_gnd_net_),
            .in3(N__53227),
            .lcout(\ppm_encoder_1.counter24_0_I_57_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_8_LC_11_2_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_8_LC_11_2_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_8_LC_11_2_5 .LUT_INIT=16'b0000000001010001;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_8_LC_11_2_5  (
            .in0(N__48976),
            .in1(N__50980),
            .in2(N__48964),
            .in3(N__48916),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94083),
            .ce(N__50379),
            .sr(N__86505));
    defparam \ppm_encoder_1.counter24_0_I_27_c_RNO_LC_11_2_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_27_c_RNO_LC_11_2_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_27_c_RNO_LC_11_2_6 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_27_c_RNO_LC_11_2_6  (
            .in0(N__53012),
            .in1(N__49885),
            .in2(N__49879),
            .in3(N__53036),
            .lcout(\ppm_encoder_1.counter24_0_I_27_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.ppm_output_reg_RNO_0_LC_11_3_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_0_LC_11_3_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_0_LC_11_3_0 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \ppm_encoder_1.ppm_output_reg_RNO_0_LC_11_3_0  (
            .in0(N__53225),
            .in1(N__52939),
            .in2(N__49798),
            .in3(N__49551),
            .lcout(\ppm_encoder_1.N_500 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNI5K08_0_LC_11_3_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNI5K08_0_LC_11_3_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNI5K08_0_LC_11_3_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \ppm_encoder_1.counter_RNI5K08_0_LC_11_3_1  (
            .in0(_gnd_net_),
            .in1(N__52622),
            .in2(_gnd_net_),
            .in3(N__52598),
            .lcout(\ppm_encoder_1.N_486_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIJMMD_LC_11_3_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIJMMD_LC_11_3_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIJMMD_LC_11_3_2 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \ppm_encoder_1.counter24_0_I_57_c_RNIJMMD_LC_11_3_2  (
            .in0(_gnd_net_),
            .in1(N__49563),
            .in2(_gnd_net_),
            .in3(N__49549),
            .lcout(\ppm_encoder_1.counter24_0_I_57_c_RNIJMMDZ0 ),
            .ltout(\ppm_encoder_1.counter24_0_I_57_c_RNIJMMDZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.ppm_output_reg_LC_11_3_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.ppm_output_reg_LC_11_3_3 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.ppm_output_reg_LC_11_3_3 .LUT_INIT=16'b1100110001001111;
    LogicCell40 \ppm_encoder_1.ppm_output_reg_LC_11_3_3  (
            .in0(N__49782),
            .in1(N__49809),
            .in2(N__49831),
            .in3(N__49828),
            .lcout(ppm_output_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94086),
            .ce(),
            .sr(N__86500));
    defparam \ppm_encoder_1.counter_RNI09RH2_18_LC_11_3_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNI09RH2_18_LC_11_3_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNI09RH2_18_LC_11_3_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \ppm_encoder_1.counter_RNI09RH2_18_LC_11_3_4  (
            .in0(N__53224),
            .in1(N__52938),
            .in2(N__49797),
            .in3(N__49781),
            .lcout(\ppm_encoder_1.N_486 ),
            .ltout(\ppm_encoder_1.N_486_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_LC_11_3_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_LC_11_3_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_LC_11_3_5 .LUT_INIT=16'b1111111111110100;
    LogicCell40 \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_LC_11_3_5  (
            .in0(N__49564),
            .in1(N__49552),
            .in2(N__49705),
            .in3(N__71057),
            .lcout(\ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIV9SJ1_LC_11_3_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIV9SJ1_LC_11_3_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIV9SJ1_LC_11_3_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_57_c_RNIV9SJ1_LC_11_3_6  (
            .in0(N__49697),
            .in1(N__49562),
            .in2(N__50598),
            .in3(N__49550),
            .lcout(\ppm_encoder_1.N_374 ),
            .ltout(\ppm_encoder_1.N_374_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_0_LC_11_3_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_0_LC_11_3_7 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_0_LC_11_3_7 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \ppm_encoder_1.init_pulses_0_LC_11_3_7  (
            .in0(N__49394),
            .in1(N__49273),
            .in2(N__49261),
            .in3(N__49258),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94086),
            .ce(),
            .sr(N__86500));
    defparam \ppm_encoder_1.counter24_0_I_1_c_RNO_LC_11_4_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_1_c_RNO_LC_11_4_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_1_c_RNO_LC_11_4_0 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_1_c_RNO_LC_11_4_0  (
            .in0(N__52624),
            .in1(N__50203),
            .in2(N__52603),
            .in3(N__50041),
            .lcout(\ppm_encoder_1.counter24_0_I_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_1_LC_11_4_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_1_LC_11_4_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_1_LC_11_4_2 .LUT_INIT=16'b1111111011101110;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_1_LC_11_4_2  (
            .in0(N__50452),
            .in1(N__50257),
            .in2(N__50245),
            .in3(N__50482),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94091),
            .ce(N__50385),
            .sr(N__86493));
    defparam \ppm_encoder_1.pulses2count_esr_11_LC_11_4_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_11_LC_11_4_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_11_LC_11_4_3 .LUT_INIT=16'b1111111011101110;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_11_LC_11_4_3  (
            .in0(N__50451),
            .in1(N__50197),
            .in2(N__50491),
            .in3(N__50185),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94091),
            .ce(N__50385),
            .sr(N__86493));
    defparam \ppm_encoder_1.counter24_0_I_33_c_RNO_LC_11_4_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_33_c_RNO_LC_11_4_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_33_c_RNO_LC_11_4_4 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_33_c_RNO_LC_11_4_4  (
            .in0(N__50065),
            .in1(N__53417),
            .in2(N__50152),
            .in3(N__52988),
            .lcout(\ppm_encoder_1.counter24_0_I_33_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_10_LC_11_4_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_10_LC_11_4_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_10_LC_11_4_5 .LUT_INIT=16'b0000000001010001;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_10_LC_11_4_5  (
            .in0(N__50134),
            .in1(N__50950),
            .in2(N__50122),
            .in3(N__50077),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94091),
            .ce(N__50385),
            .sr(N__86493));
    defparam \ppm_encoder_1.pulses2count_esr_0_LC_11_5_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_0_LC_11_5_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_0_LC_11_5_0 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_0_LC_11_5_0  (
            .in0(N__53507),
            .in1(N__50059),
            .in2(_gnd_net_),
            .in3(N__50047),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94097),
            .ce(N__50383),
            .sr(N__86490));
    defparam \ppm_encoder_1.pulses2count_esr_4_LC_11_5_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_4_LC_11_5_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_4_LC_11_5_2 .LUT_INIT=16'b0000010100000001;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_4_LC_11_5_2  (
            .in0(N__50035),
            .in1(N__50957),
            .in2(N__50026),
            .in3(N__50017),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94097),
            .ce(N__50383),
            .sr(N__86490));
    defparam \ppm_encoder_1.pulses2count_esr_5_LC_11_5_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_5_LC_11_5_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_5_LC_11_5_6 .LUT_INIT=16'b0000000000001101;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_5_LC_11_5_6  (
            .in0(N__50958),
            .in1(N__49960),
            .in2(N__53818),
            .in3(N__49921),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94097),
            .ce(N__50383),
            .sr(N__86490));
    defparam \ppm_encoder_1.pulses2count_esr_13_LC_11_6_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_13_LC_11_6_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_13_LC_11_6_1 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_13_LC_11_6_1  (
            .in0(N__53517),
            .in1(N__50755),
            .in2(_gnd_net_),
            .in3(N__50743),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94104),
            .ce(N__50386),
            .sr(N__86482));
    defparam \ppm_encoder_1.pulses2count_esr_12_LC_11_6_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_12_LC_11_6_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_12_LC_11_6_2 .LUT_INIT=16'b1111111011101110;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_12_LC_11_6_2  (
            .in0(N__50437),
            .in1(N__50812),
            .in2(N__50497),
            .in3(N__50701),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94104),
            .ce(N__50386),
            .sr(N__86482));
    defparam \ppm_encoder_1.pulses2count_esr_2_LC_11_6_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_2_LC_11_6_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_2_LC_11_6_3 .LUT_INIT=16'b0000000000110001;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_2_LC_11_6_3  (
            .in0(N__50495),
            .in1(N__50659),
            .in2(N__50644),
            .in3(N__50438),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94104),
            .ce(N__50386),
            .sr(N__86482));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_3_LC_11_6_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_3_LC_11_6_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_3_LC_11_6_4 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_3_LC_11_6_4  (
            .in0(N__50611),
            .in1(N__50584),
            .in2(_gnd_net_),
            .in3(N__50530),
            .lcout(),
            .ltout(\ppm_encoder_1.pulses2count_9_0_0_3_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_3_LC_11_6_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_3_LC_11_6_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_3_LC_11_6_5 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_3_LC_11_6_5  (
            .in0(N__50496),
            .in1(N__50439),
            .in2(N__50422),
            .in3(N__50418),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94104),
            .ce(N__50386),
            .sr(N__86482));
    defparam \ppm_encoder_1.counter24_0_I_9_c_RNO_LC_11_6_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_9_c_RNO_LC_11_6_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_9_c_RNO_LC_11_6_6 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_9_c_RNO_LC_11_6_6  (
            .in0(N__53158),
            .in1(N__50317),
            .in2(N__50311),
            .in3(N__52576),
            .lcout(\ppm_encoder_1.counter24_0_I_9_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_7_LC_11_7_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_7_LC_11_7_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_7_LC_11_7_6 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.elevator_7_LC_11_7_6  (
            .in0(N__54571),
            .in1(N__50290),
            .in2(N__51369),
            .in3(N__50280),
            .lcout(\ppm_encoder_1.elevatorZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94110),
            .ce(),
            .sr(N__86473));
    defparam \pid_side.error_i_reg_3_LC_11_8_0 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_3_LC_11_8_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_3_LC_11_8_0 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \pid_side.error_i_reg_3_LC_11_8_0  (
            .in0(N__65485),
            .in1(N__82086),
            .in2(N__62422),
            .in3(N__80722),
            .lcout(\pid_side.error_i_regZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94117),
            .ce(),
            .sr(N__86597));
    defparam \pid_side.state_RNI1OVK_0_LC_11_8_1 .C_ON=1'b0;
    defparam \pid_side.state_RNI1OVK_0_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.state_RNI1OVK_0_LC_11_8_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pid_side.state_RNI1OVK_0_LC_11_8_1  (
            .in0(_gnd_net_),
            .in1(N__65484),
            .in2(_gnd_net_),
            .in3(N__86596),
            .lcout(\pid_side.state_ns_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_13_LC_11_8_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_13_LC_11_8_3 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_13_LC_11_8_3 .LUT_INIT=16'b1101100001110010;
    LogicCell40 \ppm_encoder_1.aileron_13_LC_11_8_3  (
            .in0(N__51327),
            .in1(N__51412),
            .in2(N__51403),
            .in3(N__53931),
            .lcout(\ppm_encoder_1.aileronZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94117),
            .ce(),
            .sr(N__86597));
    defparam \ppm_encoder_1.elevator_5_LC_11_8_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_5_LC_11_8_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_5_LC_11_8_6 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.elevator_5_LC_11_8_6  (
            .in0(N__51385),
            .in1(N__52534),
            .in2(N__51063),
            .in3(N__51328),
            .lcout(\ppm_encoder_1.elevatorZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94117),
            .ce(),
            .sr(N__86597));
    defparam \uart_drone.timer_Count_1_LC_11_9_0 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_1_LC_11_9_0 .SEQ_MODE=4'b1000;
    defparam \uart_drone.timer_Count_1_LC_11_9_0 .LUT_INIT=16'b0100010001000000;
    LogicCell40 \uart_drone.timer_Count_1_LC_11_9_0  (
            .in0(N__70811),
            .in1(N__51043),
            .in2(N__51562),
            .in3(N__50796),
            .lcout(\uart_drone.timer_CountZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94127),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNIU8TV1_3_LC_11_9_3 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNIU8TV1_3_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNIU8TV1_3_LC_11_9_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uart_drone.timer_Count_RNIU8TV1_3_LC_11_9_3  (
            .in0(N__56756),
            .in1(N__51520),
            .in2(_gnd_net_),
            .in3(N__54783),
            .lcout(\uart_drone.N_144_1 ),
            .ltout(\uart_drone.N_144_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_3_LC_11_9_4 .C_ON=1'b0;
    defparam \uart_drone.state_3_LC_11_9_4 .SEQ_MODE=4'b1000;
    defparam \uart_drone.state_3_LC_11_9_4 .LUT_INIT=16'b0000000001000101;
    LogicCell40 \uart_drone.state_3_LC_11_9_4  (
            .in0(N__70810),
            .in1(N__51591),
            .in2(N__51001),
            .in3(N__50998),
            .lcout(\uart_drone.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94127),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_12_LC_11_9_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_12_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_12_LC_11_9_7 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_12_LC_11_9_7  (
            .in0(N__50992),
            .in1(N__50956),
            .in2(N__50869),
            .in3(N__50851),
            .lcout(\ppm_encoder_1.pulses2count_9_0_3_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_4_LC_11_10_0 .C_ON=1'b0;
    defparam \uart_drone.state_4_LC_11_10_0 .SEQ_MODE=4'b1000;
    defparam \uart_drone.state_4_LC_11_10_0 .LUT_INIT=16'b1111001011110000;
    LogicCell40 \uart_drone.state_4_LC_11_10_0  (
            .in0(N__50803),
            .in1(N__70804),
            .in2(N__50797),
            .in3(N__53973),
            .lcout(\uart_drone.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94135),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNO_0_2_LC_11_10_2 .C_ON=1'b0;
    defparam \uart_drone.state_RNO_0_2_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNO_0_2_LC_11_10_2 .LUT_INIT=16'b0000001100100010;
    LogicCell40 \uart_drone.state_RNO_0_2_LC_11_10_2  (
            .in0(N__51590),
            .in1(N__70803),
            .in2(N__56876),
            .in3(N__51440),
            .lcout(),
            .ltout(\uart_drone.state_srsts_i_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_2_LC_11_10_3 .C_ON=1'b0;
    defparam \uart_drone.state_2_LC_11_10_3 .SEQ_MODE=4'b1000;
    defparam \uart_drone.state_2_LC_11_10_3 .LUT_INIT=16'b1011000011110000;
    LogicCell40 \uart_drone.state_2_LC_11_10_3  (
            .in0(N__51441),
            .in1(N__51518),
            .in2(N__51634),
            .in3(N__54775),
            .lcout(\uart_drone.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94135),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIRSI31_11_LC_11_10_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIRSI31_11_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIRSI31_11_LC_11_10_4 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \Commands_frame_decoder.state_RNIRSI31_11_LC_11_10_4  (
            .in0(N__51631),
            .in1(N__70802),
            .in2(_gnd_net_),
            .in3(N__55253),
            .lcout(\Commands_frame_decoder.state_RNIRSI31Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNI40411_2_LC_11_10_5 .C_ON=1'b0;
    defparam \uart_drone.state_RNI40411_2_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNI40411_2_LC_11_10_5 .LUT_INIT=16'b0101010011111100;
    LogicCell40 \uart_drone.state_RNI40411_2_LC_11_10_5  (
            .in0(N__51514),
            .in1(N__51589),
            .in2(N__53984),
            .in3(N__54774),
            .lcout(\uart_drone.timer_Count_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNI62411_4_LC_11_10_7 .C_ON=1'b0;
    defparam \uart_drone.state_RNI62411_4_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNI62411_4_LC_11_10_7 .LUT_INIT=16'b0010001100000011;
    LogicCell40 \uart_drone.state_RNI62411_4_LC_11_10_7  (
            .in0(N__51513),
            .in1(N__54812),
            .in2(N__53983),
            .in3(N__54773),
            .lcout(\uart_drone.un1_state_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_1_LC_11_11_0 .C_ON=1'b0;
    defparam \uart_drone.state_1_LC_11_11_0 .SEQ_MODE=4'b1000;
    defparam \uart_drone.state_1_LC_11_11_0 .LUT_INIT=16'b0000000011001000;
    LogicCell40 \uart_drone.state_1_LC_11_11_0  (
            .in0(N__51445),
            .in1(N__56827),
            .in2(N__54709),
            .in3(N__70753),
            .lcout(\uart_drone.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94142),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNIP8RT_10_LC_11_11_1 .C_ON=1'b0;
    defparam \reset_module_System.count_RNIP8RT_10_LC_11_11_1 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNIP8RT_10_LC_11_11_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \reset_module_System.count_RNIP8RT_10_LC_11_11_1  (
            .in0(_gnd_net_),
            .in1(N__51877),
            .in2(_gnd_net_),
            .in3(N__51895),
            .lcout(\reset_module_System.reset6_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone_sync.aux_3__0__0_LC_11_11_2 .C_ON=1'b0;
    defparam \uart_drone_sync.aux_3__0__0_LC_11_11_2 .SEQ_MODE=4'b1000;
    defparam \uart_drone_sync.aux_3__0__0_LC_11_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone_sync.aux_3__0__0_LC_11_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51427),
            .lcout(\uart_drone_sync.aux_3__0__0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94142),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone_sync.Q_0__0_LC_11_11_3 .C_ON=1'b0;
    defparam \uart_drone_sync.Q_0__0_LC_11_11_3 .SEQ_MODE=4'b1000;
    defparam \uart_drone_sync.Q_0__0_LC_11_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone_sync.Q_0__0_LC_11_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51418),
            .lcout(debug_CH0_16A_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94142),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_6_LC_11_11_5 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_6_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_6_LC_11_11_5 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \uart_drone.data_Aux_RNO_0_6_LC_11_11_5  (
            .in0(N__56493),
            .in1(N__56556),
            .in2(_gnd_net_),
            .in3(N__56622),
            .lcout(\uart_drone.data_Auxce_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNI9ADK1_4_LC_11_11_6 .C_ON=1'b0;
    defparam \uart_drone.state_RNI9ADK1_4_LC_11_11_6 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNI9ADK1_4_LC_11_11_6 .LUT_INIT=16'b1111111100101010;
    LogicCell40 \uart_drone.state_RNI9ADK1_4_LC_11_11_6  (
            .in0(N__53985),
            .in1(N__54723),
            .in2(N__51670),
            .in3(N__54813),
            .lcout(\uart_drone.un1_state_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_4_LC_11_11_7 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_4_LC_11_11_7 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_4_LC_11_11_7 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \uart_drone.data_Aux_RNO_0_4_LC_11_11_7  (
            .in0(N__56492),
            .in1(N__56555),
            .in2(_gnd_net_),
            .in3(N__56621),
            .lcout(\uart_drone.data_Auxce_0_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_0_LC_11_12_0 .C_ON=1'b0;
    defparam \reset_module_System.count_0_LC_11_12_0 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_0_LC_11_12_0 .LUT_INIT=16'b1101010101010101;
    LogicCell40 \reset_module_System.count_0_LC_11_12_0  (
            .in0(N__51777),
            .in1(N__55029),
            .in2(N__54945),
            .in3(N__54919),
            .lcout(\reset_module_System.countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94155),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNI10J41_1_LC_11_12_1 .C_ON=1'b0;
    defparam \reset_module_System.count_RNI10J41_1_LC_11_12_1 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNI10J41_1_LC_11_12_1 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \reset_module_System.count_RNI10J41_1_LC_11_12_1  (
            .in0(N__51730),
            .in1(N__51973),
            .in2(N__51814),
            .in3(N__51752),
            .lcout(\reset_module_System.reset6_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNO_0_1_LC_11_12_2 .C_ON=1'b0;
    defparam \reset_module_System.count_RNO_0_1_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNO_0_1_LC_11_12_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \reset_module_System.count_RNO_0_1_LC_11_12_2  (
            .in0(N__51753),
            .in1(_gnd_net_),
            .in2(N__51778),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\reset_module_System.count_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_1_LC_11_12_3 .C_ON=1'b0;
    defparam \reset_module_System.count_1_LC_11_12_3 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_1_LC_11_12_3 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \reset_module_System.count_1_LC_11_12_3  (
            .in0(N__55030),
            .in1(N__54916),
            .in2(N__51661),
            .in3(N__54940),
            .lcout(\reset_module_System.countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94155),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNIN3HK3_12_LC_11_12_4 .C_ON=1'b0;
    defparam \reset_module_System.count_RNIN3HK3_12_LC_11_12_4 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNIN3HK3_12_LC_11_12_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \reset_module_System.count_RNIN3HK3_12_LC_11_12_4  (
            .in0(N__51773),
            .in1(N__54835),
            .in2(N__51859),
            .in3(N__51784),
            .lcout(\reset_module_System.reset6_19 ),
            .ltout(\reset_module_System.reset6_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.reset_iso_LC_11_12_5 .C_ON=1'b0;
    defparam \reset_module_System.reset_iso_LC_11_12_5 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.reset_iso_LC_11_12_5 .LUT_INIT=16'b0101111111111111;
    LogicCell40 \reset_module_System.reset_iso_LC_11_12_5  (
            .in0(N__55028),
            .in1(_gnd_net_),
            .in2(N__51658),
            .in3(N__54936),
            .lcout(\reset_module_System.reset_isoZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94155),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNI97FD_5_LC_11_12_6 .C_ON=1'b0;
    defparam \reset_module_System.count_RNI97FD_5_LC_11_12_6 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNI97FD_5_LC_11_12_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \reset_module_System.count_RNI97FD_5_LC_11_12_6  (
            .in0(N__51714),
            .in1(N__51681),
            .in2(N__51916),
            .in3(N__51696),
            .lcout(),
            .ltout(\reset_module_System.reset6_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNI53692_14_LC_11_12_7 .C_ON=1'b0;
    defparam \reset_module_System.count_RNI53692_14_LC_11_12_7 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNI53692_14_LC_11_12_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \reset_module_System.count_RNI53692_14_LC_11_12_7  (
            .in0(N__51991),
            .in1(N__51835),
            .in2(N__51793),
            .in3(N__51790),
            .lcout(\reset_module_System.reset6_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_1_cry_1_c_LC_11_13_0 .C_ON=1'b1;
    defparam \reset_module_System.count_1_cry_1_c_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_1_cry_1_c_LC_11_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \reset_module_System.count_1_cry_1_c_LC_11_13_0  (
            .in0(_gnd_net_),
            .in1(N__51772),
            .in2(N__51757),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_13_0_),
            .carryout(\reset_module_System.count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNO_0_2_LC_11_13_1 .C_ON=1'b1;
    defparam \reset_module_System.count_RNO_0_2_LC_11_13_1 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNO_0_2_LC_11_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_RNO_0_2_LC_11_13_1  (
            .in0(_gnd_net_),
            .in1(N__54849),
            .in2(_gnd_net_),
            .in3(N__51736),
            .lcout(\reset_module_System.count_1_2 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_1 ),
            .carryout(\reset_module_System.count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_3_LC_11_13_2 .C_ON=1'b1;
    defparam \reset_module_System.count_3_LC_11_13_2 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_3_LC_11_13_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_3_LC_11_13_2  (
            .in0(_gnd_net_),
            .in1(N__54883),
            .in2(_gnd_net_),
            .in3(N__51733),
            .lcout(\reset_module_System.countZ0Z_3 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_2 ),
            .carryout(\reset_module_System.count_1_cry_3 ),
            .clk(N__94167),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_4_LC_11_13_3 .C_ON=1'b1;
    defparam \reset_module_System.count_4_LC_11_13_3 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_4_LC_11_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_4_LC_11_13_3  (
            .in0(_gnd_net_),
            .in1(N__51729),
            .in2(_gnd_net_),
            .in3(N__51718),
            .lcout(\reset_module_System.countZ0Z_4 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_3 ),
            .carryout(\reset_module_System.count_1_cry_4 ),
            .clk(N__94167),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_5_LC_11_13_4 .C_ON=1'b1;
    defparam \reset_module_System.count_5_LC_11_13_4 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_5_LC_11_13_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_5_LC_11_13_4  (
            .in0(_gnd_net_),
            .in1(N__51715),
            .in2(_gnd_net_),
            .in3(N__51703),
            .lcout(\reset_module_System.countZ0Z_5 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_4 ),
            .carryout(\reset_module_System.count_1_cry_5 ),
            .clk(N__94167),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_6_LC_11_13_5 .C_ON=1'b1;
    defparam \reset_module_System.count_6_LC_11_13_5 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_6_LC_11_13_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_6_LC_11_13_5  (
            .in0(_gnd_net_),
            .in1(N__54897),
            .in2(_gnd_net_),
            .in3(N__51700),
            .lcout(\reset_module_System.countZ0Z_6 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_5 ),
            .carryout(\reset_module_System.count_1_cry_6 ),
            .clk(N__94167),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_7_LC_11_13_6 .C_ON=1'b1;
    defparam \reset_module_System.count_7_LC_11_13_6 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_7_LC_11_13_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_7_LC_11_13_6  (
            .in0(_gnd_net_),
            .in1(N__51697),
            .in2(_gnd_net_),
            .in3(N__51685),
            .lcout(\reset_module_System.countZ0Z_7 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_6 ),
            .carryout(\reset_module_System.count_1_cry_7 ),
            .clk(N__94167),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_8_LC_11_13_7 .C_ON=1'b1;
    defparam \reset_module_System.count_8_LC_11_13_7 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_8_LC_11_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_8_LC_11_13_7  (
            .in0(_gnd_net_),
            .in1(N__51682),
            .in2(_gnd_net_),
            .in3(N__51919),
            .lcout(\reset_module_System.countZ0Z_8 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_7 ),
            .carryout(\reset_module_System.count_1_cry_8 ),
            .clk(N__94167),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_9_LC_11_14_0 .C_ON=1'b1;
    defparam \reset_module_System.count_9_LC_11_14_0 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_9_LC_11_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_9_LC_11_14_0  (
            .in0(_gnd_net_),
            .in1(N__51912),
            .in2(_gnd_net_),
            .in3(N__51898),
            .lcout(\reset_module_System.countZ0Z_9 ),
            .ltout(),
            .carryin(bfn_11_14_0_),
            .carryout(\reset_module_System.count_1_cry_9 ),
            .clk(N__94180),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_10_LC_11_14_1 .C_ON=1'b1;
    defparam \reset_module_System.count_10_LC_11_14_1 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_10_LC_11_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_10_LC_11_14_1  (
            .in0(_gnd_net_),
            .in1(N__51894),
            .in2(_gnd_net_),
            .in3(N__51880),
            .lcout(\reset_module_System.countZ0Z_10 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_9 ),
            .carryout(\reset_module_System.count_1_cry_10 ),
            .clk(N__94180),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_11_LC_11_14_2 .C_ON=1'b1;
    defparam \reset_module_System.count_11_LC_11_14_2 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_11_LC_11_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_11_LC_11_14_2  (
            .in0(_gnd_net_),
            .in1(N__51876),
            .in2(_gnd_net_),
            .in3(N__51862),
            .lcout(\reset_module_System.countZ0Z_11 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_10 ),
            .carryout(\reset_module_System.count_1_cry_11 ),
            .clk(N__94180),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_12_LC_11_14_3 .C_ON=1'b1;
    defparam \reset_module_System.count_12_LC_11_14_3 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_12_LC_11_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_12_LC_11_14_3  (
            .in0(_gnd_net_),
            .in1(N__51852),
            .in2(_gnd_net_),
            .in3(N__51841),
            .lcout(\reset_module_System.countZ0Z_12 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_11 ),
            .carryout(\reset_module_System.count_1_cry_12 ),
            .clk(N__94180),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_13_LC_11_14_4 .C_ON=1'b1;
    defparam \reset_module_System.count_13_LC_11_14_4 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_13_LC_11_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_13_LC_11_14_4  (
            .in0(_gnd_net_),
            .in1(N__55041),
            .in2(_gnd_net_),
            .in3(N__51838),
            .lcout(\reset_module_System.countZ0Z_13 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_12 ),
            .carryout(\reset_module_System.count_1_cry_13 ),
            .clk(N__94180),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_14_LC_11_14_5 .C_ON=1'b1;
    defparam \reset_module_System.count_14_LC_11_14_5 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_14_LC_11_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_14_LC_11_14_5  (
            .in0(_gnd_net_),
            .in1(N__51834),
            .in2(_gnd_net_),
            .in3(N__51820),
            .lcout(\reset_module_System.countZ0Z_14 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_13 ),
            .carryout(\reset_module_System.count_1_cry_14 ),
            .clk(N__94180),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_15_LC_11_14_6 .C_ON=1'b1;
    defparam \reset_module_System.count_15_LC_11_14_6 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_15_LC_11_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_15_LC_11_14_6  (
            .in0(_gnd_net_),
            .in1(N__55068),
            .in2(_gnd_net_),
            .in3(N__51817),
            .lcout(\reset_module_System.countZ0Z_15 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_14 ),
            .carryout(\reset_module_System.count_1_cry_15 ),
            .clk(N__94180),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_16_LC_11_14_7 .C_ON=1'b1;
    defparam \reset_module_System.count_16_LC_11_14_7 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_16_LC_11_14_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_16_LC_11_14_7  (
            .in0(_gnd_net_),
            .in1(N__51807),
            .in2(_gnd_net_),
            .in3(N__51796),
            .lcout(\reset_module_System.countZ0Z_16 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_15 ),
            .carryout(\reset_module_System.count_1_cry_16 ),
            .clk(N__94180),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_17_LC_11_15_0 .C_ON=1'b1;
    defparam \reset_module_System.count_17_LC_11_15_0 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_17_LC_11_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_17_LC_11_15_0  (
            .in0(_gnd_net_),
            .in1(N__51990),
            .in2(_gnd_net_),
            .in3(N__51976),
            .lcout(\reset_module_System.countZ0Z_17 ),
            .ltout(),
            .carryin(bfn_11_15_0_),
            .carryout(\reset_module_System.count_1_cry_17 ),
            .clk(N__94193),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_18_LC_11_15_1 .C_ON=1'b1;
    defparam \reset_module_System.count_18_LC_11_15_1 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_18_LC_11_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_18_LC_11_15_1  (
            .in0(_gnd_net_),
            .in1(N__51972),
            .in2(_gnd_net_),
            .in3(N__51958),
            .lcout(\reset_module_System.countZ0Z_18 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_17 ),
            .carryout(\reset_module_System.count_1_cry_18 ),
            .clk(N__94193),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_19_LC_11_15_2 .C_ON=1'b1;
    defparam \reset_module_System.count_19_LC_11_15_2 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_19_LC_11_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_19_LC_11_15_2  (
            .in0(_gnd_net_),
            .in1(N__55081),
            .in2(_gnd_net_),
            .in3(N__51955),
            .lcout(\reset_module_System.countZ0Z_19 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_18 ),
            .carryout(\reset_module_System.count_1_cry_19 ),
            .clk(N__94193),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_20_LC_11_15_3 .C_ON=1'b1;
    defparam \reset_module_System.count_20_LC_11_15_3 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_20_LC_11_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_20_LC_11_15_3  (
            .in0(_gnd_net_),
            .in1(N__54864),
            .in2(_gnd_net_),
            .in3(N__51952),
            .lcout(\reset_module_System.countZ0Z_20 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_19 ),
            .carryout(\reset_module_System.count_1_cry_20 ),
            .clk(N__94193),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_21_LC_11_15_4 .C_ON=1'b0;
    defparam \reset_module_System.count_21_LC_11_15_4 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_21_LC_11_15_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \reset_module_System.count_21_LC_11_15_4  (
            .in0(_gnd_net_),
            .in1(N__55056),
            .in2(_gnd_net_),
            .in3(N__51949),
            .lcout(\reset_module_System.countZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94193),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIJ9P4_7_LC_11_15_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIJ9P4_7_LC_11_15_5 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIJ9P4_7_LC_11_15_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_RNIJ9P4_7_LC_11_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51946),
            .lcout(drone_H_disp_side_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIHL1J_5_LC_11_15_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIHL1J_5_LC_11_15_7 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIHL1J_5_LC_11_15_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_RNIHL1J_5_LC_11_15_7  (
            .in0(_gnd_net_),
            .in1(N__69343),
            .in2(_gnd_net_),
            .in3(N__55234),
            .lcout(\Commands_frame_decoder.source_CH4data_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_10_LC_11_16_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_10_LC_11_16_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_10_LC_11_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_10_LC_11_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57244),
            .lcout(\dron_frame_decoder_1.drone_H_disp_side_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94209),
            .ce(N__52264),
            .sr(N__86433));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_11_LC_11_16_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_11_LC_11_16_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_11_LC_11_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_11_LC_11_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58016),
            .lcout(drone_H_disp_side_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94209),
            .ce(N__52264),
            .sr(N__86433));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_12_LC_11_16_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_12_LC_11_16_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_12_LC_11_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_12_LC_11_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57938),
            .lcout(drone_H_disp_side_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94209),
            .ce(N__52264),
            .sr(N__86433));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_13_LC_11_16_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_13_LC_11_16_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_13_LC_11_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_13_LC_11_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57868),
            .lcout(drone_H_disp_side_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94209),
            .ce(N__52264),
            .sr(N__86433));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_14_LC_11_16_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_14_LC_11_16_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_14_LC_11_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_14_LC_11_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57137),
            .lcout(drone_H_disp_side_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94209),
            .ce(N__52264),
            .sr(N__86433));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_15_LC_11_16_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_15_LC_11_16_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_15_LC_11_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_15_LC_11_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57792),
            .lcout(drone_H_disp_side_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94209),
            .ce(N__52264),
            .sr(N__86433));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_8_LC_11_16_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_8_LC_11_16_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_8_LC_11_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_8_LC_11_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57722),
            .lcout(\dron_frame_decoder_1.drone_H_disp_side_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94209),
            .ce(N__52264),
            .sr(N__86433));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_9_LC_11_16_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_9_LC_11_16_7 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_9_LC_11_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_9_LC_11_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57317),
            .lcout(\dron_frame_decoder_1.drone_H_disp_side_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94209),
            .ce(N__52264),
            .sr(N__86433));
    defparam \uart_pc.data_rdy_LC_11_17_1 .C_ON=1'b0;
    defparam \uart_pc.data_rdy_LC_11_17_1 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_rdy_LC_11_17_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uart_pc.data_rdy_LC_11_17_1  (
            .in0(N__52230),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52132),
            .lcout(uart_pc_data_rdy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94226),
            .ce(),
            .sr(N__86425));
    defparam \Commands_frame_decoder.source_alt_kp_4_LC_11_17_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_4_LC_11_17_2 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_alt_kp_4_LC_11_17_2 .LUT_INIT=16'b1011111110000000;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_4_LC_11_17_2  (
            .in0(N__88829),
            .in1(N__52108),
            .in2(N__55208),
            .in3(N__52071),
            .lcout(alt_kp_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94226),
            .ce(),
            .sr(N__86425));
    defparam \Commands_frame_decoder.source_xy_kp_4_LC_11_17_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kp_4_LC_11_17_3 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_xy_kp_4_LC_11_17_3 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \Commands_frame_decoder.source_xy_kp_4_LC_11_17_3  (
            .in0(N__52010),
            .in1(N__55158),
            .in2(N__52057),
            .in3(N__88830),
            .lcout(xy_kp_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94226),
            .ce(),
            .sr(N__86425));
    defparam \Commands_frame_decoder.state_3_LC_11_17_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_3_LC_11_17_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_3_LC_11_17_5 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \Commands_frame_decoder.state_3_LC_11_17_5  (
            .in0(N__52419),
            .in1(N__52457),
            .in2(_gnd_net_),
            .in3(N__69392),
            .lcout(\Commands_frame_decoder.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94226),
            .ce(),
            .sr(N__86425));
    defparam \Commands_frame_decoder.state_4_LC_11_17_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_4_LC_11_17_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_4_LC_11_17_6 .LUT_INIT=16'b1111111110100000;
    LogicCell40 \Commands_frame_decoder.state_4_LC_11_17_6  (
            .in0(N__69393),
            .in1(_gnd_net_),
            .in2(N__52384),
            .in3(N__52405),
            .lcout(\Commands_frame_decoder.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94226),
            .ce(),
            .sr(N__86425));
    defparam \Commands_frame_decoder.state_RNIGK1J_4_LC_11_17_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIGK1J_4_LC_11_17_7 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIGK1J_4_LC_11_17_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_RNIGK1J_4_LC_11_17_7  (
            .in0(_gnd_net_),
            .in1(N__52380),
            .in2(_gnd_net_),
            .in3(N__55157),
            .lcout(\Commands_frame_decoder.source_CH3data_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_axb_13_LC_11_18_0 .C_ON=1'b0;
    defparam \pid_alt.error_axb_13_LC_11_18_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_axb_13_LC_11_18_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_axb_13_LC_11_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52357),
            .lcout(\pid_alt.error_axbZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_13_LC_11_18_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_13_LC_11_18_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_13_LC_11_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_13_LC_11_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57872),
            .lcout(drone_altitude_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94243),
            .ce(N__52330),
            .sr(N__86414));
    defparam \pid_alt.error_axb_14_LC_11_18_2 .C_ON=1'b0;
    defparam \pid_alt.error_axb_14_LC_11_18_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_axb_14_LC_11_18_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_axb_14_LC_11_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52336),
            .lcout(\pid_alt.error_axbZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_14_LC_11_18_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_14_LC_11_18_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_14_LC_11_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_14_LC_11_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57147),
            .lcout(drone_altitude_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94243),
            .ce(N__52330),
            .sr(N__86414));
    defparam \pid_alt.error_axb_2_LC_11_18_4 .C_ON=1'b0;
    defparam \pid_alt.error_axb_2_LC_11_18_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_axb_2_LC_11_18_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_axb_2_LC_11_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52306),
            .lcout(\pid_alt.error_axbZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_axb_3_LC_11_18_5 .C_ON=1'b0;
    defparam \pid_alt.error_axb_3_LC_11_18_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_axb_3_LC_11_18_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_axb_3_LC_11_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52291),
            .lcout(\pid_alt.error_axbZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_axb_1_LC_11_18_6 .C_ON=1'b0;
    defparam \pid_front.error_axb_1_LC_11_18_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_axb_1_LC_11_18_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_front.error_axb_1_LC_11_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52495),
            .lcout(\pid_front.error_axbZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_axb_2_LC_11_18_7 .C_ON=1'b0;
    defparam \pid_front.error_axb_2_LC_11_18_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_axb_2_LC_11_18_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_front.error_axb_2_LC_11_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55363),
            .lcout(\pid_front.error_axbZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_0_LC_11_19_0 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_0_LC_11_19_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_0_LC_11_19_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_0_LC_11_19_0  (
            .in0(_gnd_net_),
            .in1(N__66289),
            .in2(_gnd_net_),
            .in3(N__66373),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94260),
            .ce(N__75321),
            .sr(N__86403));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIVIR9_11_LC_11_19_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIVIR9_11_LC_11_19_2 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIVIR9_11_LC_11_19_2 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNIVIR9_11_LC_11_19_2  (
            .in0(_gnd_net_),
            .in1(N__52489),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(drone_altitude_i_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNI1A23_10_LC_11_19_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNI1A23_10_LC_11_19_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNI1A23_10_LC_11_19_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_RNI1A23_10_LC_11_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55570),
            .lcout(drone_H_disp_front_i_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNI4D23_13_LC_11_19_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNI4D23_13_LC_11_19_4 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNI4D23_13_LC_11_19_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_RNI4D23_13_LC_11_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57814),
            .lcout(drone_H_disp_front_i_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIK7V3_4_LC_11_19_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIK7V3_4_LC_11_19_5 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIK7V3_4_LC_11_19_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_RNIK7V3_4_LC_11_19_5  (
            .in0(N__55357),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(drone_H_disp_front_i_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIL8V3_5_LC_11_19_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIL8V3_5_LC_11_19_6 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIL8V3_5_LC_11_19_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_RNIL8V3_5_LC_11_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52471),
            .lcout(drone_H_disp_front_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIM9V3_6_LC_11_19_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIM9V3_6_LC_11_19_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIM9V3_6_LC_11_19_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_RNIM9V3_6_LC_11_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52501),
            .lcout(drone_H_disp_front_i_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_5_LC_11_20_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_5_LC_11_20_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_5_LC_11_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_5_LC_11_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57873),
            .lcout(\dron_frame_decoder_1.drone_H_disp_front_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94279),
            .ce(N__57399),
            .sr(N__86394));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_6_LC_11_20_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_6_LC_11_20_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_6_LC_11_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_6_LC_11_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57149),
            .lcout(\dron_frame_decoder_1.drone_H_disp_front_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94279),
            .ce(N__57399),
            .sr(N__86394));
    defparam \pid_front.error_i_acumm_13_LC_11_21_0 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_13_LC_11_21_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_13_LC_11_21_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_front.error_i_acumm_13_LC_11_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70117),
            .lcout(\pid_front.error_i_acummZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94294),
            .ce(N__75769),
            .sr(_gnd_net_));
    defparam \pid_front.un11lto30_i_a2_0_c_LC_11_22_0 .C_ON=1'b1;
    defparam \pid_front.un11lto30_i_a2_0_c_LC_11_22_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.un11lto30_i_a2_0_c_LC_11_22_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_front.un11lto30_i_a2_0_c_LC_11_22_0  (
            .in0(_gnd_net_),
            .in1(N__58057),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_22_0_),
            .carryout(\pid_front.un11lto30_i_a2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un11lto30_i_a2_1_c_LC_11_22_1 .C_ON=1'b1;
    defparam \pid_front.un11lto30_i_a2_1_c_LC_11_22_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.un11lto30_i_a2_1_c_LC_11_22_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_front.un11lto30_i_a2_1_c_LC_11_22_1  (
            .in0(_gnd_net_),
            .in1(N__52546),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_front.un11lto30_i_a2 ),
            .carryout(\pid_front.un11lto30_i_a2_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un11lto30_i_a2_2_c_LC_11_22_2 .C_ON=1'b1;
    defparam \pid_front.un11lto30_i_a2_2_c_LC_11_22_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.un11lto30_i_a2_2_c_LC_11_22_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_front.un11lto30_i_a2_2_c_LC_11_22_2  (
            .in0(_gnd_net_),
            .in1(N__52510),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_front.un11lto30_i_a2_0 ),
            .carryout(\pid_front.un11lto30_i_a2_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un11lto30_i_a2_3_c_LC_11_22_3 .C_ON=1'b1;
    defparam \pid_front.un11lto30_i_a2_3_c_LC_11_22_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.un11lto30_i_a2_3_c_LC_11_22_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_front.un11lto30_i_a2_3_c_LC_11_22_3  (
            .in0(_gnd_net_),
            .in1(N__55807),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_front.un11lto30_i_a2_1 ),
            .carryout(\pid_front.un11lto30_i_a2_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un11lto30_i_a2_4_c_LC_11_22_4 .C_ON=1'b1;
    defparam \pid_front.un11lto30_i_a2_4_c_LC_11_22_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.un11lto30_i_a2_4_c_LC_11_22_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_front.un11lto30_i_a2_4_c_LC_11_22_4  (
            .in0(_gnd_net_),
            .in1(N__55828),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_front.un11lto30_i_a2_2 ),
            .carryout(\pid_front.un11lto30_i_a2_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un11lto30_i_a2_5_c_LC_11_22_5 .C_ON=1'b1;
    defparam \pid_front.un11lto30_i_a2_5_c_LC_11_22_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.un11lto30_i_a2_5_c_LC_11_22_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_front.un11lto30_i_a2_5_c_LC_11_22_5  (
            .in0(_gnd_net_),
            .in1(N__55557),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_front.un11lto30_i_a2_3 ),
            .carryout(\pid_front.un11lto30_i_a2_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un11lto30_i_a2_6_c_LC_11_22_6 .C_ON=1'b1;
    defparam \pid_front.un11lto30_i_a2_6_c_LC_11_22_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.un11lto30_i_a2_6_c_LC_11_22_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_front.un11lto30_i_a2_6_c_LC_11_22_6  (
            .in0(_gnd_net_),
            .in1(N__55927),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_front.un11lto30_i_a2_4 ),
            .carryout(\pid_front.un11lto30_i_a2_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un11lto30_i_a2_7_c_LC_11_22_7 .C_ON=1'b1;
    defparam \pid_front.un11lto30_i_a2_7_c_LC_11_22_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.un11lto30_i_a2_7_c_LC_11_22_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_front.un11lto30_i_a2_7_c_LC_11_22_7  (
            .in0(_gnd_net_),
            .in1(N__55852),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_front.un11lto30_i_a2_5 ),
            .carryout(\pid_front.un11lto30_i_a2_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un11lto30_i_a2_7_c_RNIQ1JH6_LC_11_23_0 .C_ON=1'b0;
    defparam \pid_front.un11lto30_i_a2_7_c_RNIQ1JH6_LC_11_23_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.un11lto30_i_a2_7_c_RNIQ1JH6_LC_11_23_0 .LUT_INIT=16'b1110111011111111;
    LogicCell40 \pid_front.un11lto30_i_a2_7_c_RNIQ1JH6_LC_11_23_0  (
            .in0(N__55777),
            .in1(N__55764),
            .in2(_gnd_net_),
            .in3(N__52549),
            .lcout(\pid_front.N_291 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNI3Q532_4_LC_11_23_2 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNI3Q532_4_LC_11_23_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNI3Q532_4_LC_11_23_2 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \pid_front.pid_prereg_esr_RNI3Q532_4_LC_11_23_2  (
            .in0(N__58464),
            .in1(N__58866),
            .in2(N__55537),
            .in3(N__58431),
            .lcout(\pid_front.N_631 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un11lto30_i_a2_1_c_RNO_LC_11_23_3 .C_ON=1'b0;
    defparam \pid_front.un11lto30_i_a2_1_c_RNO_LC_11_23_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.un11lto30_i_a2_1_c_RNO_LC_11_23_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_front.un11lto30_i_a2_1_c_RNO_LC_11_23_3  (
            .in0(N__58430),
            .in1(N__58394),
            .in2(N__58368),
            .in3(N__58463),
            .lcout(\pid_front.un11lto30_i_a2_0_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNI211A1_20_LC_11_24_0 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNI211A1_20_LC_11_24_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNI211A1_20_LC_11_24_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_front.pid_prereg_esr_RNI211A1_20_LC_11_24_0  (
            .in0(N__58750),
            .in1(N__58726),
            .in2(N__58711),
            .in3(N__58783),
            .lcout(\pid_front.un11lto30_i_a2_4_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNIRM2N_6_LC_11_24_1 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNIRM2N_6_LC_11_24_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNIRM2N_6_LC_11_24_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_front.pid_prereg_esr_RNIRM2N_6_LC_11_24_1  (
            .in0(N__58200),
            .in1(N__58230),
            .in2(N__58364),
            .in3(N__58401),
            .lcout(),
            .ltout(\pid_front.un1_reset_i_a2_3_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNIOL7G1_8_LC_11_24_2 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNIOL7G1_8_LC_11_24_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNIOL7G1_8_LC_11_24_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_front.pid_prereg_esr_RNIOL7G1_8_LC_11_24_2  (
            .in0(N__58284),
            .in1(N__58649),
            .in2(N__52540),
            .in3(N__58578),
            .lcout(\pid_front.N_593 ),
            .ltout(\pid_front.N_593_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.source_pid_1_esr_5_LC_11_24_3 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_esr_5_LC_11_24_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_esr_5_LC_11_24_3 .LUT_INIT=16'b0100010100000000;
    LogicCell40 \pid_front.source_pid_1_esr_5_LC_11_24_3  (
            .in0(N__60149),
            .in1(N__58872),
            .in2(N__52537),
            .in3(N__58435),
            .lcout(front_order_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94342),
            .ce(N__60029),
            .sr(N__59971));
    defparam \pid_front.un11lto30_i_a2_2_c_RNO_LC_11_24_5 .C_ON=1'b0;
    defparam \pid_front.un11lto30_i_a2_2_c_RNO_LC_11_24_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.un11lto30_i_a2_2_c_RNO_LC_11_24_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_front.un11lto30_i_a2_2_c_RNO_LC_11_24_5  (
            .in0(N__58199),
            .in1(N__58229),
            .in2(N__58653),
            .in3(N__58283),
            .lcout(\pid_front.N_11_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_45_c_RNO_LC_12_1_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_45_c_RNO_LC_12_1_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_45_c_RNO_LC_12_1_0 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_45_c_RNO_LC_12_1_0  (
            .in0(N__53313),
            .in1(N__52969),
            .in2(N__52963),
            .in3(N__53334),
            .lcout(\ppm_encoder_1.counter24_0_I_45_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNIS9KG_8_LC_12_1_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNIS9KG_8_LC_12_1_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNIS9KG_8_LC_12_1_1 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \ppm_encoder_1.counter_RNIS9KG_8_LC_12_1_1  (
            .in0(N__52993),
            .in1(N__53017),
            .in2(N__53425),
            .in3(N__53041),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_a2_18_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNIG7H22_2_LC_12_1_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNIG7H22_2_LC_12_1_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNIG7H22_2_LC_12_1_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ppm_encoder_1.counter_RNIG7H22_2_LC_12_1_2  (
            .in0(N__52912),
            .in1(N__52918),
            .in2(N__52942),
            .in3(N__52924),
            .lcout(\ppm_encoder_1.N_486_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNIS9KG_2_LC_12_1_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNIS9KG_2_LC_12_1_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNIS9KG_2_LC_12_1_3 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \ppm_encoder_1.counter_RNIS9KG_2_LC_12_1_3  (
            .in0(N__53293),
            .in1(N__53153),
            .in2(N__53263),
            .in3(N__52571),
            .lcout(\ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_a2_18_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNIQM6H_12_LC_12_1_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNIQM6H_12_LC_12_1_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNIQM6H_12_LC_12_1_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \ppm_encoder_1.counter_RNIQM6H_12_LC_12_1_4  (
            .in0(N__53314),
            .in1(N__53364),
            .in2(N__53398),
            .in3(N__53335),
            .lcout(\ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_a2_18_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNIUS1G_4_LC_12_1_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNIUS1G_4_LC_12_1_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNIUS1G_4_LC_12_1_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \ppm_encoder_1.counter_RNIUS1G_4_LC_12_1_5  (
            .in0(N__53088),
            .in1(N__53109),
            .in2(N__53068),
            .in3(N__53130),
            .lcout(\ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_a2_18_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_0_LC_12_2_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_0_LC_12_2_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_0_LC_12_2_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_0_LC_12_2_0  (
            .in0(_gnd_net_),
            .in1(N__52623),
            .in2(N__52905),
            .in3(N__52899),
            .lcout(\ppm_encoder_1.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_12_2_0_),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_0 ),
            .clk(N__94081),
            .ce(),
            .sr(N__53202));
    defparam \ppm_encoder_1.counter_1_LC_12_2_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_1_LC_12_2_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_1_LC_12_2_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_1_LC_12_2_1  (
            .in0(_gnd_net_),
            .in1(N__52599),
            .in2(_gnd_net_),
            .in3(N__52579),
            .lcout(\ppm_encoder_1.counterZ0Z_1 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_0 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_1 ),
            .clk(N__94081),
            .ce(),
            .sr(N__53202));
    defparam \ppm_encoder_1.counter_2_LC_12_2_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_2_LC_12_2_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_2_LC_12_2_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_2_LC_12_2_2  (
            .in0(_gnd_net_),
            .in1(N__52575),
            .in2(_gnd_net_),
            .in3(N__52552),
            .lcout(\ppm_encoder_1.counterZ0Z_2 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_1 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_2 ),
            .clk(N__94081),
            .ce(),
            .sr(N__53202));
    defparam \ppm_encoder_1.counter_3_LC_12_2_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_3_LC_12_2_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_3_LC_12_2_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_3_LC_12_2_3  (
            .in0(_gnd_net_),
            .in1(N__53154),
            .in2(_gnd_net_),
            .in3(N__53134),
            .lcout(\ppm_encoder_1.counterZ0Z_3 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_2 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_3 ),
            .clk(N__94081),
            .ce(),
            .sr(N__53202));
    defparam \ppm_encoder_1.counter_4_LC_12_2_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_4_LC_12_2_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_4_LC_12_2_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_4_LC_12_2_4  (
            .in0(_gnd_net_),
            .in1(N__53131),
            .in2(_gnd_net_),
            .in3(N__53113),
            .lcout(\ppm_encoder_1.counterZ0Z_4 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_3 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_4 ),
            .clk(N__94081),
            .ce(),
            .sr(N__53202));
    defparam \ppm_encoder_1.counter_5_LC_12_2_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_5_LC_12_2_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_5_LC_12_2_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_5_LC_12_2_5  (
            .in0(_gnd_net_),
            .in1(N__53110),
            .in2(_gnd_net_),
            .in3(N__53092),
            .lcout(\ppm_encoder_1.counterZ0Z_5 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_4 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_5 ),
            .clk(N__94081),
            .ce(),
            .sr(N__53202));
    defparam \ppm_encoder_1.counter_6_LC_12_2_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_6_LC_12_2_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_6_LC_12_2_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_6_LC_12_2_6  (
            .in0(_gnd_net_),
            .in1(N__53089),
            .in2(_gnd_net_),
            .in3(N__53071),
            .lcout(\ppm_encoder_1.counterZ0Z_6 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_5 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_6 ),
            .clk(N__94081),
            .ce(),
            .sr(N__53202));
    defparam \ppm_encoder_1.counter_7_LC_12_2_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_7_LC_12_2_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_7_LC_12_2_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_7_LC_12_2_7  (
            .in0(_gnd_net_),
            .in1(N__53066),
            .in2(_gnd_net_),
            .in3(N__53044),
            .lcout(\ppm_encoder_1.counterZ0Z_7 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_6 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_7 ),
            .clk(N__94081),
            .ce(),
            .sr(N__53202));
    defparam \ppm_encoder_1.counter_8_LC_12_3_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_8_LC_12_3_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_8_LC_12_3_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_8_LC_12_3_0  (
            .in0(_gnd_net_),
            .in1(N__53040),
            .in2(_gnd_net_),
            .in3(N__53020),
            .lcout(\ppm_encoder_1.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_12_3_0_),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_8 ),
            .clk(N__94084),
            .ce(),
            .sr(N__53201));
    defparam \ppm_encoder_1.counter_9_LC_12_3_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_9_LC_12_3_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_9_LC_12_3_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_9_LC_12_3_1  (
            .in0(_gnd_net_),
            .in1(N__53016),
            .in2(_gnd_net_),
            .in3(N__52996),
            .lcout(\ppm_encoder_1.counterZ0Z_9 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_8 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_9 ),
            .clk(N__94084),
            .ce(),
            .sr(N__53201));
    defparam \ppm_encoder_1.counter_10_LC_12_3_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_10_LC_12_3_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_10_LC_12_3_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_10_LC_12_3_2  (
            .in0(_gnd_net_),
            .in1(N__52992),
            .in2(_gnd_net_),
            .in3(N__52972),
            .lcout(\ppm_encoder_1.counterZ0Z_10 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_9 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_10 ),
            .clk(N__94084),
            .ce(),
            .sr(N__53201));
    defparam \ppm_encoder_1.counter_11_LC_12_3_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_11_LC_12_3_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_11_LC_12_3_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_11_LC_12_3_3  (
            .in0(_gnd_net_),
            .in1(N__53421),
            .in2(_gnd_net_),
            .in3(N__53401),
            .lcout(\ppm_encoder_1.counterZ0Z_11 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_10 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_11 ),
            .clk(N__94084),
            .ce(),
            .sr(N__53201));
    defparam \ppm_encoder_1.counter_12_LC_12_3_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_12_LC_12_3_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_12_LC_12_3_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_12_LC_12_3_4  (
            .in0(_gnd_net_),
            .in1(N__53390),
            .in2(_gnd_net_),
            .in3(N__53368),
            .lcout(\ppm_encoder_1.counterZ0Z_12 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_11 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_12 ),
            .clk(N__94084),
            .ce(),
            .sr(N__53201));
    defparam \ppm_encoder_1.counter_13_LC_12_3_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_13_LC_12_3_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_13_LC_12_3_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_13_LC_12_3_5  (
            .in0(_gnd_net_),
            .in1(N__53360),
            .in2(_gnd_net_),
            .in3(N__53338),
            .lcout(\ppm_encoder_1.counterZ0Z_13 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_12 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_13 ),
            .clk(N__94084),
            .ce(),
            .sr(N__53201));
    defparam \ppm_encoder_1.counter_14_LC_12_3_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_14_LC_12_3_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_14_LC_12_3_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_14_LC_12_3_6  (
            .in0(_gnd_net_),
            .in1(N__53333),
            .in2(_gnd_net_),
            .in3(N__53317),
            .lcout(\ppm_encoder_1.counterZ0Z_14 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_13 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_14 ),
            .clk(N__94084),
            .ce(),
            .sr(N__53201));
    defparam \ppm_encoder_1.counter_15_LC_12_3_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_15_LC_12_3_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_15_LC_12_3_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_15_LC_12_3_7  (
            .in0(_gnd_net_),
            .in1(N__53312),
            .in2(_gnd_net_),
            .in3(N__53296),
            .lcout(\ppm_encoder_1.counterZ0Z_15 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_14 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_15 ),
            .clk(N__94084),
            .ce(),
            .sr(N__53201));
    defparam \ppm_encoder_1.counter_16_LC_12_4_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_16_LC_12_4_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_16_LC_12_4_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_16_LC_12_4_0  (
            .in0(_gnd_net_),
            .in1(N__53285),
            .in2(_gnd_net_),
            .in3(N__53266),
            .lcout(\ppm_encoder_1.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_12_4_0_),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_16 ),
            .clk(N__94087),
            .ce(),
            .sr(N__53203));
    defparam \ppm_encoder_1.counter_17_LC_12_4_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_17_LC_12_4_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_17_LC_12_4_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_17_LC_12_4_1  (
            .in0(_gnd_net_),
            .in1(N__53255),
            .in2(_gnd_net_),
            .in3(N__53233),
            .lcout(\ppm_encoder_1.counterZ0Z_17 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_16 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_17 ),
            .clk(N__94087),
            .ce(),
            .sr(N__53203));
    defparam \ppm_encoder_1.counter_18_LC_12_4_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_18_LC_12_4_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_18_LC_12_4_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.counter_18_LC_12_4_2  (
            .in0(_gnd_net_),
            .in1(N__53226),
            .in2(_gnd_net_),
            .in3(N__53230),
            .lcout(\ppm_encoder_1.counterZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94087),
            .ce(),
            .sr(N__53203));
    defparam \pid_side.source_pid_1_esr_12_LC_12_5_0 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_esr_12_LC_12_5_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_esr_12_LC_12_5_0 .LUT_INIT=16'b1111000100000000;
    LogicCell40 \pid_side.source_pid_1_esr_12_LC_12_5_0  (
            .in0(N__64803),
            .in1(N__62039),
            .in2(N__65134),
            .in3(N__64839),
            .lcout(side_order_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94092),
            .ce(N__59148),
            .sr(N__59399));
    defparam \pid_side.source_pid_1_esr_13_LC_12_5_1 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_esr_13_LC_12_5_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_esr_13_LC_12_5_1 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \pid_side.source_pid_1_esr_13_LC_12_5_1  (
            .in0(N__62040),
            .in1(N__65130),
            .in2(_gnd_net_),
            .in3(N__64802),
            .lcout(side_order_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94092),
            .ce(N__59148),
            .sr(N__59399));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_14_LC_12_5_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_14_LC_12_5_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_14_LC_12_5_2 .LUT_INIT=16'b0000010100100010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_14_LC_12_5_2  (
            .in0(N__54107),
            .in1(N__53911),
            .in2(N__53890),
            .in3(N__54231),
            .lcout(),
            .ltout(\ppm_encoder_1.pulses2count_9_i_0_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_14_LC_12_5_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_14_LC_12_5_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_14_LC_12_5_3 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_14_LC_12_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__53851),
            .in3(N__53501),
            .lcout(\ppm_encoder_1.pulses2count_9_i_1_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_5_LC_12_5_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_5_LC_12_5_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_5_LC_12_5_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_5_LC_12_5_4  (
            .in0(N__53503),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53833),
            .lcout(\ppm_encoder_1.pulses2count_9_i_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIGJLB1_1_LC_12_5_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIGJLB1_1_LC_12_5_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIGJLB1_1_LC_12_5_5 .LUT_INIT=16'b1111111010101010;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_RNIGJLB1_1_LC_12_5_5  (
            .in0(N__53798),
            .in1(N__54106),
            .in2(N__54251),
            .in3(N__53698),
            .lcout(\ppm_encoder_1.N_301 ),
            .ltout(\ppm_encoder_1.N_301_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_6_LC_12_5_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_6_LC_12_5_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_6_LC_12_5_6 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_6_LC_12_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__53557),
            .in3(N__53554),
            .lcout(\ppm_encoder_1.pulses2count_9_0_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_7_LC_12_5_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_7_LC_12_5_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_7_LC_12_5_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_7_LC_12_5_7  (
            .in0(N__53995),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53502),
            .lcout(\ppm_encoder_1.pulses2count_9_i_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.source_pid_1_10_LC_12_6_0 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_10_LC_12_6_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_10_LC_12_6_0 .LUT_INIT=16'b1110111011100010;
    LogicCell40 \pid_side.source_pid_1_10_LC_12_6_0  (
            .in0(N__53441),
            .in1(N__60746),
            .in2(N__64432),
            .in3(N__59249),
            .lcout(side_order_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94098),
            .ce(),
            .sr(N__59410));
    defparam \pid_side.source_pid_1_11_LC_12_6_1 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_11_LC_12_6_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_11_LC_12_6_1 .LUT_INIT=16'b1110111111100000;
    LogicCell40 \pid_side.source_pid_1_11_LC_12_6_1  (
            .in0(N__59242),
            .in1(N__64882),
            .in2(N__60754),
            .in3(N__54473),
            .lcout(side_order_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94098),
            .ce(),
            .sr(N__59410));
    defparam \pid_side.source_pid_1_6_LC_12_6_2 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_6_LC_12_6_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_6_LC_12_6_2 .LUT_INIT=16'b1110111011100010;
    LogicCell40 \pid_side.source_pid_1_6_LC_12_6_2  (
            .in0(N__54437),
            .in1(N__60747),
            .in2(N__64564),
            .in3(N__59250),
            .lcout(side_order_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94098),
            .ce(),
            .sr(N__59410));
    defparam \pid_side.source_pid_1_7_LC_12_6_3 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_7_LC_12_6_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_7_LC_12_6_3 .LUT_INIT=16'b1110111011100100;
    LogicCell40 \pid_side.source_pid_1_7_LC_12_6_3  (
            .in0(N__60744),
            .in1(N__54410),
            .in2(N__59256),
            .in3(N__64523),
            .lcout(side_order_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94098),
            .ce(),
            .sr(N__59410));
    defparam \pid_side.source_pid_1_8_LC_12_6_4 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_8_LC_12_6_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_8_LC_12_6_4 .LUT_INIT=16'b1110111011100010;
    LogicCell40 \pid_side.source_pid_1_8_LC_12_6_4  (
            .in0(N__54374),
            .in1(N__60748),
            .in2(N__64486),
            .in3(N__59251),
            .lcout(side_order_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94098),
            .ce(),
            .sr(N__59410));
    defparam \pid_side.source_pid_1_9_LC_12_6_5 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_9_LC_12_6_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_9_LC_12_6_5 .LUT_INIT=16'b1110111011100100;
    LogicCell40 \pid_side.source_pid_1_9_LC_12_6_5  (
            .in0(N__60745),
            .in1(N__54341),
            .in2(N__59257),
            .in3(N__64456),
            .lcout(side_order_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94098),
            .ce(),
            .sr(N__59410));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIPJL01_3_LC_12_7_4 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIPJL01_3_LC_12_7_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIPJL01_3_LC_12_7_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIPJL01_3_LC_12_7_4  (
            .in0(N__62768),
            .in1(N__59602),
            .in2(_gnd_net_),
            .in3(N__59666),
            .lcout(\pid_side.error_i_acumm_13_0_a2_3_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_7_LC_12_8_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_7_LC_12_8_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_7_LC_12_8_3 .LUT_INIT=16'b0000001101010000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_7_LC_12_8_3  (
            .in0(N__54315),
            .in1(N__54288),
            .in2(N__54261),
            .in3(N__54102),
            .lcout(\ppm_encoder_1.pulses2count_9_i_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNIOU0N_4_LC_12_9_0 .C_ON=1'b0;
    defparam \uart_drone.state_RNIOU0N_4_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNIOU0N_4_LC_12_9_0 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \uart_drone.state_RNIOU0N_4_LC_12_9_0  (
            .in0(N__53979),
            .in1(N__54814),
            .in2(_gnd_net_),
            .in3(N__70805),
            .lcout(\uart_drone.state_RNIOU0NZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNO_0_0_LC_12_9_2 .C_ON=1'b0;
    defparam \uart_drone.state_RNO_0_0_LC_12_9_2 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNO_0_0_LC_12_9_2 .LUT_INIT=16'b0000000011011101;
    LogicCell40 \uart_drone.state_RNO_0_0_LC_12_9_2  (
            .in0(N__54699),
            .in1(N__56862),
            .in2(_gnd_net_),
            .in3(N__70806),
            .lcout(),
            .ltout(\uart_drone.state_srsts_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_0_LC_12_9_3 .C_ON=1'b0;
    defparam \uart_drone.state_0_LC_12_9_3 .SEQ_MODE=4'b1000;
    defparam \uart_drone.state_0_LC_12_9_3 .LUT_INIT=16'b1010111110001111;
    LogicCell40 \uart_drone.state_0_LC_12_9_3  (
            .in0(N__54815),
            .in1(N__54784),
            .in2(N__54730),
            .in3(N__54727),
            .lcout(\uart_drone.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94118),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNI2U6A8_3_LC_12_9_5 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNI2U6A8_3_LC_12_9_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNI2U6A8_3_LC_12_9_5 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNI2U6A8_3_LC_12_9_5  (
            .in0(N__56401),
            .in1(N__60430),
            .in2(N__54688),
            .in3(N__59715),
            .lcout(\pid_side.N_634 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.source_pid_1_10_LC_12_10_0 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_10_LC_12_10_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_10_LC_12_10_0 .LUT_INIT=16'b1111110010111000;
    LogicCell40 \pid_front.source_pid_1_10_LC_12_10_0  (
            .in0(N__60181),
            .in1(N__70520),
            .in2(N__54671),
            .in3(N__58207),
            .lcout(front_order_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94128),
            .ce(),
            .sr(N__59991));
    defparam \pid_front.source_pid_1_11_LC_12_10_1 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_11_LC_12_10_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_11_LC_12_10_1 .LUT_INIT=16'b1111101011011000;
    LogicCell40 \pid_front.source_pid_1_11_LC_12_10_1  (
            .in0(N__70517),
            .in1(N__60182),
            .in2(N__54641),
            .in3(N__58654),
            .lcout(front_order_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94128),
            .ce(),
            .sr(N__59991));
    defparam \pid_front.source_pid_1_6_LC_12_10_2 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_6_LC_12_10_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_6_LC_12_10_2 .LUT_INIT=16'b1111110010111000;
    LogicCell40 \pid_front.source_pid_1_6_LC_12_10_2  (
            .in0(N__60183),
            .in1(N__70521),
            .in2(N__54602),
            .in3(N__58405),
            .lcout(front_order_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94128),
            .ce(),
            .sr(N__59991));
    defparam \pid_front.source_pid_1_7_LC_12_10_3 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_7_LC_12_10_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_7_LC_12_10_3 .LUT_INIT=16'b1111101011011000;
    LogicCell40 \pid_front.source_pid_1_7_LC_12_10_3  (
            .in0(N__70518),
            .in1(N__60184),
            .in2(N__54569),
            .in3(N__58369),
            .lcout(front_order_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94128),
            .ce(),
            .sr(N__59991));
    defparam \pid_front.source_pid_1_8_LC_12_10_4 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_8_LC_12_10_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_8_LC_12_10_4 .LUT_INIT=16'b1111101111001000;
    LogicCell40 \pid_front.source_pid_1_8_LC_12_10_4  (
            .in0(N__60185),
            .in1(N__70522),
            .in2(N__58297),
            .in3(N__54536),
            .lcout(front_order_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94128),
            .ce(),
            .sr(N__59991));
    defparam \pid_front.source_pid_1_9_LC_12_10_5 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_9_LC_12_10_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_9_LC_12_10_5 .LUT_INIT=16'b1111101011011000;
    LogicCell40 \pid_front.source_pid_1_9_LC_12_10_5  (
            .in0(N__70519),
            .in1(N__60186),
            .in2(N__54509),
            .in3(N__58240),
            .lcout(front_order_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94128),
            .ce(),
            .sr(N__59991));
    defparam \pid_side.error_d_reg_esr_RNI2OIO_13_LC_12_10_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_RNI2OIO_13_LC_12_10_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_esr_RNI2OIO_13_LC_12_10_6 .LUT_INIT=16'b1101110101000100;
    LogicCell40 \pid_side.error_d_reg_esr_RNI2OIO_13_LC_12_10_6  (
            .in0(N__79122),
            .in1(N__90918),
            .in2(_gnd_net_),
            .in3(N__91494),
            .lcout(\pid_side.error_d_reg_esr_RNI2OIOZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_esr_RNI2OIO_1_13_LC_12_10_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_RNI2OIO_1_13_LC_12_10_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_esr_RNI2OIO_1_13_LC_12_10_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_side.error_d_reg_esr_RNI2OIO_1_13_LC_12_10_7  (
            .in0(N__91495),
            .in1(_gnd_net_),
            .in2(N__90922),
            .in3(N__79123),
            .lcout(\pid_side.N_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.source_pid_1_esr_1_LC_12_11_0 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_esr_1_LC_12_11_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_esr_1_LC_12_11_0 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \pid_front.source_pid_1_esr_1_LC_12_11_0  (
            .in0(N__60179),
            .in1(N__60122),
            .in2(_gnd_net_),
            .in3(N__58165),
            .lcout(front_order_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94136),
            .ce(N__60036),
            .sr(N__59990));
    defparam \pid_front.source_pid_1_esr_4_LC_12_11_5 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_esr_4_LC_12_11_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_esr_4_LC_12_11_5 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \pid_front.source_pid_1_esr_4_LC_12_11_5  (
            .in0(N__60123),
            .in1(N__60180),
            .in2(_gnd_net_),
            .in3(N__58471),
            .lcout(front_order_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94136),
            .ce(N__60036),
            .sr(N__59990));
    defparam \reset_module_System.count_2_LC_12_12_0 .C_ON=1'b0;
    defparam \reset_module_System.count_2_LC_12_12_0 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_2_LC_12_12_0 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \reset_module_System.count_2_LC_12_12_0  (
            .in0(N__54917),
            .in1(N__55027),
            .in2(N__54946),
            .in3(N__54952),
            .lcout(\reset_module_System.countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94143),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.state_RNIM6IF_1_LC_12_12_2 .C_ON=1'b0;
    defparam \pid_side.state_RNIM6IF_1_LC_12_12_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.state_RNIM6IF_1_LC_12_12_2 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \pid_side.state_RNIM6IF_1_LC_12_12_2  (
            .in0(_gnd_net_),
            .in1(N__60715),
            .in2(_gnd_net_),
            .in3(N__70704),
            .lcout(\pid_side.N_205 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.state_RNIVIRQ_0_LC_12_12_3 .C_ON=1'b0;
    defparam \pid_front.state_RNIVIRQ_0_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.state_RNIVIRQ_0_LC_12_12_3 .LUT_INIT=16'b1010101110101010;
    LogicCell40 \pid_front.state_RNIVIRQ_0_LC_12_12_3  (
            .in0(N__70705),
            .in1(N__70604),
            .in2(N__70516),
            .in3(N__69183),
            .lcout(\pid_front.state_RNIVIRQZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.reset_LC_12_12_5 .C_ON=1'b0;
    defparam \reset_module_System.reset_LC_12_12_5 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.reset_LC_12_12_5 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \reset_module_System.reset_LC_12_12_5  (
            .in0(N__55026),
            .in1(N__54941),
            .in2(_gnd_net_),
            .in3(N__54918),
            .lcout(reset_system),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94143),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNI9O1P_2_LC_12_13_0 .C_ON=1'b0;
    defparam \reset_module_System.count_RNI9O1P_2_LC_12_13_0 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNI9O1P_2_LC_12_13_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \reset_module_System.count_RNI9O1P_2_LC_12_13_0  (
            .in0(N__54898),
            .in1(N__54882),
            .in2(N__54868),
            .in3(N__54850),
            .lcout(\reset_module_System.reset6_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.state_RNISV141_0_LC_12_13_1 .C_ON=1'b0;
    defparam \pid_front.state_RNISV141_0_LC_12_13_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.state_RNISV141_0_LC_12_13_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pid_front.state_RNISV141_0_LC_12_13_1  (
            .in0(_gnd_net_),
            .in1(N__54829),
            .in2(_gnd_net_),
            .in3(N__93124),
            .lcout(\pid_front.N_787_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.un1_state57_i_LC_12_13_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.un1_state57_i_LC_12_13_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.un1_state57_i_LC_12_13_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \Commands_frame_decoder.un1_state57_i_LC_12_13_2  (
            .in0(N__70731),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55278),
            .lcout(\Commands_frame_decoder.un1_state57_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.N_27_0_i_i_a2_2_LC_12_13_3 .C_ON=1'b0;
    defparam \pid_side.N_27_0_i_i_a2_2_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.N_27_0_i_i_a2_2_LC_12_13_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \pid_side.N_27_0_i_i_a2_2_LC_12_13_3  (
            .in0(_gnd_net_),
            .in1(N__83183),
            .in2(_gnd_net_),
            .in3(N__82257),
            .lcout(pid_side_N_493),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.state_RNIQLTD_1_LC_12_13_5 .C_ON=1'b0;
    defparam \pid_front.state_RNIQLTD_1_LC_12_13_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.state_RNIQLTD_1_LC_12_13_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \pid_front.state_RNIQLTD_1_LC_12_13_5  (
            .in0(_gnd_net_),
            .in1(N__70498),
            .in2(_gnd_net_),
            .in3(N__70729),
            .lcout(\pid_front.N_205 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.state_RNINK4U_0_LC_12_13_6 .C_ON=1'b0;
    defparam \pid_side.state_RNINK4U_0_LC_12_13_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.state_RNINK4U_0_LC_12_13_6 .LUT_INIT=16'b1010101010111010;
    LogicCell40 \pid_side.state_RNINK4U_0_LC_12_13_6  (
            .in0(N__70730),
            .in1(N__60711),
            .in2(N__69191),
            .in3(N__60798),
            .lcout(),
            .ltout(\pid_side.state_RNINK4UZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.state_RNIK1B71_0_LC_12_13_7 .C_ON=1'b0;
    defparam \pid_side.state_RNIK1B71_0_LC_12_13_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.state_RNIK1B71_0_LC_12_13_7 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \pid_side.state_RNIK1B71_0_LC_12_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__55084),
            .in3(N__93125),
            .lcout(\pid_side.N_868_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_2_c_RNIFP8G1_LC_12_14_5 .C_ON=1'b0;
    defparam \pid_front.error_cry_2_c_RNIFP8G1_LC_12_14_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_2_c_RNIFP8G1_LC_12_14_5 .LUT_INIT=16'b0010010101110101;
    LogicCell40 \pid_front.error_cry_2_c_RNIFP8G1_LC_12_14_5  (
            .in0(N__82686),
            .in1(N__74076),
            .in2(N__79654),
            .in3(N__79856),
            .lcout(\pid_front.error_cry_2_c_RNIFP8GZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNI34OR1_21_LC_12_14_6 .C_ON=1'b0;
    defparam \reset_module_System.count_RNI34OR1_21_LC_12_14_6 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNI34OR1_21_LC_12_14_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \reset_module_System.count_RNI34OR1_21_LC_12_14_6  (
            .in0(N__55080),
            .in1(N__55069),
            .in2(N__55057),
            .in3(N__55042),
            .lcout(\reset_module_System.reset6_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_9_LC_12_15_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_9_LC_12_15_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_9_LC_12_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_9_LC_12_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57319),
            .lcout(\dron_frame_decoder_1.drone_H_disp_front_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94181),
            .ce(N__57655),
            .sr(N__86434));
    defparam \pid_front.error_cry_0_c_RNIVSLV_LC_12_16_0 .C_ON=1'b0;
    defparam \pid_front.error_cry_0_c_RNIVSLV_LC_12_16_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_c_RNIVSLV_LC_12_16_0 .LUT_INIT=16'b0000101011001110;
    LogicCell40 \pid_front.error_cry_0_c_RNIVSLV_LC_12_16_0  (
            .in0(N__83167),
            .in1(N__82255),
            .in2(N__84660),
            .in3(N__74133),
            .lcout(\pid_front.m64_i_o2_0 ),
            .ltout(\pid_front.m64_i_o2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_4_14_LC_12_16_1 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_4_14_LC_12_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_4_14_LC_12_16_1 .LUT_INIT=16'b1111100011111001;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_4_14_LC_12_16_1  (
            .in0(N__90646),
            .in1(N__82688),
            .in2(N__55306),
            .in3(N__79972),
            .lcout(),
            .ltout(\pid_front.error_i_reg_esr_RNO_4_0_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_2_14_LC_12_16_2 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_2_14_LC_12_16_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_2_14_LC_12_16_2 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_2_14_LC_12_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__55303),
            .in3(N__84836),
            .lcout(\pid_front.N_111 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_1_c_RNILQ1F2_LC_12_16_3 .C_ON=1'b0;
    defparam \pid_front.error_cry_1_c_RNILQ1F2_LC_12_16_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_1_c_RNILQ1F2_LC_12_16_3 .LUT_INIT=16'b0011000000010000;
    LogicCell40 \pid_front.error_cry_1_c_RNILQ1F2_LC_12_16_3  (
            .in0(N__81309),
            .in1(N__55300),
            .in2(N__87803),
            .in3(N__79973),
            .lcout(\pid_front.error_cry_1_c_RNILQ1FZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_c_RNIVSLV_0_LC_12_16_4 .C_ON=1'b0;
    defparam \pid_front.error_cry_0_c_RNIVSLV_0_LC_12_16_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_c_RNIVSLV_0_LC_12_16_4 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \pid_front.error_cry_0_c_RNIVSLV_0_LC_12_16_4  (
            .in0(N__83166),
            .in1(N__82254),
            .in2(N__84659),
            .in3(N__74132),
            .lcout(\pid_front.m1_0_03 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_1_c_RNIR72C1_LC_12_16_5 .C_ON=1'b0;
    defparam \pid_front.error_cry_1_c_RNIR72C1_LC_12_16_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_1_c_RNIR72C1_LC_12_16_5 .LUT_INIT=16'b0111011101011111;
    LogicCell40 \pid_front.error_cry_1_c_RNIR72C1_LC_12_16_5  (
            .in0(N__82256),
            .in1(N__79971),
            .in2(N__79890),
            .in3(N__83168),
            .lcout(),
            .ltout(\pid_front.m9_2_03_3_i_0_o2_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_1_c_RNI624A3_LC_12_16_6 .C_ON=1'b0;
    defparam \pid_front.error_cry_1_c_RNI624A3_LC_12_16_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_1_c_RNI624A3_LC_12_16_6 .LUT_INIT=16'b1010111000001100;
    LogicCell40 \pid_front.error_cry_1_c_RNI624A3_LC_12_16_6  (
            .in0(N__74958),
            .in1(N__83475),
            .in2(N__55294),
            .in3(N__69552),
            .lcout(),
            .ltout(\pid_front.m9_2_03_3_i_0_o2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_2_c_RNI46SR4_LC_12_16_7 .C_ON=1'b0;
    defparam \pid_front.error_cry_2_c_RNI46SR4_LC_12_16_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_2_c_RNI46SR4_LC_12_16_7 .LUT_INIT=16'b1111110011110000;
    LogicCell40 \pid_front.error_cry_2_c_RNI46SR4_LC_12_16_7  (
            .in0(_gnd_net_),
            .in1(N__60652),
            .in2(N__55291),
            .in3(N__74062),
            .lcout(\pid_front.m9_2_03_3_i_0_o2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_axb_3_LC_12_17_0 .C_ON=1'b0;
    defparam \pid_front.error_axb_3_LC_12_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_axb_3_LC_12_17_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_front.error_axb_3_LC_12_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55288),
            .lcout(\pid_front.error_axbZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_3_LC_12_17_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_3_LC_12_17_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_3_LC_12_17_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_3_LC_12_17_1  (
            .in0(N__58012),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(drone_H_disp_front_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94210),
            .ce(N__57414),
            .sr(N__86415));
    defparam \pid_side.error_axb_1_LC_12_17_2 .C_ON=1'b0;
    defparam \pid_side.error_axb_1_LC_12_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_axb_1_LC_12_17_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_side.error_axb_1_LC_12_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57256),
            .lcout(\pid_side.error_axbZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_axb_2_LC_12_17_3 .C_ON=1'b0;
    defparam \pid_side.error_axb_2_LC_12_17_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_axb_2_LC_12_17_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_side.error_axb_2_LC_12_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57184),
            .lcout(\pid_side.error_axbZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_axb_3_LC_12_17_4 .C_ON=1'b0;
    defparam \pid_side.error_axb_3_LC_12_17_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_axb_3_LC_12_17_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_side.error_axb_3_LC_12_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57178),
            .lcout(\pid_side.error_axbZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_2_LC_12_17_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_2_LC_12_17_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_2_LC_12_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_2_LC_12_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57243),
            .lcout(drone_H_disp_front_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94210),
            .ce(N__57414),
            .sr(N__86415));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_4_LC_12_17_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_4_LC_12_17_7 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_4_LC_12_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_4_LC_12_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57948),
            .lcout(\dron_frame_decoder_1.drone_H_disp_front_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94210),
            .ce(N__57414),
            .sr(N__86415));
    defparam \pid_front.error_cry_0_c_inv_LC_12_18_0 .C_ON=1'b1;
    defparam \pid_front.error_cry_0_c_inv_LC_12_18_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_c_inv_LC_12_18_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_front.error_cry_0_c_inv_LC_12_18_0  (
            .in0(_gnd_net_),
            .in1(N__55348),
            .in2(_gnd_net_),
            .in3(N__57424),
            .lcout(\pid_front.error_axb_0 ),
            .ltout(),
            .carryin(bfn_12_18_0_),
            .carryout(\pid_front.error_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_c_RNIC7KB_LC_12_18_1 .C_ON=1'b1;
    defparam \pid_front.error_cry_0_c_RNIC7KB_LC_12_18_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_c_RNIC7KB_LC_12_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_cry_0_c_RNIC7KB_LC_12_18_1  (
            .in0(_gnd_net_),
            .in1(N__55342),
            .in2(_gnd_net_),
            .in3(N__55336),
            .lcout(\pid_front.error_1 ),
            .ltout(),
            .carryin(\pid_front.error_cry_0 ),
            .carryout(\pid_front.error_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_1_c_RNIEALB_LC_12_18_2 .C_ON=1'b1;
    defparam \pid_front.error_cry_1_c_RNIEALB_LC_12_18_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_1_c_RNIEALB_LC_12_18_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_cry_1_c_RNIEALB_LC_12_18_2  (
            .in0(_gnd_net_),
            .in1(N__55333),
            .in2(_gnd_net_),
            .in3(N__55327),
            .lcout(\pid_front.error_2 ),
            .ltout(),
            .carryin(\pid_front.error_cry_1 ),
            .carryout(\pid_front.error_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_2_c_RNIGDMB_LC_12_18_3 .C_ON=1'b1;
    defparam \pid_front.error_cry_2_c_RNIGDMB_LC_12_18_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_2_c_RNIGDMB_LC_12_18_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_cry_2_c_RNIGDMB_LC_12_18_3  (
            .in0(_gnd_net_),
            .in1(N__55324),
            .in2(_gnd_net_),
            .in3(N__55318),
            .lcout(\pid_front.error_3 ),
            .ltout(),
            .carryin(\pid_front.error_cry_2 ),
            .carryout(\pid_front.error_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_3_c_RNIABAG_LC_12_18_4 .C_ON=1'b1;
    defparam \pid_front.error_cry_3_c_RNIABAG_LC_12_18_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_3_c_RNIABAG_LC_12_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_3_c_RNIABAG_LC_12_18_4  (
            .in0(_gnd_net_),
            .in1(N__55315),
            .in2(N__55483),
            .in3(N__55309),
            .lcout(\pid_front.error_4 ),
            .ltout(),
            .carryin(\pid_front.error_cry_3 ),
            .carryout(\pid_front.error_cry_0_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_0_c_RNIOQKB_LC_12_18_5 .C_ON=1'b1;
    defparam \pid_front.error_cry_0_0_c_RNIOQKB_LC_12_18_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_0_c_RNIOQKB_LC_12_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_0_0_c_RNIOQKB_LC_12_18_5  (
            .in0(_gnd_net_),
            .in1(N__55408),
            .in2(N__55471),
            .in3(N__55402),
            .lcout(\pid_front.error_5 ),
            .ltout(),
            .carryin(\pid_front.error_cry_0_0 ),
            .carryout(\pid_front.error_cry_1_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_1_0_c_RNIR0RF_LC_12_18_6 .C_ON=1'b1;
    defparam \pid_front.error_cry_1_0_c_RNIR0RF_LC_12_18_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_1_0_c_RNIR0RF_LC_12_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_1_0_c_RNIR0RF_LC_12_18_6  (
            .in0(_gnd_net_),
            .in1(N__55399),
            .in2(N__55459),
            .in3(N__55393),
            .lcout(\pid_front.error_6 ),
            .ltout(),
            .carryin(\pid_front.error_cry_1_0 ),
            .carryout(\pid_front.error_cry_2_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_2_0_c_RNIU61K_LC_12_18_7 .C_ON=1'b1;
    defparam \pid_front.error_cry_2_0_c_RNIU61K_LC_12_18_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_2_0_c_RNIU61K_LC_12_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_2_0_c_RNIU61K_LC_12_18_7  (
            .in0(_gnd_net_),
            .in1(N__57043),
            .in2(N__55447),
            .in3(N__55390),
            .lcout(\pid_front.error_7 ),
            .ltout(),
            .carryin(\pid_front.error_cry_2_0 ),
            .carryout(\pid_front.error_cry_3_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_3_0_c_RNI1D7O_LC_12_19_0 .C_ON=1'b1;
    defparam \pid_front.error_cry_3_0_c_RNI1D7O_LC_12_19_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_3_0_c_RNI1D7O_LC_12_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_3_0_c_RNI1D7O_LC_12_19_0  (
            .in0(_gnd_net_),
            .in1(N__55435),
            .in2(N__57034),
            .in3(N__55387),
            .lcout(\pid_front.error_8 ),
            .ltout(),
            .carryin(bfn_12_19_0_),
            .carryout(\pid_front.error_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_4_c_RNILNBG_LC_12_19_1 .C_ON=1'b1;
    defparam \pid_front.error_cry_4_c_RNILNBG_LC_12_19_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_4_c_RNILNBG_LC_12_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_4_c_RNILNBG_LC_12_19_1  (
            .in0(_gnd_net_),
            .in1(N__57016),
            .in2(N__55429),
            .in3(N__55384),
            .lcout(\pid_front.error_9 ),
            .ltout(),
            .carryin(\pid_front.error_cry_4 ),
            .carryout(\pid_front.error_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_5_c_RNIVNFF_LC_12_19_2 .C_ON=1'b1;
    defparam \pid_front.error_cry_5_c_RNIVNFF_LC_12_19_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_5_c_RNIVNFF_LC_12_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_5_c_RNIVNFF_LC_12_19_2  (
            .in0(_gnd_net_),
            .in1(N__55381),
            .in2(N__55420),
            .in3(N__55375),
            .lcout(\pid_front.error_10 ),
            .ltout(),
            .carryin(\pid_front.error_cry_5 ),
            .carryout(\pid_front.error_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_6_c_RNI3VJG_LC_12_19_3 .C_ON=1'b1;
    defparam \pid_front.error_cry_6_c_RNI3VJG_LC_12_19_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_6_c_RNI3VJG_LC_12_19_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_front.error_cry_6_c_RNI3VJG_LC_12_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__58102),
            .in3(N__55372),
            .lcout(\pid_front.error_11 ),
            .ltout(),
            .carryin(\pid_front.error_cry_6 ),
            .carryout(\pid_front.error_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_7_c_RNIAPPM_LC_12_19_4 .C_ON=1'b1;
    defparam \pid_front.error_cry_7_c_RNIAPPM_LC_12_19_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_7_c_RNIAPPM_LC_12_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_7_c_RNIAPPM_LC_12_19_4  (
            .in0(_gnd_net_),
            .in1(N__57436),
            .in2(N__58090),
            .in3(N__55369),
            .lcout(\pid_front.error_12 ),
            .ltout(),
            .carryin(\pid_front.error_cry_7 ),
            .carryout(\pid_front.error_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_8_c_RNIAC2E_LC_12_19_5 .C_ON=1'b1;
    defparam \pid_front.error_cry_8_c_RNIAC2E_LC_12_19_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_8_c_RNIAC2E_LC_12_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_8_c_RNIAC2E_LC_12_19_5  (
            .in0(_gnd_net_),
            .in1(N__58072),
            .in2(N__57813),
            .in3(N__55366),
            .lcout(\pid_front.error_13 ),
            .ltout(),
            .carryin(\pid_front.error_cry_8 ),
            .carryout(\pid_front.error_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_9_c_RNIDG3E_LC_12_19_6 .C_ON=1'b1;
    defparam \pid_front.error_cry_9_c_RNIDG3E_LC_12_19_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_9_c_RNIDG3E_LC_12_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_9_c_RNIDG3E_LC_12_19_6  (
            .in0(_gnd_net_),
            .in1(N__55581),
            .in2(N__55498),
            .in3(N__55489),
            .lcout(\pid_front.error_14 ),
            .ltout(),
            .carryin(\pid_front.error_cry_9 ),
            .carryout(\pid_front.error_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_10_c_RNINTDI_LC_12_19_7 .C_ON=1'b0;
    defparam \pid_front.error_cry_10_c_RNINTDI_LC_12_19_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_10_c_RNINTDI_LC_12_19_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_cry_10_c_RNINTDI_LC_12_19_7  (
            .in0(N__55582),
            .in1(N__57733),
            .in2(_gnd_net_),
            .in3(N__55486),
            .lcout(\pid_front.error_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH3data_esr_0_LC_12_20_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_0_LC_12_20_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_0_LC_12_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_0_LC_12_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88261),
            .lcout(front_command_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94261),
            .ce(N__55600),
            .sr(N__86384));
    defparam \Commands_frame_decoder.source_CH3data_esr_1_LC_12_20_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_1_LC_12_20_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_1_LC_12_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_1_LC_12_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85485),
            .lcout(front_command_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94261),
            .ce(N__55600),
            .sr(N__86384));
    defparam \Commands_frame_decoder.source_CH3data_esr_2_LC_12_20_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_2_LC_12_20_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_2_LC_12_20_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_2_LC_12_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__92509),
            .lcout(front_command_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94261),
            .ce(N__55600),
            .sr(N__86384));
    defparam \Commands_frame_decoder.source_CH3data_esr_3_LC_12_20_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_3_LC_12_20_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_3_LC_12_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_3_LC_12_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__92287),
            .lcout(front_command_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94261),
            .ce(N__55600),
            .sr(N__86384));
    defparam \Commands_frame_decoder.source_CH3data_esr_4_LC_12_20_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_4_LC_12_20_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_4_LC_12_20_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_4_LC_12_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88846),
            .lcout(front_command_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94261),
            .ce(N__55600),
            .sr(N__86384));
    defparam \Commands_frame_decoder.source_CH3data_esr_5_LC_12_20_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_5_LC_12_20_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_5_LC_12_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_5_LC_12_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88665),
            .lcout(front_command_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94261),
            .ce(N__55600),
            .sr(N__86384));
    defparam \Commands_frame_decoder.source_CH3data_esr_6_LC_12_20_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_6_LC_12_20_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_6_LC_12_20_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_6_LC_12_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88482),
            .lcout(front_command_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94261),
            .ce(N__55600),
            .sr(N__86384));
    defparam \Commands_frame_decoder.source_CH3data_ess_7_LC_12_20_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_ess_7_LC_12_20_7 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_CH3data_ess_7_LC_12_20_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_ess_7_LC_12_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__92122),
            .lcout(front_command_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94261),
            .ce(N__55600),
            .sr(N__86384));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_14_LC_12_21_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_14_LC_12_21_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_14_LC_12_21_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_14_LC_12_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57148),
            .lcout(drone_H_disp_front_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94280),
            .ce(N__57648),
            .sr(N__86377));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_10_LC_12_21_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_10_LC_12_21_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_10_LC_12_21_5 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_10_LC_12_21_5  (
            .in0(_gnd_net_),
            .in1(N__57250),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\dron_frame_decoder_1.drone_H_disp_front_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94280),
            .ce(N__57648),
            .sr(N__86377));
    defparam \pid_front.pid_prereg_esr_RNI1CIT4_16_LC_12_22_0 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNI1CIT4_16_LC_12_22_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNI1CIT4_16_LC_12_22_0 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \pid_front.pid_prereg_esr_RNI1CIT4_16_LC_12_22_0  (
            .in0(N__55926),
            .in1(N__55558),
            .in2(N__55851),
            .in3(N__55827),
            .lcout(\pid_front.N_175 ),
            .ltout(\pid_front.N_175_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNID3QC5_15_LC_12_22_1 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNID3QC5_15_LC_12_22_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNID3QC5_15_LC_12_22_1 .LUT_INIT=16'b1111111111111010;
    LogicCell40 \pid_front.pid_prereg_esr_RNID3QC5_15_LC_12_22_1  (
            .in0(N__58540),
            .in1(_gnd_net_),
            .in2(N__55540),
            .in3(N__55798),
            .lcout(\pid_front.N_277 ),
            .ltout(\pid_front.N_277_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNI7FE58_0_LC_12_22_2 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNI7FE58_0_LC_12_22_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNI7FE58_0_LC_12_22_2 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \pid_front.pid_prereg_esr_RNI7FE58_0_LC_12_22_2  (
            .in0(N__55533),
            .in1(N__58063),
            .in2(N__55519),
            .in3(N__58048),
            .lcout(\pid_front.N_342 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNIC02A7_30_LC_12_22_3 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNIC02A7_30_LC_12_22_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNIC02A7_30_LC_12_22_3 .LUT_INIT=16'b0001010100000101;
    LogicCell40 \pid_front.pid_prereg_esr_RNIC02A7_30_LC_12_22_3  (
            .in0(N__70972),
            .in1(N__58867),
            .in2(N__70482),
            .in3(N__55516),
            .lcout(),
            .ltout(\pid_front.un1_reset_i_o3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNIJMSRH_30_LC_12_22_4 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNIJMSRH_30_LC_12_22_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNIJMSRH_30_LC_12_22_4 .LUT_INIT=16'b1111111100001011;
    LogicCell40 \pid_front.pid_prereg_esr_RNIJMSRH_30_LC_12_22_4  (
            .in0(N__70973),
            .in1(N__60108),
            .in2(N__55510),
            .in3(N__55507),
            .lcout(\pid_front.un1_reset_0_i_3 ),
            .ltout(\pid_front.un1_reset_0_i_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.state_RNIGVJ0I_1_LC_12_22_5 .C_ON=1'b0;
    defparam \pid_front.state_RNIGVJ0I_1_LC_12_22_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.state_RNIGVJ0I_1_LC_12_22_5 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \pid_front.state_RNIGVJ0I_1_LC_12_22_5  (
            .in0(N__70461),
            .in1(_gnd_net_),
            .in2(N__55501),
            .in3(_gnd_net_),
            .lcout(\pid_front.state_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.source_pid_1_esr_13_LC_12_22_6 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_esr_13_LC_12_22_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_esr_13_LC_12_22_6 .LUT_INIT=16'b1111111100001010;
    LogicCell40 \pid_front.source_pid_1_esr_13_LC_12_22_6  (
            .in0(N__55714),
            .in1(_gnd_net_),
            .in2(N__58873),
            .in3(N__58584),
            .lcout(front_order_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94295),
            .ce(N__60020),
            .sr(N__59950));
    defparam \pid_front.source_pid_1_esr_12_LC_12_22_7 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_esr_12_LC_12_22_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_esr_12_LC_12_22_7 .LUT_INIT=16'b1000100010001010;
    LogicCell40 \pid_front.source_pid_1_esr_12_LC_12_22_7  (
            .in0(N__58617),
            .in1(N__58871),
            .in2(N__58588),
            .in3(N__55713),
            .lcout(front_order_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94295),
            .ce(N__60020),
            .sr(N__59950));
    defparam \pid_front.error_p_reg_esr_RNIPC5D1_7_LC_12_23_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIPC5D1_7_LC_12_23_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIPC5D1_7_LC_12_23_0 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIPC5D1_7_LC_12_23_0  (
            .in0(N__55657),
            .in1(N__55651),
            .in2(_gnd_net_),
            .in3(N__75381),
            .lcout(\pid_front.error_p_reg_esr_RNIPC5D1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIGL6F_0_8_LC_12_23_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIGL6F_0_8_LC_12_23_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIGL6F_0_8_LC_12_23_1 .LUT_INIT=16'b0110001110011100;
    LogicCell40 \pid_front.error_p_reg_esr_RNIGL6F_0_8_LC_12_23_1  (
            .in0(N__94616),
            .in1(N__61254),
            .in2(N__55639),
            .in3(N__55620),
            .lcout(\pid_front.error_p_reg_esr_RNIGL6F_0Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNI6UN6_7_LC_12_23_2 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNI6UN6_7_LC_12_23_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNI6UN6_7_LC_12_23_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNI6UN6_7_LC_12_23_2  (
            .in0(_gnd_net_),
            .in1(N__55634),
            .in2(_gnd_net_),
            .in3(N__94615),
            .lcout(\pid_front.N_2364_i ),
            .ltout(\pid_front.N_2364_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIBG6F_7_LC_12_23_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIBG6F_7_LC_12_23_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIBG6F_7_LC_12_23_3 .LUT_INIT=16'b1010111100101011;
    LogicCell40 \pid_front.error_p_reg_esr_RNIBG6F_7_LC_12_23_3  (
            .in0(N__55893),
            .in1(N__59086),
            .in2(N__55660),
            .in3(N__81751),
            .lcout(\pid_front.error_p_reg_esr_RNIBG6FZ0Z_7 ),
            .ltout(\pid_front.error_p_reg_esr_RNIBG6FZ0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIS0F23_7_LC_12_23_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIS0F23_7_LC_12_23_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIS0F23_7_LC_12_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_p_reg_esr_RNIS0F23_7_LC_12_23_4  (
            .in0(N__58326),
            .in1(N__55650),
            .in2(N__55642),
            .in3(N__75380),
            .lcout(\pid_front.error_p_reg_esr_RNIS0F23Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_7_LC_12_23_5 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_7_LC_12_23_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_7_LC_12_23_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_7_LC_12_23_5  (
            .in0(N__94618),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prevZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94310),
            .ce(N__71786),
            .sr(N__71629));
    defparam \pid_front.error_p_reg_esr_RNIGL6F_8_LC_12_23_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIGL6F_8_LC_12_23_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIGL6F_8_LC_12_23_6 .LUT_INIT=16'b1111010101110001;
    LogicCell40 \pid_front.error_p_reg_esr_RNIGL6F_8_LC_12_23_6  (
            .in0(N__61255),
            .in1(N__55638),
            .in2(N__55624),
            .in3(N__94617),
            .lcout(\pid_front.error_p_reg_esr_RNIGL6FZ0Z_8 ),
            .ltout(\pid_front.error_p_reg_esr_RNIGL6FZ0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIV7CQ2_8_LC_12_23_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIV7CQ2_8_LC_12_23_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIV7CQ2_8_LC_12_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_p_reg_esr_RNIV7CQ2_8_LC_12_23_7  (
            .in0(N__58254),
            .in1(N__71290),
            .in2(N__55831),
            .in3(N__66920),
            .lcout(\pid_front.error_p_reg_esr_RNIV7CQ2Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNIMHT91_16_LC_12_24_1 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNIMHT91_16_LC_12_24_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNIMHT91_16_LC_12_24_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_front.pid_prereg_esr_RNIMHT91_16_LC_12_24_1  (
            .in0(N__58504),
            .in1(N__58495),
            .in2(N__58486),
            .in3(N__58513),
            .lcout(\pid_front.un11lto30_i_a2_3_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un11lto30_i_a2_3_c_RNO_LC_12_24_3 .C_ON=1'b0;
    defparam \pid_front.un11lto30_i_a2_3_c_RNO_LC_12_24_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.un11lto30_i_a2_3_c_RNO_LC_12_24_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_front.un11lto30_i_a2_3_c_RNO_LC_12_24_3  (
            .in0(N__58570),
            .in1(N__55792),
            .in2(N__58538),
            .in3(N__58606),
            .lcout(\pid_front.un11lto30_i_a2_2_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_14_LC_12_24_4 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_14_LC_12_24_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_14_LC_12_24_4 .LUT_INIT=16'b0011101011001010;
    LogicCell40 \pid_front.pid_prereg_14_LC_12_24_4  (
            .in0(N__55794),
            .in1(N__58948),
            .in2(N__70611),
            .in3(N__58549),
            .lcout(\pid_front.pid_preregZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94327),
            .ce(),
            .sr(N__86365));
    defparam \pid_front.pid_prereg_esr_RNIT5641_15_LC_12_24_5 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNIT5641_15_LC_12_24_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNIT5641_15_LC_12_24_5 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \pid_front.pid_prereg_esr_RNIT5641_15_LC_12_24_5  (
            .in0(N__58571),
            .in1(N__55793),
            .in2(N__58539),
            .in3(N__58607),
            .lcout(\pid_front.source_pid_9_i_0_o3_0_11 ),
            .ltout(\pid_front.source_pid_9_i_0_o3_0_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNIMQ9C6_30_LC_12_24_6 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNIMQ9C6_30_LC_12_24_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNIMQ9C6_30_LC_12_24_6 .LUT_INIT=16'b0101010101010000;
    LogicCell40 \pid_front.pid_prereg_esr_RNIMQ9C6_30_LC_12_24_6  (
            .in0(N__58862),
            .in1(_gnd_net_),
            .in2(N__55771),
            .in3(N__55768),
            .lcout(\pid_front.N_386 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI1VPN6_19_LC_12_25_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI1VPN6_19_LC_12_25_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI1VPN6_19_LC_12_25_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_front.error_p_reg_esr_RNI1VPN6_19_LC_12_25_0  (
            .in0(_gnd_net_),
            .in1(N__61065),
            .in2(_gnd_net_),
            .in3(N__61092),
            .lcout(\pid_front.error_p_reg_esr_RNI1VPN6Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIF0FB3_0_19_LC_12_25_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIF0FB3_0_19_LC_12_25_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIF0FB3_0_19_LC_12_25_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_p_reg_esr_RNIF0FB3_0_19_LC_12_25_1  (
            .in0(N__64188),
            .in1(N__70203),
            .in2(_gnd_net_),
            .in3(N__71432),
            .lcout(\pid_front.un1_pid_prereg_0_9 ),
            .ltout(\pid_front.un1_pid_prereg_0_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIQOPM6_18_LC_12_25_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIQOPM6_18_LC_12_25_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIQOPM6_18_LC_12_25_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIQOPM6_18_LC_12_25_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__55753),
            .in3(N__55950),
            .lcout(\pid_front.error_p_reg_esr_RNIQOPM6Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIF0FB3_19_LC_12_25_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIF0FB3_19_LC_12_25_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIF0FB3_19_LC_12_25_3 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIF0FB3_19_LC_12_25_3  (
            .in0(N__64189),
            .in1(N__70204),
            .in2(_gnd_net_),
            .in3(N__71433),
            .lcout(\pid_front.un1_pid_prereg_0_10 ),
            .ltout(\pid_front.un1_pid_prereg_0_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIRNJED_18_LC_12_25_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIRNJED_18_LC_12_25_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIRNJED_18_LC_12_25_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIRNJED_18_LC_12_25_4  (
            .in0(N__55951),
            .in1(N__55936),
            .in2(N__55954),
            .in3(N__61091),
            .lcout(\pid_front.error_p_reg_esr_RNIRNJEDZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIBOAB3_18_LC_12_25_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIBOAB3_18_LC_12_25_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIBOAB3_18_LC_12_25_5 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIBOAB3_18_LC_12_25_5  (
            .in0(N__72091),
            .in1(N__76147),
            .in2(_gnd_net_),
            .in3(N__72061),
            .lcout(\pid_front.un1_pid_prereg_0_8 ),
            .ltout(\pid_front.un1_pid_prereg_0_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI80EDD_17_LC_12_25_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI80EDD_17_LC_12_25_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI80EDD_17_LC_12_25_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_front.error_p_reg_esr_RNI80EDD_17_LC_12_25_6  (
            .in0(N__72034),
            .in1(N__72013),
            .in2(N__55939),
            .in3(N__55935),
            .lcout(\pid_front.error_p_reg_esr_RNI80EDDZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIIUAC3_0_20_LC_12_25_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIIUAC3_0_20_LC_12_25_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIIUAC3_0_20_LC_12_25_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIIUAC3_0_20_LC_12_25_7  (
            .in0(N__66621),
            .in1(N__64173),
            .in2(_gnd_net_),
            .in3(N__71397),
            .lcout(\pid_front.un1_pid_prereg_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNIIH1A1_24_LC_12_26_0 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNIIH1A1_24_LC_12_26_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNIIH1A1_24_LC_12_26_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_front.pid_prereg_esr_RNIIH1A1_24_LC_12_26_0  (
            .in0(N__58675),
            .in1(N__58684),
            .in2(N__58666),
            .in3(N__58693),
            .lcout(\pid_front.un11lto30_i_a2_5_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIBG6F_0_7_LC_12_26_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIBG6F_0_7_LC_12_26_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIBG6F_0_7_LC_12_26_3 .LUT_INIT=16'b0101101010010110;
    LogicCell40 \pid_front.error_p_reg_esr_RNIBG6F_0_7_LC_12_26_3  (
            .in0(N__55906),
            .in1(N__59079),
            .in2(N__55897),
            .in3(N__81726),
            .lcout(\pid_front.error_p_reg_esr_RNIBG6F_0Z0Z_7 ),
            .ltout(\pid_front.error_p_reg_esr_RNIBG6F_0Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI3K9L1_6_LC_12_26_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI3K9L1_6_LC_12_26_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI3K9L1_6_LC_12_26_4 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_front.error_p_reg_esr_RNI3K9L1_6_LC_12_26_4  (
            .in0(N__58816),
            .in1(_gnd_net_),
            .in2(N__55855),
            .in3(N__75450),
            .lcout(\pid_front.error_p_reg_esr_RNI3K9L1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNIN7IV_28_LC_12_26_7 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNIN7IV_28_LC_12_26_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNIN7IV_28_LC_12_26_7 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \pid_front.pid_prereg_esr_RNIN7IV_28_LC_12_26_7  (
            .in0(N__58839),
            .in1(N__58885),
            .in2(_gnd_net_),
            .in3(N__58894),
            .lcout(\pid_front.un11lto30_i_a2_6_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIQHN6_1_LC_12_27_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIQHN6_1_LC_12_27_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIQHN6_1_LC_12_27_1 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIQHN6_1_LC_12_27_1  (
            .in0(N__61364),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61336),
            .lcout(),
            .ltout(\pid_front.error_d_reg_prev_esr_RNIQHN6Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNID19M1_1_LC_12_27_2 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNID19M1_1_LC_12_27_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNID19M1_1_LC_12_27_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNID19M1_1_LC_12_27_2  (
            .in0(N__75568),
            .in1(N__63616),
            .in2(N__55981),
            .in3(N__61302),
            .lcout(\pid_front.error_d_reg_prev_esr_RNID19M1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI2BC9_1_LC_12_27_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI2BC9_1_LC_12_27_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI2BC9_1_LC_12_27_3 .LUT_INIT=16'b1111110011010100;
    LogicCell40 \pid_front.error_p_reg_esr_RNI2BC9_1_LC_12_27_3  (
            .in0(N__58987),
            .in1(N__61334),
            .in2(N__59040),
            .in3(N__58911),
            .lcout(\pid_front.error_p_reg_esr_RNI2BC9Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_0_LC_12_27_4 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_0_LC_12_27_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_0_LC_12_27_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_0_LC_12_27_4  (
            .in0(N__58913),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prevZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94366),
            .ce(N__71805),
            .sr(N__71707));
    defparam \pid_front.error_p_reg_esr_RNI2BC9_0_1_LC_12_27_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI2BC9_0_1_LC_12_27_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI2BC9_0_1_LC_12_27_5 .LUT_INIT=16'b1111001101110001;
    LogicCell40 \pid_front.error_p_reg_esr_RNI2BC9_0_1_LC_12_27_5  (
            .in0(N__58988),
            .in1(N__61335),
            .in2(N__59041),
            .in3(N__58912),
            .lcout(),
            .ltout(\pid_front.error_p_reg_esr_RNI2BC9_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIFSHO_1_LC_12_27_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIFSHO_1_LC_12_27_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIFSHO_1_LC_12_27_6 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIFSHO_1_LC_12_27_6  (
            .in0(_gnd_net_),
            .in1(N__61363),
            .in2(N__55978),
            .in3(N__55975),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIFSHOZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_1_LC_12_27_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_1_LC_12_27_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_1_LC_12_27_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_1_LC_12_27_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61337),
            .lcout(\pid_front.error_d_reg_prevZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94366),
            .ce(N__71805),
            .sr(N__71707));
    defparam \pid_front.error_p_reg_esr_6_LC_12_28_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_6_LC_12_28_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_6_LC_12_28_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_6_LC_12_28_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55969),
            .lcout(\pid_front.error_p_regZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94373),
            .ce(N__93317),
            .sr(N__93003));
    defparam \pid_side.un11lto30_i_a2_1_c_RNO_LC_13_2_0 .C_ON=1'b0;
    defparam \pid_side.un11lto30_i_a2_1_c_RNO_LC_13_2_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.un11lto30_i_a2_1_c_RNO_LC_13_2_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_side.un11lto30_i_a2_1_c_RNO_LC_13_2_0  (
            .in0(N__64598),
            .in1(N__64559),
            .in2(N__64525),
            .in3(N__64634),
            .lcout(\pid_side.un11lto30_i_a2_0_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIQGO21_14_LC_13_3_2 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIQGO21_14_LC_13_3_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIQGO21_14_LC_13_3_2 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIQGO21_14_LC_13_3_2  (
            .in0(N__61921),
            .in1(N__61936),
            .in2(_gnd_net_),
            .in3(N__62017),
            .lcout(),
            .ltout(\pid_side.error_i_acumm_13_i_o2_0_7_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNI5LOD5_0_13_LC_13_3_3 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNI5LOD5_0_13_LC_13_3_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNI5LOD5_0_13_LC_13_3_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNI5LOD5_0_13_LC_13_3_3  (
            .in0(N__60610),
            .in1(N__62131),
            .in2(N__56071),
            .in3(N__61906),
            .lcout(\pid_side.N_227 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNI0NAP5_12_LC_13_3_5 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNI0NAP5_12_LC_13_3_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNI0NAP5_12_LC_13_3_5 .LUT_INIT=16'b1101110111011101;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNI0NAP5_12_LC_13_3_5  (
            .in0(N__59782),
            .in1(N__61966),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.N_285 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNI22KG1_1_LC_13_4_1 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNI22KG1_1_LC_13_4_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNI22KG1_1_LC_13_4_1 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \pid_side.pid_prereg_esr_RNI22KG1_1_LC_13_4_1  (
            .in0(N__64659),
            .in1(N__64251),
            .in2(N__60753),
            .in3(N__64272),
            .lcout(),
            .ltout(\pid_side.un1_reset_i_a2_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNI7BMH5_0_LC_13_4_2 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNI7BMH5_0_LC_13_4_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNI7BMH5_0_LC_13_4_2 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \pid_side.pid_prereg_esr_RNI7BMH5_0_LC_13_4_2  (
            .in0(N__59353),
            .in1(N__59307),
            .in2(N__56068),
            .in3(N__62041),
            .lcout(),
            .ltout(\pid_side.N_342_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNIJUV5A_30_LC_13_4_3 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNIJUV5A_30_LC_13_4_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNIJUV5A_30_LC_13_4_3 .LUT_INIT=16'b1111000011111011;
    LogicCell40 \pid_side.pid_prereg_esr_RNIJUV5A_30_LC_13_4_3  (
            .in0(N__70966),
            .in1(N__59193),
            .in2(N__56065),
            .in3(N__59341),
            .lcout(\pid_side.un1_reset_0_i_3 ),
            .ltout(\pid_side.un1_reset_0_i_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.state_RNICOBCA_1_LC_13_4_4 .C_ON=1'b0;
    defparam \pid_side.state_RNICOBCA_1_LC_13_4_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.state_RNICOBCA_1_LC_13_4_4 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \pid_side.state_RNICOBCA_1_LC_13_4_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__56062),
            .in3(N__60743),
            .lcout(\pid_side.state_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.source_pid_1_esr_1_LC_13_4_5 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_esr_1_LC_13_4_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_esr_1_LC_13_4_5 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \pid_side.source_pid_1_esr_1_LC_13_4_5  (
            .in0(N__59237),
            .in1(N__59194),
            .in2(_gnd_net_),
            .in3(N__64273),
            .lcout(side_order_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94082),
            .ce(N__59141),
            .sr(N__59395));
    defparam \pid_side.source_pid_1_esr_2_LC_13_4_6 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_esr_2_LC_13_4_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_esr_2_LC_13_4_6 .LUT_INIT=16'b0000000000001010;
    LogicCell40 \pid_side.source_pid_1_esr_2_LC_13_4_6  (
            .in0(N__64252),
            .in1(_gnd_net_),
            .in2(N__59200),
            .in3(N__59241),
            .lcout(side_order_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94082),
            .ce(N__59141),
            .sr(N__59395));
    defparam \pid_side.source_pid_1_esr_3_LC_13_4_7 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_esr_3_LC_13_4_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_esr_3_LC_13_4_7 .LUT_INIT=16'b0000000000001010;
    LogicCell40 \pid_side.source_pid_1_esr_3_LC_13_4_7  (
            .in0(N__64660),
            .in1(_gnd_net_),
            .in2(N__59255),
            .in3(N__59198),
            .lcout(side_order_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94082),
            .ce(N__59141),
            .sr(N__59395));
    defparam \pid_side.state_RNIV8D6_0_LC_13_5_0 .C_ON=1'b0;
    defparam \pid_side.state_RNIV8D6_0_LC_13_5_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.state_RNIV8D6_0_LC_13_5_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pid_side.state_RNIV8D6_0_LC_13_5_0  (
            .in0(_gnd_net_),
            .in1(N__86582),
            .in2(_gnd_net_),
            .in3(N__60804),
            .lcout(\pid_side.state_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_14_LC_13_5_1 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_14_LC_13_5_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_14_LC_13_5_1 .LUT_INIT=16'b0011101011001010;
    LogicCell40 \pid_side.pid_prereg_14_LC_13_5_1  (
            .in0(N__62065),
            .in1(N__65350),
            .in2(N__60808),
            .in3(N__64768),
            .lcout(\pid_side.pid_preregZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94085),
            .ce(),
            .sr(N__86474));
    defparam \pid_side.un11lto30_i_a2_3_c_RNO_LC_13_5_2 .C_ON=1'b0;
    defparam \pid_side.un11lto30_i_a2_3_c_RNO_LC_13_5_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.un11lto30_i_a2_3_c_RNO_LC_13_5_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_side.un11lto30_i_a2_3_c_RNO_LC_13_5_2  (
            .in0(N__62056),
            .in1(N__64797),
            .in2(N__64756),
            .in3(N__64834),
            .lcout(\pid_side.un11lto30_i_a2_2_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNIDPVG_15_LC_13_5_3 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNIDPVG_15_LC_13_5_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNIDPVG_15_LC_13_5_3 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \pid_side.pid_prereg_esr_RNIDPVG_15_LC_13_5_3  (
            .in0(N__64835),
            .in1(N__64755),
            .in2(N__64804),
            .in3(N__62057),
            .lcout(\pid_side.source_pid_9_i_0_o3_0_11 ),
            .ltout(\pid_side.source_pid_9_i_0_o3_0_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNI6SNT_30_LC_13_5_4 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNI6SNT_30_LC_13_5_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNI6SNT_30_LC_13_5_4 .LUT_INIT=16'b0101010101010000;
    LogicCell40 \pid_side.pid_prereg_esr_RNI6SNT_30_LC_13_5_4  (
            .in0(N__65128),
            .in1(_gnd_net_),
            .in2(N__56329),
            .in3(N__62083),
            .lcout(\pid_side.N_386 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNI86E35_2_LC_13_5_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNI86E35_2_LC_13_5_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNI86E35_2_LC_13_5_6 .LUT_INIT=16'b0011001110011100;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_RNI86E35_2_LC_13_5_6  (
            .in0(N__56297),
            .in1(N__56152),
            .in2(N__56140),
            .in3(N__56125),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_0_axb_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNI1TA86_2_LC_13_5_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNI1TA86_2_LC_13_5_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNI1TA86_2_LC_13_5_7 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_RNI1TA86_2_LC_13_5_7  (
            .in0(_gnd_net_),
            .in1(N__56100),
            .in2(N__56086),
            .in3(_gnd_net_),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_RNI1TA86Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIGSJV_7_LC_13_6_1 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIGSJV_7_LC_13_6_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIGSJV_7_LC_13_6_1 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIGSJV_7_LC_13_6_1  (
            .in0(N__59492),
            .in1(N__59468),
            .in2(_gnd_net_),
            .in3(N__59426),
            .lcout(\pid_side.N_177 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIE2M21_12_LC_13_6_2 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIE2M21_12_LC_13_6_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIE2M21_12_LC_13_6_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIE2M21_12_LC_13_6_2  (
            .in0(_gnd_net_),
            .in1(N__59752),
            .in2(_gnd_net_),
            .in3(N__59451),
            .lcout(),
            .ltout(\pid_side.N_531_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIB8KB7_28_LC_13_6_3 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIB8KB7_28_LC_13_6_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIB8KB7_28_LC_13_6_3 .LUT_INIT=16'b1110111011101100;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIB8KB7_28_LC_13_6_3  (
            .in0(N__62792),
            .in1(N__60445),
            .in2(N__56350),
            .in3(N__61972),
            .lcout(\pid_side.N_255 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIEE6C1_5_LC_13_7_0 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIEE6C1_5_LC_13_7_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIEE6C1_5_LC_13_7_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIEE6C1_5_LC_13_7_0  (
            .in0(N__59816),
            .in1(N__59619),
            .in2(N__60332),
            .in3(N__59637),
            .lcout(\pid_side.N_603 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_6_LC_13_7_1 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_6_LC_13_7_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_6_LC_13_7_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_6_LC_13_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67852),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94095),
            .ce(N__65072),
            .sr(N__86460));
    defparam \pid_side.error_i_acumm_prereg_esr_5_LC_13_7_2 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_5_LC_13_7_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_5_LC_13_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_5_LC_13_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76059),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94095),
            .ce(N__65072),
            .sr(N__86460));
    defparam \pid_side.error_i_acumm_prereg_esr_11_LC_13_7_3 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_11_LC_13_7_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_11_LC_13_7_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_11_LC_13_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72566),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94095),
            .ce(N__65072),
            .sr(N__86460));
    defparam \pid_side.error_i_acumm_prereg_esr_10_LC_13_7_4 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_10_LC_13_7_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_10_LC_13_7_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_10_LC_13_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73180),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94095),
            .ce(N__65072),
            .sr(N__86460));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIJ04N_0_10_LC_13_7_5 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIJ04N_0_10_LC_13_7_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIJ04N_0_10_LC_13_7_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIJ04N_0_10_LC_13_7_5  (
            .in0(_gnd_net_),
            .in1(N__60322),
            .in2(_gnd_net_),
            .in3(N__59815),
            .lcout(\pid_side.N_544 ),
            .ltout(\pid_side.N_544_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIL12S6_12_LC_13_7_6 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIL12S6_12_LC_13_7_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIL12S6_12_LC_13_7_6 .LUT_INIT=16'b1010101011111011;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIL12S6_12_LC_13_7_6  (
            .in0(N__62769),
            .in1(N__59767),
            .in2(N__56347),
            .in3(N__59701),
            .lcout(\pid_side.error_i_acumm_13_i_0_tz_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_12_LC_13_7_7 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_12_LC_13_7_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_12_LC_13_7_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_12_LC_13_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68374),
            .lcout(\pid_side.un10lto12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94095),
            .ce(N__65072),
            .sr(N__86460));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIUU922_10_LC_13_8_0 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIUU922_10_LC_13_8_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIUU922_10_LC_13_8_0 .LUT_INIT=16'b0001111100001111;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIUU922_10_LC_13_8_0  (
            .in0(N__60326),
            .in1(N__59817),
            .in2(N__59768),
            .in3(N__56373),
            .lcout(\pid_side.N_181 ),
            .ltout(\pid_side.N_181_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_RNO_1_3_LC_13_8_1 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_RNO_1_3_LC_13_8_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_RNO_1_3_LC_13_8_1 .LUT_INIT=16'b0000000011110100;
    LogicCell40 \pid_side.error_i_acumm_RNO_1_3_LC_13_8_1  (
            .in0(N__59600),
            .in1(N__56394),
            .in2(N__56383),
            .in3(N__59700),
            .lcout(),
            .ltout(\pid_side.error_i_acumm_13_i_0_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_RNO_0_3_LC_13_8_2 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_RNO_0_3_LC_13_8_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_RNO_0_3_LC_13_8_2 .LUT_INIT=16'b1111111100010000;
    LogicCell40 \pid_side.error_i_acumm_RNO_0_3_LC_13_8_2  (
            .in0(N__62788),
            .in1(N__59667),
            .in2(N__56380),
            .in3(N__60452),
            .lcout(),
            .ltout(\pid_side.error_i_acumm_13_i_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_3_LC_13_8_3 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_3_LC_13_8_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_3_LC_13_8_3 .LUT_INIT=16'b0000101100001111;
    LogicCell40 \pid_side.error_i_acumm_3_LC_13_8_3  (
            .in0(N__59668),
            .in1(N__62789),
            .in2(N__56377),
            .in3(N__59915),
            .lcout(\pid_side.error_i_acummZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94102),
            .ce(N__60537),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNI3K2G7_12_LC_13_8_5 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNI3K2G7_12_LC_13_8_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNI3K2G7_12_LC_13_8_5 .LUT_INIT=16'b1111111101110000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNI3K2G7_12_LC_13_8_5  (
            .in0(N__56374),
            .in1(N__56362),
            .in2(N__59781),
            .in3(N__59699),
            .lcout(),
            .ltout(\pid_side.N_233_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIR48B8_28_LC_13_8_6 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIR48B8_28_LC_13_8_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIR48B8_28_LC_13_8_6 .LUT_INIT=16'b1111111101010000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIR48B8_28_LC_13_8_6  (
            .in0(N__62787),
            .in1(_gnd_net_),
            .in2(N__56356),
            .in3(N__60451),
            .lcout(\pid_side.N_251 ),
            .ltout(\pid_side.N_251_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_4_LC_13_8_7 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_4_LC_13_8_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_4_LC_13_8_7 .LUT_INIT=16'b0000101000001110;
    LogicCell40 \pid_side.error_i_acumm_4_LC_13_8_7  (
            .in0(N__59601),
            .in1(N__62790),
            .in2(N__56353),
            .in3(N__59916),
            .lcout(\pid_side.error_i_acummZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94102),
            .ce(N__60537),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_8_LC_13_9_0 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_8_LC_13_9_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_8_LC_13_9_0 .LUT_INIT=16'b0011001100010001;
    LogicCell40 \pid_side.error_i_acumm_8_LC_13_9_0  (
            .in0(N__59544),
            .in1(N__59562),
            .in2(_gnd_net_),
            .in3(N__59479),
            .lcout(\pid_side.error_i_acummZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94108),
            .ce(N__60549),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_9_LC_13_9_1 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_9_LC_13_9_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_9_LC_13_9_1 .LUT_INIT=16'b0000101000001111;
    LogicCell40 \pid_side.error_i_acumm_9_LC_13_9_1  (
            .in0(N__59500),
            .in1(_gnd_net_),
            .in2(N__59566),
            .in3(N__59545),
            .lcout(\pid_side.error_i_acummZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94108),
            .ce(N__60549),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_2_LC_13_9_2 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_2_LC_13_9_2 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_2_LC_13_9_2 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \uart_drone.data_Aux_RNO_0_2_LC_13_9_2  (
            .in0(N__56544),
            .in1(N__56479),
            .in2(_gnd_net_),
            .in3(N__56610),
            .lcout(\uart_drone.data_Auxce_0_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_3_LC_13_9_3 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_3_LC_13_9_3 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_3_LC_13_9_3 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \uart_drone.data_Aux_RNO_0_3_LC_13_9_3  (
            .in0(N__56611),
            .in1(_gnd_net_),
            .in2(N__56491),
            .in3(N__56545),
            .lcout(\uart_drone.data_Auxce_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_0_LC_13_10_2 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_0_LC_13_10_2 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_0_LC_13_10_2 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \uart_drone.data_Aux_RNO_0_0_LC_13_10_2  (
            .in0(N__56501),
            .in1(N__56564),
            .in2(_gnd_net_),
            .in3(N__56630),
            .lcout(\uart_drone.data_Auxce_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_1_LC_13_10_4 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_1_LC_13_10_4 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_1_LC_13_10_4 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \uart_drone.data_Aux_RNO_0_1_LC_13_10_4  (
            .in0(N__56502),
            .in1(N__56565),
            .in2(_gnd_net_),
            .in3(N__56631),
            .lcout(\uart_drone.data_Auxce_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_5_LC_13_10_7 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_5_LC_13_10_7 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_5_LC_13_10_7 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \uart_drone.data_Aux_RNO_0_5_LC_13_10_7  (
            .in0(N__56632),
            .in1(_gnd_net_),
            .in2(N__56569),
            .in3(N__56503),
            .lcout(\uart_drone.data_Auxce_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_0_LC_13_11_0 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_0_LC_13_11_0 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_0_LC_13_11_0 .LUT_INIT=16'b1010101011100010;
    LogicCell40 \uart_drone.data_Aux_0_LC_13_11_0  (
            .in0(N__56727),
            .in1(N__56446),
            .in2(N__56866),
            .in3(N__56901),
            .lcout(\uart_drone.data_AuxZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94125),
            .ce(),
            .sr(N__56743));
    defparam \uart_drone.data_Aux_1_LC_13_11_1 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_1_LC_13_11_1 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_1_LC_13_11_1 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \uart_drone.data_Aux_1_LC_13_11_1  (
            .in0(N__56902),
            .in1(N__56440),
            .in2(N__56715),
            .in3(N__56853),
            .lcout(\uart_drone.data_AuxZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94125),
            .ce(),
            .sr(N__56743));
    defparam \uart_drone.data_Aux_2_LC_13_11_2 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_2_LC_13_11_2 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_2_LC_13_11_2 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \uart_drone.data_Aux_2_LC_13_11_2  (
            .in0(N__56434),
            .in1(N__56694),
            .in2(N__56867),
            .in3(N__56903),
            .lcout(\uart_drone.data_AuxZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94125),
            .ce(),
            .sr(N__56743));
    defparam \uart_drone.data_Aux_3_LC_13_11_3 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_3_LC_13_11_3 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_3_LC_13_11_3 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \uart_drone.data_Aux_3_LC_13_11_3  (
            .in0(N__56904),
            .in1(N__56425),
            .in2(N__56682),
            .in3(N__56854),
            .lcout(\uart_drone.data_AuxZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94125),
            .ce(),
            .sr(N__56743));
    defparam \uart_drone.data_Aux_4_LC_13_11_4 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_4_LC_13_11_4 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_4_LC_13_11_4 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \uart_drone.data_Aux_4_LC_13_11_4  (
            .in0(N__56416),
            .in1(N__56661),
            .in2(N__56868),
            .in3(N__56905),
            .lcout(\uart_drone.data_AuxZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94125),
            .ce(),
            .sr(N__56743));
    defparam \uart_drone.data_Aux_5_LC_13_11_5 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_5_LC_13_11_5 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_5_LC_13_11_5 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \uart_drone.data_Aux_5_LC_13_11_5  (
            .in0(N__56906),
            .in1(N__56407),
            .in2(N__56649),
            .in3(N__56855),
            .lcout(\uart_drone.data_AuxZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94125),
            .ce(),
            .sr(N__56743));
    defparam \uart_drone.data_Aux_6_LC_13_11_6 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_6_LC_13_11_6 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_6_LC_13_11_6 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \uart_drone.data_Aux_6_LC_13_11_6  (
            .in0(N__56920),
            .in1(N__57003),
            .in2(N__56869),
            .in3(N__56907),
            .lcout(\uart_drone.data_AuxZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94125),
            .ce(),
            .sr(N__56743));
    defparam \uart_drone.data_Aux_7_LC_13_11_7 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_7_LC_13_11_7 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_7_LC_13_11_7 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \uart_drone.data_Aux_7_LC_13_11_7  (
            .in0(N__56908),
            .in1(N__56852),
            .in2(N__56991),
            .in3(N__56769),
            .lcout(\uart_drone.data_AuxZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94125),
            .ce(),
            .sr(N__56743));
    defparam \pid_side.error_i_reg_esr_RNO_4_27_LC_13_12_6 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_4_27_LC_13_12_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_4_27_LC_13_12_6 .LUT_INIT=16'b0000000100110001;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_4_27_LC_13_12_6  (
            .in0(N__76655),
            .in1(N__87804),
            .in2(N__84168),
            .in3(N__83676),
            .lcout(\pid_side.N_338 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_esr_0_LC_13_13_0 .C_ON=1'b0;
    defparam \uart_drone.data_esr_0_LC_13_13_0 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_0_LC_13_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_0_LC_13_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56731),
            .lcout(uart_drone_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94141),
            .ce(N__56974),
            .sr(N__56956));
    defparam \uart_drone.data_esr_1_LC_13_13_1 .C_ON=1'b0;
    defparam \uart_drone.data_esr_1_LC_13_13_1 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_1_LC_13_13_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart_drone.data_esr_1_LC_13_13_1  (
            .in0(N__56716),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(uart_drone_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94141),
            .ce(N__56974),
            .sr(N__56956));
    defparam \uart_drone.data_esr_2_LC_13_13_2 .C_ON=1'b0;
    defparam \uart_drone.data_esr_2_LC_13_13_2 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_2_LC_13_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_2_LC_13_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56698),
            .lcout(uart_drone_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94141),
            .ce(N__56974),
            .sr(N__56956));
    defparam \uart_drone.data_esr_3_LC_13_13_3 .C_ON=1'b0;
    defparam \uart_drone.data_esr_3_LC_13_13_3 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_3_LC_13_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_3_LC_13_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56683),
            .lcout(uart_drone_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94141),
            .ce(N__56974),
            .sr(N__56956));
    defparam \uart_drone.data_esr_4_LC_13_13_4 .C_ON=1'b0;
    defparam \uart_drone.data_esr_4_LC_13_13_4 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_4_LC_13_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_4_LC_13_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56665),
            .lcout(uart_drone_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94141),
            .ce(N__56974),
            .sr(N__56956));
    defparam \uart_drone.data_esr_5_LC_13_13_5 .C_ON=1'b0;
    defparam \uart_drone.data_esr_5_LC_13_13_5 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_5_LC_13_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_5_LC_13_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56650),
            .lcout(uart_drone_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94141),
            .ce(N__56974),
            .sr(N__56956));
    defparam \uart_drone.data_esr_6_LC_13_13_6 .C_ON=1'b0;
    defparam \uart_drone.data_esr_6_LC_13_13_6 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_6_LC_13_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_6_LC_13_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57007),
            .lcout(uart_drone_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94141),
            .ce(N__56974),
            .sr(N__56956));
    defparam \uart_drone.data_esr_7_LC_13_13_7 .C_ON=1'b0;
    defparam \uart_drone.data_esr_7_LC_13_13_7 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_7_LC_13_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_7_LC_13_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56992),
            .lcout(uart_drone_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94141),
            .ce(N__56974),
            .sr(N__56956));
    defparam \pid_front.error_cry_6_c_RNIGTNV2_LC_13_14_1 .C_ON=1'b0;
    defparam \pid_front.error_cry_6_c_RNIGTNV2_LC_13_14_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_6_c_RNIGTNV2_LC_13_14_1 .LUT_INIT=16'b0011000011101110;
    LogicCell40 \pid_front.error_cry_6_c_RNIGTNV2_LC_13_14_1  (
            .in0(N__74495),
            .in1(N__78510),
            .in2(N__74317),
            .in3(N__56938),
            .lcout(\pid_front.N_187 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_3_22_LC_13_14_2 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_3_22_LC_13_14_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_3_22_LC_13_14_2 .LUT_INIT=16'b0001010110110101;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_3_22_LC_13_14_2  (
            .in0(N__82687),
            .in1(N__74300),
            .in2(N__90653),
            .in3(N__74494),
            .lcout(),
            .ltout(\pid_front.m26_2_03_0_m2_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_2_22_LC_13_14_3 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_2_22_LC_13_14_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_2_22_LC_13_14_3 .LUT_INIT=16'b0101111000001110;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_2_22_LC_13_14_3  (
            .in0(N__89066),
            .in1(N__73898),
            .in2(N__56932),
            .in3(N__78307),
            .lcout(\pid_front.N_297 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_2_23_LC_13_14_4 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_2_23_LC_13_14_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_2_23_LC_13_14_4 .LUT_INIT=16'b0100010011110100;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_2_23_LC_13_14_4  (
            .in0(N__73899),
            .in1(N__76955),
            .in2(N__76981),
            .in3(N__80659),
            .lcout(),
            .ltout(\pid_front.m27_2_03_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_0_23_LC_13_14_5 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_23_LC_13_14_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_23_LC_13_14_5 .LUT_INIT=16'b1111000011111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_23_LC_13_14_5  (
            .in0(_gnd_net_),
            .in1(N__73279),
            .in2(N__56929),
            .in3(N__56926),
            .lcout(\pid_front.m27_2_03_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_1_23_LC_13_14_6 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_1_23_LC_13_14_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_1_23_LC_13_14_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_1_23_LC_13_14_6  (
            .in0(N__78306),
            .in1(N__89065),
            .in2(_gnd_net_),
            .in3(N__74304),
            .lcout(\pid_front.N_253 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_7_LC_13_15_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_7_LC_13_15_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_7_LC_13_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_7_LC_13_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57781),
            .lcout(\dron_frame_decoder_1.drone_H_disp_front_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94165),
            .ce(N__57418),
            .sr(N__86426));
    defparam \pid_side.error_i_acumm_prereg_esr_0_LC_13_16_0 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_0_LC_13_16_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_0_LC_13_16_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_0_LC_13_16_0  (
            .in0(_gnd_net_),
            .in1(N__63016),
            .in2(_gnd_net_),
            .in3(N__62461),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94178),
            .ce(N__65080),
            .sr(N__86416));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNINAV3_7_LC_13_16_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNINAV3_7_LC_13_16_1 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNINAV3_7_LC_13_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_RNINAV3_7_LC_13_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57049),
            .lcout(drone_H_disp_front_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIOBV3_8_LC_13_16_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIOBV3_8_LC_13_16_2 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIOBV3_8_LC_13_16_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_RNIOBV3_8_LC_13_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57664),
            .lcout(drone_H_disp_front_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIPCV3_9_LC_13_16_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIPCV3_9_LC_13_16_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIPCV3_9_LC_13_16_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_RNIPCV3_9_LC_13_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57022),
            .lcout(drone_H_disp_front_i_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNI08RD_13_LC_13_16_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNI08RD_13_LC_13_16_4 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNI08RD_13_LC_13_16_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_RNI08RD_13_LC_13_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77427),
            .lcout(drone_H_disp_side_i_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIG6P4_4_LC_13_16_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIG6P4_4_LC_13_16_5 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIG6P4_4_LC_13_16_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_RNIG6P4_4_LC_13_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57172),
            .lcout(drone_H_disp_side_i_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIH7P4_5_LC_13_16_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIH7P4_5_LC_13_16_6 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIH7P4_5_LC_13_16_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_RNIH7P4_5_LC_13_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57166),
            .lcout(drone_H_disp_side_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNII8P4_6_LC_13_16_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNII8P4_6_LC_13_16_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNII8P4_6_LC_13_16_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_RNII8P4_6_LC_13_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57082),
            .lcout(drone_H_disp_side_i_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_0_LC_13_17_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_0_LC_13_17_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_0_LC_13_17_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_0_LC_13_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57707),
            .lcout(drone_H_disp_side_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94192),
            .ce(N__57076),
            .sr(N__86404));
    defparam \dron_frame_decoder_1.source_H_disp_side_fast_esr_0_LC_13_17_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_fast_esr_0_LC_13_17_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_fast_esr_0_LC_13_17_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_fast_esr_0_LC_13_17_1  (
            .in0(N__57708),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(dron_frame_decoder_1_source_H_disp_side_fast_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94192),
            .ce(N__57076),
            .sr(N__86404));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_1_LC_13_17_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_1_LC_13_17_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_1_LC_13_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_1_LC_13_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57327),
            .lcout(drone_H_disp_side_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94192),
            .ce(N__57076),
            .sr(N__86404));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_2_LC_13_17_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_2_LC_13_17_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_2_LC_13_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_2_LC_13_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57226),
            .lcout(drone_H_disp_side_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94192),
            .ce(N__57076),
            .sr(N__86404));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_3_LC_13_17_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_3_LC_13_17_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_3_LC_13_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_3_LC_13_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58011),
            .lcout(drone_H_disp_side_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94192),
            .ce(N__57076),
            .sr(N__86404));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_4_LC_13_17_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_4_LC_13_17_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_4_LC_13_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_4_LC_13_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57947),
            .lcout(\dron_frame_decoder_1.drone_H_disp_side_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94192),
            .ce(N__57076),
            .sr(N__86404));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_5_LC_13_17_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_5_LC_13_17_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_5_LC_13_17_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_5_LC_13_17_6  (
            .in0(N__57874),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\dron_frame_decoder_1.drone_H_disp_side_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94192),
            .ce(N__57076),
            .sr(N__86404));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_6_LC_13_17_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_6_LC_13_17_7 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_6_LC_13_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_6_LC_13_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57150),
            .lcout(\dron_frame_decoder_1.drone_H_disp_side_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94192),
            .ce(N__57076),
            .sr(N__86404));
    defparam \pid_front.error_cry_3_0_c_RNI3DE21_LC_13_18_0 .C_ON=1'b0;
    defparam \pid_front.error_cry_3_0_c_RNI3DE21_LC_13_18_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_3_0_c_RNI3DE21_LC_13_18_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \pid_front.error_cry_3_0_c_RNI3DE21_LC_13_18_0  (
            .in0(N__79655),
            .in1(N__84628),
            .in2(_gnd_net_),
            .in3(N__74791),
            .lcout(\pid_front.N_156 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_6_12_LC_13_18_1 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_6_12_LC_13_18_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_6_12_LC_13_18_1 .LUT_INIT=16'b0001010110110101;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_6_12_LC_13_18_1  (
            .in0(N__90412),
            .in1(N__82859),
            .in2(N__79660),
            .in3(N__81112),
            .lcout(),
            .ltout(\pid_side.error_i_reg_esr_RNO_6Z0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_4_12_LC_13_18_2 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_4_12_LC_13_18_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_4_12_LC_13_18_2 .LUT_INIT=16'b0100111101001010;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_4_12_LC_13_18_2  (
            .in0(N__78514),
            .in1(N__81647),
            .in2(N__57052),
            .in3(N__81534),
            .lcout(\pid_side.N_228_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_0_LC_13_18_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_0_LC_13_18_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_0_LC_13_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_0_LC_13_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57709),
            .lcout(drone_H_disp_front_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94207),
            .ce(N__57412),
            .sr(N__86395));
    defparam \dron_frame_decoder_1.source_H_disp_front_fast_esr_0_LC_13_18_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_fast_esr_0_LC_13_18_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_fast_esr_0_LC_13_18_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_fast_esr_0_LC_13_18_4  (
            .in0(N__57710),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(dron_frame_decoder_1_source_H_disp_front_fast_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94207),
            .ce(N__57412),
            .sr(N__86395));
    defparam \pid_side.error_i_reg_esr_RNO_4_16_LC_13_18_5 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_4_16_LC_13_18_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_4_16_LC_13_18_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_4_16_LC_13_18_5  (
            .in0(N__86938),
            .in1(N__89098),
            .in2(N__89821),
            .in3(N__84543),
            .lcout(\pid_side.error_i_reg_9_1_sn_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_0_18_LC_13_18_6 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_18_LC_13_18_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_18_LC_13_18_6 .LUT_INIT=16'b0010001001010101;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_18_LC_13_18_6  (
            .in0(N__84545),
            .in1(N__89345),
            .in2(_gnd_net_),
            .in3(N__86940),
            .lcout(\pid_front.error_i_reg_9_1_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_15_LC_13_18_7 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_15_LC_13_18_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_15_LC_13_18_7 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_15_LC_13_18_7  (
            .in0(N__86939),
            .in1(N__84544),
            .in2(_gnd_net_),
            .in3(N__70252),
            .lcout(\pid_side.error_i_reg_9_rn_1_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_2_0_c_RNISPUJ1_LC_13_19_0 .C_ON=1'b0;
    defparam \pid_front.error_cry_2_0_c_RNISPUJ1_LC_13_19_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_2_0_c_RNISPUJ1_LC_13_19_0 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \pid_front.error_cry_2_0_c_RNISPUJ1_LC_13_19_0  (
            .in0(N__82277),
            .in1(N__77783),
            .in2(N__83185),
            .in3(N__77684),
            .lcout(\pid_front.N_510 ),
            .ltout(\pid_front.N_510_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_3_0_c_RNI7FBC3_LC_13_19_1 .C_ON=1'b0;
    defparam \pid_front.error_cry_3_0_c_RNI7FBC3_LC_13_19_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_3_0_c_RNI7FBC3_LC_13_19_1 .LUT_INIT=16'b0101010001010000;
    LogicCell40 \pid_front.error_cry_3_0_c_RNI7FBC3_LC_13_19_1  (
            .in0(N__84832),
            .in1(N__76895),
            .in2(N__57349),
            .in3(N__74839),
            .lcout(),
            .ltout(\pid_front.N_596_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_2_c_RNILUC3A_LC_13_19_2 .C_ON=1'b0;
    defparam \pid_front.error_cry_2_c_RNILUC3A_LC_13_19_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_2_c_RNILUC3A_LC_13_19_2 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \pid_front.error_cry_2_c_RNILUC3A_LC_13_19_2  (
            .in0(N__81334),
            .in1(N__66072),
            .in2(N__57346),
            .in3(N__57343),
            .lcout(\pid_front.m9_2_03_3_i_3 ),
            .ltout(\pid_front.m9_2_03_3_i_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_5_LC_13_19_3 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_5_LC_13_19_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_5_LC_13_19_3 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \pid_front.error_i_reg_5_LC_13_19_3  (
            .in0(N__63339),
            .in1(N__83380),
            .in2(N__57331),
            .in3(N__82130),
            .lcout(\pid_front.error_i_regZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94224),
            .ce(),
            .sr(N__86385));
    defparam \pid_front.error_cry_2_0_c_RNIAGTB1_LC_13_19_4 .C_ON=1'b0;
    defparam \pid_front.error_cry_2_0_c_RNIAGTB1_LC_13_19_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_2_0_c_RNIAGTB1_LC_13_19_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \pid_front.error_cry_2_0_c_RNIAGTB1_LC_13_19_4  (
            .in0(N__82276),
            .in1(N__77782),
            .in2(_gnd_net_),
            .in3(N__77683),
            .lcout(),
            .ltout(\pid_front.N_162_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_9_c_RNIUR1D2_LC_13_19_5 .C_ON=1'b0;
    defparam \pid_front.error_cry_9_c_RNIUR1D2_LC_13_19_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_9_c_RNIUR1D2_LC_13_19_5 .LUT_INIT=16'b0000110000101110;
    LogicCell40 \pid_front.error_cry_9_c_RNIUR1D2_LC_13_19_5  (
            .in0(N__83028),
            .in1(N__90252),
            .in2(N__58039),
            .in3(N__78281),
            .lcout(\pid_front.N_231 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_11_LC_13_20_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_11_LC_13_20_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_11_LC_13_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_11_LC_13_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58028),
            .lcout(drone_H_disp_front_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94241),
            .ce(N__57641),
            .sr(N__86378));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_12_LC_13_20_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_12_LC_13_20_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_12_LC_13_20_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_12_LC_13_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57940),
            .lcout(drone_H_disp_front_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94241),
            .ce(N__57641),
            .sr(N__86378));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_13_LC_13_20_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_13_LC_13_20_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_13_LC_13_20_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_13_LC_13_20_3  (
            .in0(N__57870),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(drone_H_disp_front_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94241),
            .ce(N__57641),
            .sr(N__86378));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_15_LC_13_20_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_15_LC_13_20_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_15_LC_13_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_15_LC_13_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57785),
            .lcout(drone_H_disp_front_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94241),
            .ce(N__57641),
            .sr(N__86378));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_8_LC_13_20_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_8_LC_13_20_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_8_LC_13_20_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_8_LC_13_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57711),
            .lcout(\dron_frame_decoder_1.drone_H_disp_front_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94241),
            .ce(N__57641),
            .sr(N__86378));
    defparam \pid_alt.error_i_acumm_esr_13_LC_13_21_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_esr_13_LC_13_21_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_esr_13_LC_13_21_0 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \pid_alt.error_i_acumm_esr_13_LC_13_21_0  (
            .in0(N__57616),
            .in1(N__57580),
            .in2(_gnd_net_),
            .in3(N__57562),
            .lcout(\pid_alt.error_i_acummZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94258),
            .ce(N__57526),
            .sr(N__57490));
    defparam \pid_front.error_axb_8_l_ofx_LC_13_21_1 .C_ON=1'b0;
    defparam \pid_front.error_axb_8_l_ofx_LC_13_21_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_axb_8_l_ofx_LC_13_21_1 .LUT_INIT=16'b1111010111110101;
    LogicCell40 \pid_front.error_axb_8_l_ofx_LC_13_21_1  (
            .in0(N__58123),
            .in1(_gnd_net_),
            .in2(N__58114),
            .in3(N__58086),
            .lcout(\pid_front.error_axb_8_l_ofx_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_axb_7_LC_13_21_2 .C_ON=1'b0;
    defparam \pid_front.error_axb_7_LC_13_21_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_axb_7_LC_13_21_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_front.error_axb_7_LC_13_21_2  (
            .in0(_gnd_net_),
            .in1(N__58122),
            .in2(_gnd_net_),
            .in3(N__58110),
            .lcout(\pid_front.error_axbZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNI3C23_12_LC_13_21_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNI3C23_12_LC_13_21_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNI3C23_12_LC_13_21_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_RNI3C23_12_LC_13_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58085),
            .lcout(drone_H_disp_front_i_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_2_c_RNIB1241_LC_13_21_4 .C_ON=1'b0;
    defparam \pid_front.error_cry_2_c_RNIB1241_LC_13_21_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_2_c_RNIB1241_LC_13_21_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \pid_front.error_cry_2_c_RNIB1241_LC_13_21_4  (
            .in0(N__82278),
            .in1(N__74052),
            .in2(_gnd_net_),
            .in3(N__79855),
            .lcout(\pid_front.N_232 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_2_c_RNIJVOR_LC_13_21_5 .C_ON=1'b0;
    defparam \pid_front.error_cry_2_c_RNIJVOR_LC_13_21_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_2_c_RNIJVOR_LC_13_21_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \pid_front.error_cry_2_c_RNIJVOR_LC_13_21_5  (
            .in0(N__74051),
            .in1(N__83178),
            .in2(_gnd_net_),
            .in3(N__82279),
            .lcout(\pid_front.N_524 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_esr_RNIETB61_13_LC_13_21_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_RNIETB61_13_LC_13_21_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_esr_RNIETB61_13_LC_13_21_6 .LUT_INIT=16'b1000100011101110;
    LogicCell40 \pid_front.error_d_reg_esr_RNIETB61_13_LC_13_21_6  (
            .in0(N__64362),
            .in1(N__67698),
            .in2(_gnd_net_),
            .in3(N__67647),
            .lcout(\pid_front.error_d_reg_esr_RNIETB61Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_esr_RNIETB61_1_13_LC_13_21_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_RNIETB61_1_13_LC_13_21_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_esr_RNIETB61_1_13_LC_13_21_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_front.error_d_reg_esr_RNIETB61_1_13_LC_13_21_7  (
            .in0(N__67648),
            .in1(_gnd_net_),
            .in2(N__67702),
            .in3(N__64363),
            .lcout(\pid_front.N_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNIGB2N_0_LC_13_22_0 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNIGB2N_0_LC_13_22_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNIGB2N_0_LC_13_22_0 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \pid_front.pid_prereg_esr_RNIGB2N_0_LC_13_22_0  (
            .in0(N__60285),
            .in1(N__58429),
            .in2(N__58618),
            .in3(N__58459),
            .lcout(\pid_front.un1_reset_i_a2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un11lto30_i_a2_0_c_RNO_LC_13_22_1 .C_ON=1'b0;
    defparam \pid_front.un11lto30_i_a2_0_c_RNO_LC_13_22_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.un11lto30_i_a2_0_c_RNO_LC_13_22_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_front.un11lto30_i_a2_0_c_RNO_LC_13_22_1  (
            .in0(N__58154),
            .in1(N__60239),
            .in2(N__60081),
            .in3(N__60284),
            .lcout(\pid_front.source_pid10lt4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNIIAAH_1_LC_13_22_2 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNIIAAH_1_LC_13_22_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNIIAAH_1_LC_13_22_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \pid_front.pid_prereg_esr_RNIIAAH_1_LC_13_22_2  (
            .in0(N__60240),
            .in1(N__60077),
            .in2(N__70469),
            .in3(N__58155),
            .lcout(\pid_front.un1_reset_i_a2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.state_1_LC_13_22_3 .C_ON=1'b0;
    defparam \pid_front.state_1_LC_13_22_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.state_1_LC_13_22_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.state_1_LC_13_22_3  (
            .in0(N__70558),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94277),
            .ce(),
            .sr(N__86369));
    defparam \pid_front.state_0_LC_13_22_4 .C_ON=1'b0;
    defparam \pid_front.state_0_LC_13_22_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.state_0_LC_13_22_4 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \pid_front.state_0_LC_13_22_4  (
            .in0(N__70447),
            .in1(N__70559),
            .in2(_gnd_net_),
            .in3(N__69150),
            .lcout(\pid_front.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94277),
            .ce(),
            .sr(N__86369));
    defparam \pid_front.state_RNIM14N_0_LC_13_22_5 .C_ON=1'b0;
    defparam \pid_front.state_RNIM14N_0_LC_13_22_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.state_RNIM14N_0_LC_13_22_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_front.state_RNIM14N_0_LC_13_22_5  (
            .in0(_gnd_net_),
            .in1(N__58177),
            .in2(_gnd_net_),
            .in3(N__93123),
            .lcout(\pid_front.state_RNIM14NZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.state_RNIPKTD_0_LC_13_22_6 .C_ON=1'b0;
    defparam \pid_front.state_RNIPKTD_0_LC_13_22_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.state_RNIPKTD_0_LC_13_22_6 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \pid_front.state_RNIPKTD_0_LC_13_22_6  (
            .in0(N__71018),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70557),
            .lcout(\pid_front.state_RNIPKTDZ0Z_0 ),
            .ltout(\pid_front.state_RNIPKTDZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.state_RNIFM151_0_LC_13_22_7 .C_ON=1'b0;
    defparam \pid_front.state_RNIFM151_0_LC_13_22_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.state_RNIFM151_0_LC_13_22_7 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \pid_front.state_RNIFM151_0_LC_13_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__58171),
            .in3(N__71627),
            .lcout(\pid_front.N_763_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_13_23_0 .C_ON=1'b1;
    defparam \pid_front.un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_13_23_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_13_23_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_front.un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_13_23_0  (
            .in0(_gnd_net_),
            .in1(N__67389),
            .in2(N__67393),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_23_0_),
            .carryout(\pid_front.un1_pid_prereg_0_cry_0_c_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_0_LC_13_23_1 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_0_LC_13_23_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_0_LC_13_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_0_LC_13_23_1  (
            .in0(_gnd_net_),
            .in1(N__58972),
            .in2(N__63213),
            .in3(N__58168),
            .lcout(\pid_front.pid_preregZ0Z_0 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_0_c_THRU_CO ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_0 ),
            .clk(N__94293),
            .ce(N__75320),
            .sr(N__86366));
    defparam \pid_front.pid_prereg_esr_1_LC_13_23_2 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_1_LC_13_23_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_1_LC_13_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_1_LC_13_23_2  (
            .in0(_gnd_net_),
            .in1(N__75614),
            .in2(N__59017),
            .in3(N__58141),
            .lcout(\pid_front.pid_preregZ0Z_1 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_0 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_1 ),
            .clk(N__94293),
            .ce(N__75320),
            .sr(N__86366));
    defparam \pid_front.pid_prereg_esr_2_LC_13_23_3 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_2_LC_13_23_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_2_LC_13_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_2_LC_13_23_3  (
            .in0(_gnd_net_),
            .in1(N__58138),
            .in2(N__75564),
            .in3(N__58126),
            .lcout(\pid_front.pid_preregZ0Z_2 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_1 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_2 ),
            .clk(N__94293),
            .ce(N__75320),
            .sr(N__86366));
    defparam \pid_front.pid_prereg_esr_3_LC_13_23_4 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_3_LC_13_23_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_3_LC_13_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_3_LC_13_23_4  (
            .in0(_gnd_net_),
            .in1(N__61290),
            .in2(N__61387),
            .in3(N__58474),
            .lcout(\pid_front.pid_preregZ0Z_3 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_2 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_3 ),
            .clk(N__94293),
            .ce(N__75320),
            .sr(N__86366));
    defparam \pid_front.pid_prereg_esr_4_LC_13_23_5 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_4_LC_13_23_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_4_LC_13_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_4_LC_13_23_5  (
            .in0(_gnd_net_),
            .in1(N__61165),
            .in2(N__61444),
            .in3(N__58438),
            .lcout(\pid_front.pid_preregZ0Z_4 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_3 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_4 ),
            .clk(N__94293),
            .ce(N__75320),
            .sr(N__86366));
    defparam \pid_front.pid_prereg_esr_5_LC_13_23_6 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_5_LC_13_23_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_5_LC_13_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_5_LC_13_23_6  (
            .in0(_gnd_net_),
            .in1(N__61633),
            .in2(N__61186),
            .in3(N__58408),
            .lcout(\pid_front.pid_preregZ0Z_5 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_4 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_5 ),
            .clk(N__94293),
            .ce(N__75320),
            .sr(N__86366));
    defparam \pid_front.pid_prereg_esr_6_LC_13_23_7 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_6_LC_13_23_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_6_LC_13_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_6_LC_13_23_7  (
            .in0(_gnd_net_),
            .in1(N__61726),
            .in2(N__61507),
            .in3(N__58372),
            .lcout(\pid_front.pid_preregZ0Z_6 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_5 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_6 ),
            .clk(N__94293),
            .ce(N__75320),
            .sr(N__86366));
    defparam \pid_front.pid_prereg_esr_7_LC_13_24_0 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_7_LC_13_24_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_7_LC_13_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_7_LC_13_24_0  (
            .in0(_gnd_net_),
            .in1(N__58801),
            .in2(N__61753),
            .in3(N__58330),
            .lcout(\pid_front.pid_preregZ0Z_7 ),
            .ltout(),
            .carryin(bfn_13_24_0_),
            .carryout(\pid_front.un1_pid_prereg_0_cry_7 ),
            .clk(N__94308),
            .ce(N__75318),
            .sr(N__86361));
    defparam \pid_front.pid_prereg_esr_8_LC_13_24_1 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_8_LC_13_24_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_8_LC_13_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_8_LC_13_24_1  (
            .in0(_gnd_net_),
            .in1(N__58327),
            .in2(N__58306),
            .in3(N__58264),
            .lcout(\pid_front.pid_preregZ0Z_8 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_7 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_8 ),
            .clk(N__94308),
            .ce(N__75318),
            .sr(N__86361));
    defparam \pid_front.pid_prereg_esr_9_LC_13_24_2 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_9_LC_13_24_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_9_LC_13_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_9_LC_13_24_2  (
            .in0(_gnd_net_),
            .in1(N__58261),
            .in2(N__58255),
            .in3(N__58210),
            .lcout(\pid_front.pid_preregZ0Z_9 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_8 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_9 ),
            .clk(N__94308),
            .ce(N__75318),
            .sr(N__86361));
    defparam \pid_front.pid_prereg_esr_10_LC_13_24_3 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_10_LC_13_24_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_10_LC_13_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_10_LC_13_24_3  (
            .in0(_gnd_net_),
            .in1(N__70345),
            .in2(N__70369),
            .in3(N__58180),
            .lcout(\pid_front.pid_preregZ0Z_10 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_9 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_10 ),
            .clk(N__94308),
            .ce(N__75318),
            .sr(N__86361));
    defparam \pid_front.pid_prereg_esr_11_LC_13_24_4 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_11_LC_13_24_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_11_LC_13_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_11_LC_13_24_4  (
            .in0(_gnd_net_),
            .in1(N__70314),
            .in2(N__70297),
            .in3(N__58621),
            .lcout(\pid_front.pid_preregZ0Z_11 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_10 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_11 ),
            .clk(N__94308),
            .ce(N__75318),
            .sr(N__86361));
    defparam \pid_front.pid_prereg_esr_12_LC_13_24_5 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_12_LC_13_24_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_12_LC_13_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_12_LC_13_24_5  (
            .in0(_gnd_net_),
            .in1(N__61612),
            .in2(N__61264),
            .in3(N__58591),
            .lcout(\pid_front.pid_preregZ0Z_12 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_11 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_12 ),
            .clk(N__94308),
            .ce(N__75318),
            .sr(N__86361));
    defparam \pid_front.pid_prereg_esr_13_LC_13_24_6 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_13_LC_13_24_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_13_LC_13_24_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_13_LC_13_24_6  (
            .in0(_gnd_net_),
            .in1(N__64015),
            .in2(N__63928),
            .in3(N__58552),
            .lcout(\pid_front.pid_preregZ0Z_13 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_12 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_13 ),
            .clk(N__94308),
            .ce(N__75318),
            .sr(N__86361));
    defparam \pid_front.un1_pid_prereg_0_cry_13_THRU_LUT4_0_LC_13_24_7 .C_ON=1'b1;
    defparam \pid_front.un1_pid_prereg_0_cry_13_THRU_LUT4_0_LC_13_24_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_pid_prereg_0_cry_13_THRU_LUT4_0_LC_13_24_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.un1_pid_prereg_0_cry_13_THRU_LUT4_0_LC_13_24_7  (
            .in0(_gnd_net_),
            .in1(N__58944),
            .in2(_gnd_net_),
            .in3(N__58543),
            .lcout(\pid_front.un1_pid_prereg_0_cry_13_THRU_CO ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_13 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_15_LC_13_25_0 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_15_LC_13_25_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_15_LC_13_25_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_15_LC_13_25_0  (
            .in0(_gnd_net_),
            .in1(N__71530),
            .in2(N__71595),
            .in3(N__58516),
            .lcout(\pid_front.pid_preregZ0Z_15 ),
            .ltout(),
            .carryin(bfn_13_25_0_),
            .carryout(\pid_front.un1_pid_prereg_0_cry_15 ),
            .clk(N__94326),
            .ce(N__75317),
            .sr(N__86359));
    defparam \pid_front.pid_prereg_esr_16_LC_13_25_1 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_16_LC_13_25_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_16_LC_13_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_16_LC_13_25_1  (
            .in0(_gnd_net_),
            .in1(N__68896),
            .in2(N__61456),
            .in3(N__58507),
            .lcout(\pid_front.pid_preregZ0Z_16 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_15 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_16 ),
            .clk(N__94326),
            .ce(N__75317),
            .sr(N__86359));
    defparam \pid_front.pid_prereg_esr_17_LC_13_25_2 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_17_LC_13_25_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_17_LC_13_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_17_LC_13_25_2  (
            .in0(_gnd_net_),
            .in1(N__61483),
            .in2(N__61495),
            .in3(N__58498),
            .lcout(\pid_front.pid_preregZ0Z_17 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_16 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_17 ),
            .clk(N__94326),
            .ce(N__75317),
            .sr(N__86359));
    defparam \pid_front.pid_prereg_esr_18_LC_13_25_3 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_18_LC_13_25_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_18_LC_13_25_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_18_LC_13_25_3  (
            .in0(_gnd_net_),
            .in1(N__63817),
            .in2(N__61528),
            .in3(N__58489),
            .lcout(\pid_front.pid_preregZ0Z_18 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_17 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_18 ),
            .clk(N__94326),
            .ce(N__75317),
            .sr(N__86359));
    defparam \pid_front.pid_prereg_esr_19_LC_13_25_4 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_19_LC_13_25_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_19_LC_13_25_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_19_LC_13_25_4  (
            .in0(_gnd_net_),
            .in1(N__63898),
            .in2(N__63916),
            .in3(N__58477),
            .lcout(\pid_front.pid_preregZ0Z_19 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_18 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_19 ),
            .clk(N__94326),
            .ce(N__75317),
            .sr(N__86359));
    defparam \pid_front.pid_prereg_esr_20_LC_13_25_5 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_20_LC_13_25_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_20_LC_13_25_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_20_LC_13_25_5  (
            .in0(_gnd_net_),
            .in1(N__58789),
            .in2(N__71995),
            .in3(N__58771),
            .lcout(\pid_front.pid_preregZ0Z_20 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_19 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_20 ),
            .clk(N__94326),
            .ce(N__75317),
            .sr(N__86359));
    defparam \pid_front.pid_prereg_esr_21_LC_13_25_6 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_21_LC_13_25_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_21_LC_13_25_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_21_LC_13_25_6  (
            .in0(_gnd_net_),
            .in1(N__58768),
            .in2(N__58762),
            .in3(N__58738),
            .lcout(\pid_front.pid_preregZ0Z_21 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_20 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_21 ),
            .clk(N__94326),
            .ce(N__75317),
            .sr(N__86359));
    defparam \pid_front.pid_prereg_esr_22_LC_13_25_7 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_22_LC_13_25_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_22_LC_13_25_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_22_LC_13_25_7  (
            .in0(_gnd_net_),
            .in1(N__61054),
            .in2(N__58735),
            .in3(N__58714),
            .lcout(\pid_front.pid_preregZ0Z_22 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_21 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_22 ),
            .clk(N__94326),
            .ce(N__75317),
            .sr(N__86359));
    defparam \pid_front.pid_prereg_esr_23_LC_13_26_0 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_23_LC_13_26_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_23_LC_13_26_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_23_LC_13_26_0  (
            .in0(_gnd_net_),
            .in1(N__61042),
            .in2(N__61231),
            .in3(N__58696),
            .lcout(\pid_front.pid_preregZ0Z_23 ),
            .ltout(),
            .carryin(bfn_13_26_0_),
            .carryout(\pid_front.un1_pid_prereg_0_cry_23 ),
            .clk(N__94341),
            .ce(N__75316),
            .sr(N__86357));
    defparam \pid_front.pid_prereg_esr_24_LC_13_26_1 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_24_LC_13_26_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_24_LC_13_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_24_LC_13_26_1  (
            .in0(_gnd_net_),
            .in1(N__61534),
            .in2(N__61201),
            .in3(N__58687),
            .lcout(\pid_front.pid_preregZ0Z_24 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_23 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_24 ),
            .clk(N__94341),
            .ce(N__75316),
            .sr(N__86357));
    defparam \pid_front.pid_prereg_esr_25_LC_13_26_2 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_25_LC_13_26_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_25_LC_13_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_25_LC_13_26_2  (
            .in0(_gnd_net_),
            .in1(N__61591),
            .in2(N__61603),
            .in3(N__58678),
            .lcout(\pid_front.pid_preregZ0Z_25 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_24 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_25 ),
            .clk(N__94341),
            .ce(N__75316),
            .sr(N__86357));
    defparam \pid_front.pid_prereg_esr_26_LC_13_26_3 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_26_LC_13_26_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_26_LC_13_26_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_26_LC_13_26_3  (
            .in0(_gnd_net_),
            .in1(N__61813),
            .in2(N__61516),
            .in3(N__58669),
            .lcout(\pid_front.pid_preregZ0Z_26 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_25 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_26 ),
            .clk(N__94341),
            .ce(N__75316),
            .sr(N__86357));
    defparam \pid_front.pid_prereg_esr_27_LC_13_26_4 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_27_LC_13_26_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_27_LC_13_26_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_27_LC_13_26_4  (
            .in0(_gnd_net_),
            .in1(N__61867),
            .in2(N__61879),
            .in3(N__58657),
            .lcout(\pid_front.pid_preregZ0Z_27 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_26 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_27 ),
            .clk(N__94341),
            .ce(N__75316),
            .sr(N__86357));
    defparam \pid_front.pid_prereg_esr_28_LC_13_26_5 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_28_LC_13_26_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_28_LC_13_26_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_28_LC_13_26_5  (
            .in0(_gnd_net_),
            .in1(N__66721),
            .in2(N__61804),
            .in3(N__58888),
            .lcout(\pid_front.pid_preregZ0Z_28 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_27 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_28 ),
            .clk(N__94341),
            .ce(N__75316),
            .sr(N__86357));
    defparam \pid_front.pid_prereg_esr_29_LC_13_26_6 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_29_LC_13_26_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_29_LC_13_26_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_29_LC_13_26_6  (
            .in0(_gnd_net_),
            .in1(N__66847),
            .in2(N__66877),
            .in3(N__58879),
            .lcout(\pid_front.pid_preregZ0Z_29 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_28 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_29 ),
            .clk(N__94341),
            .ce(N__75316),
            .sr(N__86357));
    defparam \pid_front.pid_prereg_esr_30_LC_13_26_7 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_30_LC_13_26_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_30_LC_13_26_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_front.pid_prereg_esr_30_LC_13_26_7  (
            .in0(_gnd_net_),
            .in1(N__66859),
            .in2(_gnd_net_),
            .in3(N__58876),
            .lcout(\pid_front.pid_preregZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94341),
            .ce(N__75316),
            .sr(N__86357));
    defparam \pid_front.error_d_reg_prev_esr_RNI4SN6_6_LC_13_27_0 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNI4SN6_6_LC_13_27_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNI4SN6_6_LC_13_27_0 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNI4SN6_6_LC_13_27_0  (
            .in0(N__81743),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59078),
            .lcout(),
            .ltout(\pid_front.N_2358_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI6B6F_6_LC_13_27_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI6B6F_6_LC_13_27_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI6B6F_6_LC_13_27_1 .LUT_INIT=16'b1010111100101011;
    LogicCell40 \pid_front.error_p_reg_esr_RNI6B6F_6_LC_13_27_1  (
            .in0(N__61778),
            .in1(N__61708),
            .in2(N__58819),
            .in3(N__94664),
            .lcout(\pid_front.error_p_reg_esr_RNI6B6FZ0Z_6 ),
            .ltout(\pid_front.error_p_reg_esr_RNI6B6FZ0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI3K9L1_0_6_LC_13_27_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI3K9L1_0_6_LC_13_27_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI3K9L1_0_6_LC_13_27_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_p_reg_esr_RNI3K9L1_0_6_LC_13_27_2  (
            .in0(_gnd_net_),
            .in1(N__58810),
            .in2(N__58804),
            .in3(N__75451),
            .lcout(\pid_front.error_p_reg_esr_RNI3K9L1_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIMVC9_6_LC_13_27_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIMVC9_6_LC_13_27_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIMVC9_6_LC_13_27_5 .LUT_INIT=16'b1100001101101001;
    LogicCell40 \pid_front.error_p_reg_esr_RNIMVC9_6_LC_13_27_5  (
            .in0(N__61707),
            .in1(N__81742),
            .in2(N__61782),
            .in3(N__94663),
            .lcout(),
            .ltout(\pid_front.error_p_reg_esr_RNIMVC9Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNISAJO_6_LC_13_27_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNISAJO_6_LC_13_27_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNISAJO_6_LC_13_27_6 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNISAJO_6_LC_13_27_6  (
            .in0(_gnd_net_),
            .in1(N__59077),
            .in2(N__58792),
            .in3(N__61759),
            .lcout(\pid_front.error_d_reg_prev_esr_RNISAJOZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_6_LC_13_27_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_6_LC_13_27_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_6_LC_13_27_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_6_LC_13_27_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81744),
            .lcout(\pid_front.error_d_reg_prevZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94355),
            .ce(N__71787),
            .sr(N__71706));
    defparam \pid_front.error_p_reg_esr_1_LC_13_28_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_1_LC_13_28_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_1_LC_13_28_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_p_reg_esr_1_LC_13_28_0  (
            .in0(N__59059),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_p_regZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94365),
            .ce(N__93390),
            .sr(N__93004));
    defparam \pid_front.error_p_reg_esr_RNIL1E8_1_LC_13_28_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIL1E8_1_LC_13_28_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIL1E8_1_LC_13_28_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_p_reg_esr_RNIL1E8_1_LC_13_28_1  (
            .in0(N__61371),
            .in1(N__59039),
            .in2(_gnd_net_),
            .in3(N__61338),
            .lcout(),
            .ltout(\pid_front.un1_pid_prereg_9_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIMRLT_0_LC_13_28_2 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIMRLT_0_LC_13_28_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIMRLT_0_LC_13_28_2 .LUT_INIT=16'b0000111111000011;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIMRLT_0_LC_13_28_2  (
            .in0(N__75616),
            .in1(N__58990),
            .in2(N__59020),
            .in3(N__58915),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIMRLTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_esr_1_LC_13_28_3 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_1_LC_13_28_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_1_LC_13_28_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_1_LC_13_28_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59005),
            .lcout(\pid_front.error_d_regZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94365),
            .ce(N__93390),
            .sr(N__93004));
    defparam \pid_front.error_d_reg_prev_esr_RNIAHDK_0_LC_13_28_4 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIAHDK_0_LC_13_28_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIAHDK_0_LC_13_28_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIAHDK_0_LC_13_28_4  (
            .in0(N__63217),
            .in1(N__58989),
            .in2(_gnd_net_),
            .in3(N__58914),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIAHDKZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI6D5L7_12_LC_13_28_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI6D5L7_12_LC_13_28_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI6D5L7_12_LC_13_28_5 .LUT_INIT=16'b0110001111000110;
    LogicCell40 \pid_front.error_p_reg_esr_RNI6D5L7_12_LC_13_28_5  (
            .in0(N__58960),
            .in1(N__64318),
            .in2(N__78649),
            .in3(N__67180),
            .lcout(),
            .ltout(\pid_front.error_p_reg_esr_RNI6D5L7Z0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIV1EFE_12_LC_13_28_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIV1EFE_12_LC_13_28_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIV1EFE_12_LC_13_28_6 .LUT_INIT=16'b1001011001011010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIV1EFE_12_LC_13_28_6  (
            .in0(N__69957),
            .in1(N__64405),
            .in2(N__58951),
            .in3(N__67228),
            .lcout(\pid_front.un1_pid_prereg_0_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_esr_0_LC_13_28_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_0_LC_13_28_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_0_LC_13_28_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_0_LC_13_28_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58930),
            .lcout(\pid_front.error_d_regZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94365),
            .ce(N__93390),
            .sr(N__93004));
    defparam \pid_side.un11lto30_i_a2_0_c_LC_14_3_0 .C_ON=1'b1;
    defparam \pid_side.un11lto30_i_a2_0_c_LC_14_3_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.un11lto30_i_a2_0_c_LC_14_3_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_side.un11lto30_i_a2_0_c_LC_14_3_0  (
            .in0(_gnd_net_),
            .in1(N__64309),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_3_0_),
            .carryout(\pid_side.un11lto30_i_a2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un11lto30_i_a2_1_c_LC_14_3_1 .C_ON=1'b1;
    defparam \pid_side.un11lto30_i_a2_1_c_LC_14_3_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.un11lto30_i_a2_1_c_LC_14_3_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_side.un11lto30_i_a2_1_c_LC_14_3_1  (
            .in0(_gnd_net_),
            .in1(N__59110),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_side.un11lto30_i_a2 ),
            .carryout(\pid_side.un11lto30_i_a2_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un11lto30_i_a2_2_c_LC_14_3_2 .C_ON=1'b1;
    defparam \pid_side.un11lto30_i_a2_2_c_LC_14_3_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.un11lto30_i_a2_2_c_LC_14_3_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_side.un11lto30_i_a2_2_c_LC_14_3_2  (
            .in0(_gnd_net_),
            .in1(N__59266),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_side.un11lto30_i_a2_0 ),
            .carryout(\pid_side.un11lto30_i_a2_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un11lto30_i_a2_3_c_LC_14_3_3 .C_ON=1'b1;
    defparam \pid_side.un11lto30_i_a2_3_c_LC_14_3_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.un11lto30_i_a2_3_c_LC_14_3_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_side.un11lto30_i_a2_3_c_LC_14_3_3  (
            .in0(_gnd_net_),
            .in1(N__59104),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_side.un11lto30_i_a2_1 ),
            .carryout(\pid_side.un11lto30_i_a2_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un11lto30_i_a2_4_c_LC_14_3_4 .C_ON=1'b1;
    defparam \pid_side.un11lto30_i_a2_4_c_LC_14_3_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.un11lto30_i_a2_4_c_LC_14_3_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_side.un11lto30_i_a2_4_c_LC_14_3_4  (
            .in0(_gnd_net_),
            .in1(N__62233),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_side.un11lto30_i_a2_2 ),
            .carryout(\pid_side.un11lto30_i_a2_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un11lto30_i_a2_5_c_LC_14_3_5 .C_ON=1'b1;
    defparam \pid_side.un11lto30_i_a2_5_c_LC_14_3_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.un11lto30_i_a2_5_c_LC_14_3_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_side.un11lto30_i_a2_5_c_LC_14_3_5  (
            .in0(_gnd_net_),
            .in1(N__62218),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_side.un11lto30_i_a2_3 ),
            .carryout(\pid_side.un11lto30_i_a2_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un11lto30_i_a2_6_c_LC_14_3_6 .C_ON=1'b1;
    defparam \pid_side.un11lto30_i_a2_6_c_LC_14_3_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.un11lto30_i_a2_6_c_LC_14_3_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_side.un11lto30_i_a2_6_c_LC_14_3_6  (
            .in0(_gnd_net_),
            .in1(N__62095),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_side.un11lto30_i_a2_4 ),
            .carryout(\pid_side.un11lto30_i_a2_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un11lto30_i_a2_7_c_LC_14_3_7 .C_ON=1'b1;
    defparam \pid_side.un11lto30_i_a2_7_c_LC_14_3_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.un11lto30_i_a2_7_c_LC_14_3_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_side.un11lto30_i_a2_7_c_LC_14_3_7  (
            .in0(_gnd_net_),
            .in1(N__62248),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_side.un11lto30_i_a2_5 ),
            .carryout(\pid_side.un11lto30_i_a2_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un11lto30_i_a2_7_c_RNIA3131_LC_14_4_0 .C_ON=1'b0;
    defparam \pid_side.un11lto30_i_a2_7_c_RNIA3131_LC_14_4_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.un11lto30_i_a2_7_c_RNIA3131_LC_14_4_0 .LUT_INIT=16'b1110111011111111;
    LogicCell40 \pid_side.un11lto30_i_a2_7_c_RNIA3131_LC_14_4_0  (
            .in0(N__59095),
            .in1(N__62079),
            .in2(_gnd_net_),
            .in3(N__59089),
            .lcout(\pid_side.N_291 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNI0R0B1_0_LC_14_4_3 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNI0R0B1_0_LC_14_4_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNI0R0B1_0_LC_14_4_3 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \pid_side.pid_prereg_esr_RNI0R0B1_0_LC_14_4_3  (
            .in0(N__64628),
            .in1(N__64592),
            .in2(N__64843),
            .in3(N__64296),
            .lcout(\pid_side.un1_reset_i_a2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNIKRDJ1_30_LC_14_4_4 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNIKRDJ1_30_LC_14_4_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNIKRDJ1_30_LC_14_4_4 .LUT_INIT=16'b0001010100000101;
    LogicCell40 \pid_side.pid_prereg_esr_RNIKRDJ1_30_LC_14_4_4  (
            .in0(N__70965),
            .in1(N__65126),
            .in2(N__60752),
            .in3(N__59347),
            .lcout(\pid_side.un1_reset_i_o3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNIRALN2_4_LC_14_5_1 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNIRALN2_4_LC_14_5_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNIRALN2_4_LC_14_5_1 .LUT_INIT=16'b0101000001000000;
    LogicCell40 \pid_side.pid_prereg_esr_RNIRALN2_4_LC_14_5_1  (
            .in0(N__65127),
            .in1(N__64599),
            .in2(N__59308),
            .in3(N__64635),
            .lcout(\pid_side.N_631 ),
            .ltout(\pid_side.N_631_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.source_pid_1_esr_4_LC_14_5_2 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_esr_4_LC_14_5_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_esr_4_LC_14_5_2 .LUT_INIT=16'b1111111111111010;
    LogicCell40 \pid_side.source_pid_1_esr_4_LC_14_5_2  (
            .in0(N__64636),
            .in1(_gnd_net_),
            .in2(N__59335),
            .in3(N__59254),
            .lcout(side_order_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94093),
            .ce(N__59149),
            .sr(N__59409));
    defparam \pid_side.pid_prereg_esr_RNIB61B1_10_LC_14_5_3 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNIB61B1_10_LC_14_5_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNIB61B1_10_LC_14_5_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_side.pid_prereg_esr_RNIB61B1_10_LC_14_5_3  (
            .in0(N__64452),
            .in1(N__64425),
            .in2(N__64524),
            .in3(N__64563),
            .lcout(),
            .ltout(\pid_side.un1_reset_i_a2_3_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNIS3LQ1_11_LC_14_5_4 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNIS3LQ1_11_LC_14_5_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNIS3LQ1_11_LC_14_5_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_side.pid_prereg_esr_RNIS3LQ1_11_LC_14_5_4  (
            .in0(N__64801),
            .in1(N__64878),
            .in2(N__59311),
            .in3(N__64479),
            .lcout(\pid_side.N_593 ),
            .ltout(\pid_side.N_593_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.source_pid_1_esr_5_LC_14_5_5 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_esr_5_LC_14_5_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_esr_5_LC_14_5_5 .LUT_INIT=16'b0100010100000000;
    LogicCell40 \pid_side.source_pid_1_esr_5_LC_14_5_5  (
            .in0(N__59253),
            .in1(N__65129),
            .in2(N__59293),
            .in3(N__64600),
            .lcout(side_order_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94093),
            .ce(N__59149),
            .sr(N__59409));
    defparam \pid_side.un11lto30_i_a2_2_c_RNO_LC_14_5_6 .C_ON=1'b0;
    defparam \pid_side.un11lto30_i_a2_2_c_RNO_LC_14_5_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.un11lto30_i_a2_2_c_RNO_LC_14_5_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_side.un11lto30_i_a2_2_c_RNO_LC_14_5_6  (
            .in0(N__64424),
            .in1(N__64451),
            .in2(N__64877),
            .in3(N__64478),
            .lcout(\pid_side.N_11_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.source_pid_1_esr_0_LC_14_5_7 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_esr_0_LC_14_5_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_esr_0_LC_14_5_7 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \pid_side.source_pid_1_esr_0_LC_14_5_7  (
            .in0(N__59252),
            .in1(N__59199),
            .in2(_gnd_net_),
            .in3(N__64300),
            .lcout(side_order_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94093),
            .ce(N__59149),
            .sr(N__59409));
    defparam \pid_side.error_i_acumm_prereg_esr_17_LC_14_6_0 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_17_LC_14_6_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_17_LC_14_6_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_17_LC_14_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62611),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94099),
            .ce(N__65073),
            .sr(N__86461));
    defparam \pid_side.error_i_acumm_prereg_esr_1_LC_14_6_1 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_1_LC_14_6_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_1_LC_14_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_1_LC_14_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72329),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94099),
            .ce(N__65073),
            .sr(N__86461));
    defparam \pid_side.error_i_acumm_prereg_esr_2_LC_14_6_2 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_2_LC_14_6_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_2_LC_14_6_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_2_LC_14_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76439),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94099),
            .ce(N__65073),
            .sr(N__86461));
    defparam \pid_side.error_i_acumm_prereg_esr_3_LC_14_6_3 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_3_LC_14_6_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_3_LC_14_6_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_3_LC_14_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78959),
            .lcout(\pid_side.error_i_acumm16lto3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94099),
            .ce(N__65073),
            .sr(N__86461));
    defparam \pid_side.error_i_acumm_prereg_esr_4_LC_14_6_4 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_4_LC_14_6_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_4_LC_14_6_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_4_LC_14_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76354),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94099),
            .ce(N__65073),
            .sr(N__86461));
    defparam \pid_side.error_i_acumm_prereg_esr_7_LC_14_6_5 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_7_LC_14_6_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_7_LC_14_6_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_7_LC_14_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72272),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94099),
            .ce(N__65073),
            .sr(N__86461));
    defparam \pid_side.error_i_acumm_prereg_esr_8_LC_14_6_6 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_8_LC_14_6_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_8_LC_14_6_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_8_LC_14_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72198),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94099),
            .ce(N__65073),
            .sr(N__86461));
    defparam \pid_side.error_i_acumm_prereg_esr_9_LC_14_6_7 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_9_LC_14_6_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_9_LC_14_6_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_9_LC_14_6_7  (
            .in0(N__72407),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94099),
            .ce(N__65073),
            .sr(N__86461));
    defparam \pid_side.error_i_acumm_5_LC_14_7_0 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_5_LC_14_7_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_5_LC_14_7_0 .LUT_INIT=16'b0000000010111010;
    LogicCell40 \pid_side.error_i_acumm_5_LC_14_7_0  (
            .in0(N__59638),
            .in1(N__59922),
            .in2(N__62793),
            .in3(N__59361),
            .lcout(\pid_side.error_i_acummZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94105),
            .ce(N__60550),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_6_LC_14_7_1 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_6_LC_14_7_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_6_LC_14_7_1 .LUT_INIT=16'b0101010100000100;
    LogicCell40 \pid_side.error_i_acumm_6_LC_14_7_1  (
            .in0(N__59362),
            .in1(N__62783),
            .in2(N__59926),
            .in3(N__59618),
            .lcout(\pid_side.error_i_acummZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94105),
            .ce(N__60550),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIIN4A1_5_LC_14_7_2 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIIN4A1_5_LC_14_7_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIIN4A1_5_LC_14_7_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIIN4A1_5_LC_14_7_2  (
            .in0(N__59651),
            .in1(N__59636),
            .in2(N__59620),
            .in3(N__59596),
            .lcout(),
            .ltout(\pid_side.error_i_acumm_13_0_a2_2_2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIT8ES2_28_LC_14_7_3 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIT8ES2_28_LC_14_7_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIT8ES2_28_LC_14_7_3 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIT8ES2_28_LC_14_7_3  (
            .in0(N__62770),
            .in1(N__60449),
            .in2(N__59569),
            .in3(N__59450),
            .lcout(\pid_side.error_i_acumm_13_0_a2_2_4_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIJ04N_10_LC_14_7_4 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIJ04N_10_LC_14_7_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIJ04N_10_LC_14_7_4 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIJ04N_10_LC_14_7_4  (
            .in0(_gnd_net_),
            .in1(N__60321),
            .in2(_gnd_net_),
            .in3(N__59814),
            .lcout(\pid_side.N_217 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_7_LC_14_7_7 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_7_LC_14_7_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_7_LC_14_7_7 .LUT_INIT=16'b0101010100010001;
    LogicCell40 \pid_side.error_i_acumm_7_LC_14_7_7  (
            .in0(N__59561),
            .in1(N__59538),
            .in2(_gnd_net_),
            .in3(N__59430),
            .lcout(\pid_side.error_i_acummZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94105),
            .ce(N__60550),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_1_LC_14_8_0 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_1_LC_14_8_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_1_LC_14_8_0 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \pid_side.error_i_acumm_1_LC_14_8_0  (
            .in0(N__59844),
            .in1(N__59856),
            .in2(N__59527),
            .in3(N__59877),
            .lcout(\pid_side.error_i_acummZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94111),
            .ce(N__60536),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIR48B8_1_28_LC_14_8_1 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIR48B8_1_28_LC_14_8_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIR48B8_1_28_LC_14_8_1 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIR48B8_1_28_LC_14_8_1  (
            .in0(N__60450),
            .in1(N__59515),
            .in2(N__62791),
            .in3(N__59716),
            .lcout(),
            .ltout(\pid_side.N_483_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIT2FLG_28_LC_14_8_2 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIT2FLG_28_LC_14_8_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIT2FLG_28_LC_14_8_2 .LUT_INIT=16'b1111010111110000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIT2FLG_28_LC_14_8_2  (
            .in0(N__61968),
            .in1(_gnd_net_),
            .in2(N__59509),
            .in3(N__59506),
            .lcout(\pid_side.error_i_acumm_13_0_tz_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNI3TNM1_7_LC_14_8_3 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNI3TNM1_7_LC_14_8_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNI3TNM1_7_LC_14_8_3 .LUT_INIT=16'b0000111100001110;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNI3TNM1_7_LC_14_8_3  (
            .in0(N__59499),
            .in1(N__59475),
            .in2(N__59452),
            .in3(N__59431),
            .lcout(),
            .ltout(\pid_side.N_488_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNI3K2G7_0_12_LC_14_8_4 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNI3K2G7_0_12_LC_14_8_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNI3K2G7_0_12_LC_14_8_4 .LUT_INIT=16'b0101010101010000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNI3K2G7_0_12_LC_14_8_4  (
            .in0(N__61967),
            .in1(_gnd_net_),
            .in2(N__59929),
            .in3(N__59769),
            .lcout(\pid_side.N_601 ),
            .ltout(\pid_side.N_601_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIR48B8_0_28_LC_14_8_5 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIR48B8_0_28_LC_14_8_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIR48B8_0_28_LC_14_8_5 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIR48B8_0_28_LC_14_8_5  (
            .in0(N__62776),
            .in1(_gnd_net_),
            .in2(N__59902),
            .in3(N__60453),
            .lcout(\pid_side.N_484 ),
            .ltout(\pid_side.N_484_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_0_LC_14_8_6 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_0_LC_14_8_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_0_LC_14_8_6 .LUT_INIT=16'b1010101010101000;
    LogicCell40 \pid_side.error_i_acumm_0_LC_14_8_6  (
            .in0(N__59899),
            .in1(N__59843),
            .in2(N__59881),
            .in3(N__59855),
            .lcout(\pid_side.error_i_acummZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94111),
            .ce(N__60536),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_2_LC_14_8_7 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_2_LC_14_8_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_2_LC_14_8_7 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \pid_side.error_i_acumm_2_LC_14_8_7  (
            .in0(N__59878),
            .in1(N__59869),
            .in2(N__59860),
            .in3(N__59845),
            .lcout(\pid_side.error_i_acummZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94111),
            .ce(N__60536),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_RNO_0_10_LC_14_9_0 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_RNO_0_10_LC_14_9_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_RNO_0_10_LC_14_9_0 .LUT_INIT=16'b0000111100001011;
    LogicCell40 \pid_side.error_i_acumm_RNO_0_10_LC_14_9_0  (
            .in0(N__59785),
            .in1(N__59823),
            .in2(N__62771),
            .in3(N__59718),
            .lcout(),
            .ltout(\pid_side.N_355_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_10_LC_14_9_1 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_10_LC_14_9_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_10_LC_14_9_1 .LUT_INIT=16'b0000001100000010;
    LogicCell40 \pid_side.error_i_acumm_10_LC_14_9_1  (
            .in0(N__59824),
            .in1(N__60442),
            .in2(N__59791),
            .in3(N__60353),
            .lcout(\pid_side.error_i_acummZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94119),
            .ce(N__60541),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_RNO_0_12_LC_14_9_2 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_RNO_0_12_LC_14_9_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_RNO_0_12_LC_14_9_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pid_side.error_i_acumm_RNO_0_12_LC_14_9_2  (
            .in0(_gnd_net_),
            .in1(N__59783),
            .in2(_gnd_net_),
            .in3(N__59717),
            .lcout(),
            .ltout(\pid_side.N_242_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_12_LC_14_9_3 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_12_LC_14_9_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_12_LC_14_9_3 .LUT_INIT=16'b0001000001010000;
    LogicCell40 \pid_side.error_i_acumm_12_LC_14_9_3  (
            .in0(N__60443),
            .in1(N__62742),
            .in2(N__59788),
            .in3(N__60355),
            .lcout(\pid_side.error_i_acummZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94119),
            .ce(N__60541),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_RNO_0_11_LC_14_9_4 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_RNO_0_11_LC_14_9_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_RNO_0_11_LC_14_9_4 .LUT_INIT=16'b0000111100001101;
    LogicCell40 \pid_side.error_i_acumm_RNO_0_11_LC_14_9_4  (
            .in0(N__60333),
            .in1(N__59784),
            .in2(N__62772),
            .in3(N__59719),
            .lcout(),
            .ltout(\pid_side.N_353_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_11_LC_14_9_5 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_11_LC_14_9_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_11_LC_14_9_5 .LUT_INIT=16'b0000010100000100;
    LogicCell40 \pid_side.error_i_acumm_11_LC_14_9_5  (
            .in0(N__60444),
            .in1(N__60354),
            .in2(N__60337),
            .in3(N__60334),
            .lcout(\pid_side.error_i_acummZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94119),
            .ce(N__60541),
            .sr(_gnd_net_));
    defparam \pid_front.source_pid_1_esr_0_LC_14_10_0 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_esr_0_LC_14_10_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_esr_0_LC_14_10_0 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \pid_front.source_pid_1_esr_0_LC_14_10_0  (
            .in0(N__60131),
            .in1(N__60194),
            .in2(_gnd_net_),
            .in3(N__60298),
            .lcout(front_order_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94129),
            .ce(N__60040),
            .sr(N__59995));
    defparam \pid_front.source_pid_1_esr_2_LC_14_10_2 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_esr_2_LC_14_10_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_esr_2_LC_14_10_2 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \pid_front.source_pid_1_esr_2_LC_14_10_2  (
            .in0(N__60132),
            .in1(N__60195),
            .in2(_gnd_net_),
            .in3(N__60250),
            .lcout(front_order_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94129),
            .ce(N__60040),
            .sr(N__59995));
    defparam \pid_front.source_pid_1_esr_3_LC_14_10_3 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_esr_3_LC_14_10_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_esr_3_LC_14_10_3 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \pid_front.source_pid_1_esr_3_LC_14_10_3  (
            .in0(N__60196),
            .in1(N__60133),
            .in2(_gnd_net_),
            .in3(N__60091),
            .lcout(front_order_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94129),
            .ce(N__60040),
            .sr(N__59995));
    defparam \pid_side.error_d_reg_fast_esr_RNIFGGE_0_13_LC_14_10_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_fast_esr_RNIFGGE_0_13_LC_14_10_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_fast_esr_RNIFGGE_0_13_LC_14_10_4 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_d_reg_fast_esr_RNIFGGE_0_13_LC_14_10_4  (
            .in0(N__90911),
            .in1(N__82324),
            .in2(_gnd_net_),
            .in3(N__79121),
            .lcout(\pid_side.error_d_reg_fast_esr_RNIFGGE_0Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI5RIO_0_14_LC_14_10_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI5RIO_0_14_LC_14_10_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI5RIO_0_14_LC_14_10_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI5RIO_0_14_LC_14_10_5  (
            .in0(N__79168),
            .in1(N__90847),
            .in2(_gnd_net_),
            .in3(N__91431),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI5RIO_0Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI5RIO_14_LC_14_10_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI5RIO_14_LC_14_10_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI5RIO_14_LC_14_10_6 .LUT_INIT=16'b1010000011111010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI5RIO_14_LC_14_10_6  (
            .in0(N__91432),
            .in1(_gnd_net_),
            .in2(N__90855),
            .in3(N__79169),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI5RIOZ0Z_14 ),
            .ltout(\pid_side.error_d_reg_prev_esr_RNI5RIOZ0Z_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI73UC2_0_14_LC_14_10_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI73UC2_0_14_LC_14_10_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI73UC2_0_14_LC_14_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI73UC2_0_14_LC_14_10_7  (
            .in0(_gnd_net_),
            .in1(N__67810),
            .in2(N__59932),
            .in3(N__62480),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI73UC2_0Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIS8JL1_0_21_LC_14_11_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIS8JL1_0_21_LC_14_11_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIS8JL1_0_21_LC_14_11_0 .LUT_INIT=16'b0001100011100111;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIS8JL1_0_21_LC_14_11_0  (
            .in0(N__91642),
            .in1(N__91329),
            .in2(N__72950),
            .in3(N__62916),
            .lcout(\pid_side.un1_pid_prereg_0_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIQ5IL1_21_LC_14_11_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIQ5IL1_21_LC_14_11_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIQ5IL1_21_LC_14_11_1 .LUT_INIT=16'b1110111100001000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIQ5IL1_21_LC_14_11_1  (
            .in0(N__91328),
            .in1(N__91643),
            .in2(N__72948),
            .in3(N__72659),
            .lcout(\pid_side.un1_pid_prereg_0_20 ),
            .ltout(\pid_side.un1_pid_prereg_0_20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI8N8M6_21_LC_14_11_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI8N8M6_21_LC_14_11_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI8N8M6_21_LC_14_11_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI8N8M6_21_LC_14_11_2  (
            .in0(N__72640),
            .in1(N__68443),
            .in2(N__60484),
            .in3(N__60468),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI8N8M6Z0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIS8JL1_21_LC_14_11_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIS8JL1_21_LC_14_11_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIS8JL1_21_LC_14_11_3 .LUT_INIT=16'b1011101010100010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIS8JL1_21_LC_14_11_3  (
            .in0(N__62915),
            .in1(N__72940),
            .in2(N__91357),
            .in3(N__91645),
            .lcout(\pid_side.un1_pid_prereg_0_22 ),
            .ltout(\pid_side.un1_pid_prereg_0_22_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIG3DM6_21_LC_14_11_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIG3DM6_21_LC_14_11_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIG3DM6_21_LC_14_11_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIG3DM6_21_LC_14_11_4  (
            .in0(N__60469),
            .in1(N__60478),
            .in2(N__60481),
            .in3(N__68318),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIG3DM6Z0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIUBKL1_0_21_LC_14_11_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIUBKL1_0_21_LC_14_11_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIUBKL1_0_21_LC_14_11_5 .LUT_INIT=16'b0001100011100111;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIUBKL1_0_21_LC_14_11_5  (
            .in0(N__91330),
            .in1(N__91644),
            .in2(N__72949),
            .in3(N__67880),
            .lcout(\pid_side.un1_pid_prereg_0_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIME5B3_21_LC_14_11_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIME5B3_21_LC_14_11_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIME5B3_21_LC_14_11_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIME5B3_21_LC_14_11_6  (
            .in0(_gnd_net_),
            .in1(N__60477),
            .in2(_gnd_net_),
            .in3(N__60467),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIME5B3Z0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIQK7B3_21_LC_14_11_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIQK7B3_21_LC_14_11_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIQK7B3_21_LC_14_11_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIQK7B3_21_LC_14_11_7  (
            .in0(N__68319),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68340),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIQK7B3Z0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNISPAE1_0_13_LC_14_12_0 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNISPAE1_0_13_LC_14_12_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNISPAE1_0_13_LC_14_12_0 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNISPAE1_0_13_LC_14_12_0  (
            .in0(N__60585),
            .in1(N__60594),
            .in2(N__60576),
            .in3(N__60618),
            .lcout(\pid_side.error_i_acumm_13_i_o2_0_10_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_13_LC_14_12_1 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_13_LC_14_12_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_13_LC_14_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_13_LC_14_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76511),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94144),
            .ce(N__65078),
            .sr(N__86439));
    defparam \pid_side.error_i_acumm_prereg_esr_RNISPAE1_13_LC_14_12_2 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNISPAE1_13_LC_14_12_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNISPAE1_13_LC_14_12_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNISPAE1_13_LC_14_12_2  (
            .in0(N__60586),
            .in1(N__60595),
            .in2(N__60577),
            .in3(N__60619),
            .lcout(\pid_side.error_i_acumm_13_i_o2_0_10_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_18_LC_14_12_3 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_18_LC_14_12_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_18_LC_14_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_18_LC_14_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65236),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94144),
            .ce(N__65078),
            .sr(N__86439));
    defparam \pid_side.error_i_acumm_prereg_esr_25_LC_14_12_4 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_25_LC_14_12_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_25_LC_14_12_4 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_25_LC_14_12_4  (
            .in0(_gnd_net_),
            .in1(N__72660),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94144),
            .ce(N__65078),
            .sr(N__86439));
    defparam \pid_side.error_i_acumm_prereg_esr_26_LC_14_12_5 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_26_LC_14_12_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_26_LC_14_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_26_LC_14_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62917),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94144),
            .ce(N__65078),
            .sr(N__86439));
    defparam \pid_side.error_d_reg_prev_esr_RNI9LLC4_12_LC_14_12_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI9LLC4_12_LC_14_12_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI9LLC4_12_LC_14_12_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI9LLC4_12_LC_14_12_6  (
            .in0(N__76510),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68542),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI9LLC4Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_27_LC_14_12_7 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_27_LC_14_12_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_27_LC_14_12_7 .LUT_INIT=16'b1100110011001110;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_27_LC_14_12_7  (
            .in0(N__81333),
            .in1(N__60562),
            .in2(N__84837),
            .in3(N__85939),
            .lcout(\pid_side.N_42_i_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_1_sqmuxa_1_i_a2_0_4_LC_14_13_0 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_1_sqmuxa_1_i_a2_0_4_LC_14_13_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_1_sqmuxa_1_i_a2_0_4_LC_14_13_0 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \pid_side.error_i_acumm_1_sqmuxa_1_i_a2_0_4_LC_14_13_0  (
            .in0(N__73367),
            .in1(N__68713),
            .in2(N__69190),
            .in3(N__84433),
            .lcout(pid_side_N_382_4),
            .ltout(pid_side_N_382_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.state_RNIU7A12_0_LC_14_13_1 .C_ON=1'b0;
    defparam \pid_side.state_RNIU7A12_0_LC_14_13_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.state_RNIU7A12_0_LC_14_13_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \pid_side.state_RNIU7A12_0_LC_14_13_1  (
            .in0(N__60789),
            .in1(N__70066),
            .in2(N__60556),
            .in3(N__70022),
            .lcout(),
            .ltout(\pid_side.N_382_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.state_RNIC78N2_0_LC_14_13_2 .C_ON=1'b0;
    defparam \pid_side.state_RNIC78N2_0_LC_14_13_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.state_RNIC78N2_0_LC_14_13_2 .LUT_INIT=16'b1111101011111110;
    LogicCell40 \pid_side.state_RNIC78N2_0_LC_14_13_2  (
            .in0(N__70851),
            .in1(N__60698),
            .in2(N__60553),
            .in3(N__60790),
            .lcout(\pid_side.N_64 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.state_RNIQ7UK_0_LC_14_13_3 .C_ON=1'b0;
    defparam \pid_side.state_RNIQ7UK_0_LC_14_13_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.state_RNIQ7UK_0_LC_14_13_3 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \pid_side.state_RNIQ7UK_0_LC_14_13_3  (
            .in0(N__69178),
            .in1(N__60691),
            .in2(_gnd_net_),
            .in3(N__60784),
            .lcout(\pid_side.state_ns_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.state_0_LC_14_13_4 .C_ON=1'b0;
    defparam \pid_side.state_0_LC_14_13_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.state_0_LC_14_13_4 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \pid_side.state_0_LC_14_13_4  (
            .in0(N__69177),
            .in1(N__60699),
            .in2(_gnd_net_),
            .in3(N__60791),
            .lcout(\pid_side.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94156),
            .ce(),
            .sr(N__86435));
    defparam \pid_side.state_RNIL5IF_0_LC_14_13_5 .C_ON=1'b0;
    defparam \pid_side.state_RNIL5IF_0_LC_14_13_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.state_RNIL5IF_0_LC_14_13_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pid_side.state_RNIL5IF_0_LC_14_13_5  (
            .in0(_gnd_net_),
            .in1(N__60783),
            .in2(_gnd_net_),
            .in3(N__70850),
            .lcout(\pid_side.state_RNIL5IFZ0Z_0 ),
            .ltout(\pid_side.state_RNIL5IFZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.state_RNIIIOO_0_LC_14_13_6 .C_ON=1'b0;
    defparam \pid_side.state_RNIIIOO_0_LC_14_13_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.state_RNIIIOO_0_LC_14_13_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_side.state_RNIIIOO_0_LC_14_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__60835),
            .in3(N__93121),
            .lcout(\pid_side.state_RNIIIOOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.state_1_LC_14_13_7 .C_ON=1'b0;
    defparam \pid_side.state_1_LC_14_13_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.state_1_LC_14_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.state_1_LC_14_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60785),
            .lcout(\pid_side.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94156),
            .ce(),
            .sr(N__86435));
    defparam \pid_front.state_RNI26LH_0_LC_14_14_1 .C_ON=1'b0;
    defparam \pid_front.state_RNI26LH_0_LC_14_14_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.state_RNI26LH_0_LC_14_14_1 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \pid_front.state_RNI26LH_0_LC_14_14_1  (
            .in0(N__70605),
            .in1(N__69182),
            .in2(_gnd_net_),
            .in3(N__70515),
            .lcout(\pid_front.state_ns_0 ),
            .ltout(\pid_front.state_ns_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.state_RNI9MMH_0_LC_14_14_2 .C_ON=1'b0;
    defparam \pid_front.state_RNI9MMH_0_LC_14_14_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.state_RNI9MMH_0_LC_14_14_2 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \pid_front.state_RNI9MMH_0_LC_14_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__60655),
            .in3(N__86587),
            .lcout(\pid_front.state_ns_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.m9_2_03_3_i_0_a2_1_0_LC_14_14_5 .C_ON=1'b0;
    defparam \pid_front.m9_2_03_3_i_0_a2_1_0_LC_14_14_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.m9_2_03_3_i_0_a2_1_0_LC_14_14_5 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \pid_front.m9_2_03_3_i_0_a2_1_0_LC_14_14_5  (
            .in0(N__90404),
            .in1(N__90156),
            .in2(N__90645),
            .in3(N__83002),
            .lcout(\pid_front.N_536_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_0_22_LC_14_14_7 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_22_LC_14_14_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_22_LC_14_14_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_22_LC_14_14_7  (
            .in0(N__81419),
            .in1(N__60640),
            .in2(_gnd_net_),
            .in3(N__80696),
            .lcout(\pid_front.N_301 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_18_LC_14_15_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_18_LC_14_15_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_18_LC_14_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_18_LC_14_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60634),
            .lcout(\pid_front.error_p_regZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94182),
            .ce(N__93258),
            .sr(N__92982));
    defparam \pid_front.error_p_reg_esr_RNIUAE8_4_LC_14_15_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIUAE8_4_LC_14_15_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIUAE8_4_LC_14_15_3 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_front.error_p_reg_esr_RNIUAE8_4_LC_14_15_3  (
            .in0(N__61152),
            .in1(N__66961),
            .in2(_gnd_net_),
            .in3(N__66977),
            .lcout(\pid_front.error_p_reg_esr_RNIUAE8Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_4_LC_14_15_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_4_LC_14_15_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_4_LC_14_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_4_LC_14_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60895),
            .lcout(\pid_front.error_p_regZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94182),
            .ce(N__93258),
            .sr(N__92982));
    defparam \pid_front.error_d_reg_esr_4_LC_14_15_5 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_4_LC_14_15_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_4_LC_14_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_4_LC_14_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60874),
            .lcout(\pid_front.error_d_regZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94182),
            .ce(N__93258),
            .sr(N__92982));
    defparam \pid_side.error_axb_8_l_ofx_LC_14_15_6 .C_ON=1'b0;
    defparam \pid_side.error_axb_8_l_ofx_LC_14_15_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_axb_8_l_ofx_LC_14_15_6 .LUT_INIT=16'b1111010111110101;
    LogicCell40 \pid_side.error_axb_8_l_ofx_LC_14_15_6  (
            .in0(N__60862),
            .in1(_gnd_net_),
            .in2(N__85279),
            .in3(N__77481),
            .lcout(\pid_side.error_axb_8_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_axb_7_LC_14_15_7 .C_ON=1'b0;
    defparam \pid_side.error_axb_7_LC_14_15_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_axb_7_LC_14_15_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_side.error_axb_7_LC_14_15_7  (
            .in0(_gnd_net_),
            .in1(N__85275),
            .in2(_gnd_net_),
            .in3(N__60861),
            .lcout(\pid_side.error_axbZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_0_c_RNIJB0R2_LC_14_16_0 .C_ON=1'b0;
    defparam \pid_front.error_cry_0_0_c_RNIJB0R2_LC_14_16_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_0_c_RNIJB0R2_LC_14_16_0 .LUT_INIT=16'b0010101000100000;
    LogicCell40 \pid_front.error_cry_0_0_c_RNIJB0R2_LC_14_16_0  (
            .in0(N__76866),
            .in1(N__74221),
            .in2(N__89374),
            .in3(N__77084),
            .lcout(\pid_front.N_581 ),
            .ltout(\pid_front.N_581_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_0_10_LC_14_16_1 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_10_LC_14_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_10_LC_14_16_1 .LUT_INIT=16'b1111110011110000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_10_LC_14_16_1  (
            .in0(_gnd_net_),
            .in1(N__81311),
            .in2(N__60847),
            .in3(N__60931),
            .lcout(),
            .ltout(\pid_front.error_i_reg_esr_RNO_0Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_10_LC_14_16_2 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_10_LC_14_16_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_10_LC_14_16_2 .LUT_INIT=16'b1100110011000000;
    LogicCell40 \pid_front.error_i_reg_esr_10_LC_14_16_2  (
            .in0(_gnd_net_),
            .in1(N__83378),
            .in2(N__60844),
            .in3(N__60975),
            .lcout(\pid_front.error_i_regZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94194),
            .ce(N__78105),
            .sr(N__86405));
    defparam \pid_front.error_i_reg_esr_26_LC_14_16_3 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_26_LC_14_16_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_26_LC_14_16_3 .LUT_INIT=16'b1110111011110000;
    LogicCell40 \pid_front.error_i_reg_esr_26_LC_14_16_3  (
            .in0(N__60976),
            .in1(N__60841),
            .in2(N__65995),
            .in3(N__60922),
            .lcout(\pid_front.error_i_regZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94194),
            .ce(N__78105),
            .sr(N__86405));
    defparam \pid_front.error_cry_1_0_c_RNII2EF1_0_LC_14_16_4 .C_ON=1'b0;
    defparam \pid_front.error_cry_1_0_c_RNII2EF1_0_LC_14_16_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_1_0_c_RNII2EF1_0_LC_14_16_4 .LUT_INIT=16'b0010001100100000;
    LogicCell40 \pid_front.error_cry_1_0_c_RNII2EF1_0_LC_14_16_4  (
            .in0(N__77855),
            .in1(N__89590),
            .in2(N__90254),
            .in3(N__78305),
            .lcout(),
            .ltout(\pid_front.error_cry_1_0_c_RNII2EF1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_1_0_c_RNIM2834_LC_14_16_5 .C_ON=1'b0;
    defparam \pid_front.error_cry_1_0_c_RNIM2834_LC_14_16_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_1_0_c_RNIM2834_LC_14_16_5 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \pid_front.error_cry_1_0_c_RNIM2834_LC_14_16_5  (
            .in0(_gnd_net_),
            .in1(N__61018),
            .in2(N__60934),
            .in3(N__60916),
            .lcout(\pid_front.N_228 ),
            .ltout(\pid_front.N_228_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_1_26_LC_14_16_6 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_1_26_LC_14_16_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_1_26_LC_14_16_6 .LUT_INIT=16'b0100110000000000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_1_26_LC_14_16_6  (
            .in0(N__81310),
            .in1(N__87098),
            .in2(N__60925),
            .in3(N__84522),
            .lcout(\pid_front.error_i_reg_9_sn_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_1_0_c_RNII2EF1_LC_14_16_7 .C_ON=1'b0;
    defparam \pid_front.error_cry_1_0_c_RNII2EF1_LC_14_16_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_1_0_c_RNII2EF1_LC_14_16_7 .LUT_INIT=16'b1111111011110010;
    LogicCell40 \pid_front.error_cry_1_0_c_RNII2EF1_LC_14_16_7  (
            .in0(N__78304),
            .in1(N__90240),
            .in2(N__89602),
            .in3(N__77854),
            .lcout(\pid_front.error_cry_1_0_c_RNII2EFZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_2_0_c_RNIANSH2_LC_14_17_0 .C_ON=1'b0;
    defparam \pid_front.error_cry_2_0_c_RNIANSH2_LC_14_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_2_0_c_RNIANSH2_LC_14_17_0 .LUT_INIT=16'b0101110100001000;
    LogicCell40 \pid_front.error_cry_2_0_c_RNIANSH2_LC_14_17_0  (
            .in0(N__82764),
            .in1(N__77732),
            .in2(N__85178),
            .in3(N__66209),
            .lcout(\pid_front.N_182 ),
            .ltout(\pid_front.N_182_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_6_c_RNI3O1T5_0_LC_14_17_1 .C_ON=1'b0;
    defparam \pid_front.error_cry_6_c_RNI3O1T5_0_LC_14_17_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_6_c_RNI3O1T5_0_LC_14_17_1 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \pid_front.error_cry_6_c_RNI3O1T5_0_LC_14_17_1  (
            .in0(N__89604),
            .in1(N__89078),
            .in2(N__60910),
            .in3(N__69702),
            .lcout(\pid_front.N_597 ),
            .ltout(\pid_front.N_597_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_0_24_LC_14_17_2 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_24_LC_14_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_24_LC_14_17_2 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_24_LC_14_17_2  (
            .in0(N__85764),
            .in1(N__63160),
            .in2(N__60907),
            .in3(N__60901),
            .lcout(),
            .ltout(\pid_front.m12_2_03_4_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_24_LC_14_17_3 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_24_LC_14_17_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_24_LC_14_17_3 .LUT_INIT=16'b1010000000100010;
    LogicCell40 \pid_front.error_i_reg_esr_24_LC_14_17_3  (
            .in0(N__87048),
            .in1(N__60967),
            .in2(N__60904),
            .in3(N__84521),
            .lcout(\pid_front.error_i_regZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94211),
            .ce(N__78146),
            .sr(N__86396));
    defparam \pid_front.error_cry_0_c_RNIT6SM2_LC_14_17_4 .C_ON=1'b0;
    defparam \pid_front.error_cry_0_c_RNIT6SM2_LC_14_17_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_c_RNIT6SM2_LC_14_17_4 .LUT_INIT=16'b0000111100001000;
    LogicCell40 \pid_front.error_cry_0_c_RNIT6SM2_LC_14_17_4  (
            .in0(N__74176),
            .in1(N__74966),
            .in2(N__87802),
            .in3(N__66073),
            .lcout(\pid_front.N_583 ),
            .ltout(\pid_front.N_583_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_0_8_LC_14_17_5 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_8_LC_14_17_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_8_LC_14_17_5 .LUT_INIT=16'b1111110011110000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_8_LC_14_17_5  (
            .in0(_gnd_net_),
            .in1(N__85763),
            .in2(N__60988),
            .in3(N__63154),
            .lcout(),
            .ltout(\pid_front.error_i_reg_esr_RNO_0Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_8_LC_14_17_6 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_8_LC_14_17_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_8_LC_14_17_6 .LUT_INIT=16'b1111110000000000;
    LogicCell40 \pid_front.error_i_reg_esr_8_LC_14_17_6  (
            .in0(_gnd_net_),
            .in1(N__60985),
            .in2(N__60979),
            .in3(N__83379),
            .lcout(\pid_front.error_i_regZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94211),
            .ce(N__78146),
            .sr(N__86396));
    defparam \pid_front.error_cry_6_c_RNI3O1T5_LC_14_17_7 .C_ON=1'b0;
    defparam \pid_front.error_cry_6_c_RNI3O1T5_LC_14_17_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_6_c_RNI3O1T5_LC_14_17_7 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \pid_front.error_cry_6_c_RNI3O1T5_LC_14_17_7  (
            .in0(N__89603),
            .in1(N__69703),
            .in2(N__73633),
            .in3(N__89079),
            .lcout(\pid_front.N_598 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_1_24_LC_14_18_0 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_1_24_LC_14_18_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_1_24_LC_14_18_0 .LUT_INIT=16'b1100110011101111;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_1_24_LC_14_18_0  (
            .in0(N__81443),
            .in1(N__60961),
            .in2(N__87448),
            .in3(N__80670),
            .lcout(\pid_front.m28_2_03_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_2_24_LC_14_18_1 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_2_24_LC_14_18_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_2_24_LC_14_18_1 .LUT_INIT=16'b0000001110101011;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_2_24_LC_14_18_1  (
            .in0(N__76954),
            .in1(N__73897),
            .in2(N__73383),
            .in3(N__78311),
            .lcout(\pid_front.m28_2_03_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_2_25_LC_14_18_2 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_2_25_LC_14_18_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_2_25_LC_14_18_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_2_25_LC_14_18_2  (
            .in0(N__78312),
            .in1(N__73379),
            .in2(_gnd_net_),
            .in3(N__80669),
            .lcout(),
            .ltout(\pid_front.N_302_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_0_25_LC_14_18_3 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_25_LC_14_18_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_25_LC_14_18_3 .LUT_INIT=16'b1010101010100000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_25_LC_14_18_3  (
            .in0(N__86991),
            .in1(_gnd_net_),
            .in2(N__60955),
            .in3(N__84516),
            .lcout(),
            .ltout(\pid_front.error_i_reg_9_rn_2_25_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_25_LC_14_18_4 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_25_LC_14_18_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_25_LC_14_18_4 .LUT_INIT=16'b1110111011110000;
    LogicCell40 \pid_front.error_i_reg_esr_25_LC_14_18_4  (
            .in0(N__63067),
            .in1(N__63268),
            .in2(N__60952),
            .in3(N__60949),
            .lcout(\pid_front.error_i_regZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94227),
            .ce(N__78148),
            .sr(N__86386));
    defparam \pid_front.error_i_reg_esr_RNO_1_25_LC_14_18_5 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_1_25_LC_14_18_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_1_25_LC_14_18_5 .LUT_INIT=16'b0000100010001000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_1_25_LC_14_18_5  (
            .in0(N__86990),
            .in1(N__84515),
            .in2(N__69504),
            .in3(N__74721),
            .lcout(\pid_front.error_i_reg_9_sn_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_21_LC_14_18_6 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_21_LC_14_18_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_21_LC_14_18_6 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \pid_front.error_i_reg_esr_21_LC_14_18_6  (
            .in0(N__84517),
            .in1(N__60994),
            .in2(N__60943),
            .in3(N__86992),
            .lcout(\pid_front.error_i_regZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94227),
            .ce(N__78148),
            .sr(N__86386));
    defparam \pid_front.error_i_reg_esr_23_LC_14_18_7 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_23_LC_14_18_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_23_LC_14_18_7 .LUT_INIT=16'b1011000000010000;
    LogicCell40 \pid_front.error_i_reg_esr_23_LC_14_18_7  (
            .in0(N__84563),
            .in1(N__61030),
            .in2(N__87055),
            .in3(N__63226),
            .lcout(\pid_front.error_i_regZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94227),
            .ce(N__78148),
            .sr(N__86386));
    defparam \pid_front.error_cry_1_0_c_RNIPIJ12_LC_14_19_0 .C_ON=1'b0;
    defparam \pid_front.error_cry_1_0_c_RNIPIJ12_LC_14_19_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_1_0_c_RNIPIJ12_LC_14_19_0 .LUT_INIT=16'b0100111001000100;
    LogicCell40 \pid_front.error_cry_1_0_c_RNIPIJ12_LC_14_19_0  (
            .in0(N__89591),
            .in1(N__61014),
            .in2(N__89375),
            .in3(N__77849),
            .lcout(\pid_front.N_207 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_5_c_RNIITB41_LC_14_19_1 .C_ON=1'b0;
    defparam \pid_front.error_cry_5_c_RNIITB41_LC_14_19_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_5_c_RNIITB41_LC_14_19_1 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \pid_front.error_cry_5_c_RNIITB41_LC_14_19_1  (
            .in0(N__80002),
            .in1(N__78376),
            .in2(N__90256),
            .in3(_gnd_net_),
            .lcout(\pid_front.N_154 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_5_c_RNILLSA1_LC_14_19_2 .C_ON=1'b0;
    defparam \pid_front.error_cry_5_c_RNILLSA1_LC_14_19_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_5_c_RNILLSA1_LC_14_19_2 .LUT_INIT=16'b0001110100000000;
    LogicCell40 \pid_front.error_cry_5_c_RNILLSA1_LC_14_19_2  (
            .in0(N__78275),
            .in1(N__90432),
            .in2(N__78395),
            .in3(N__90251),
            .lcout(\pid_front.N_225 ),
            .ltout(\pid_front.N_225_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_0_19_LC_14_19_3 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_19_LC_14_19_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_19_LC_14_19_3 .LUT_INIT=16'b0011111100010101;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_19_LC_14_19_3  (
            .in0(N__88888),
            .in1(N__76875),
            .in2(N__61003),
            .in3(N__74473),
            .lcout(\pid_front.error_i_reg_esr_RNO_0Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_1_0_c_RNIDC571_LC_14_19_4 .C_ON=1'b0;
    defparam \pid_front.error_cry_1_0_c_RNIDC571_LC_14_19_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_1_0_c_RNIDC571_LC_14_19_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \pid_front.error_cry_1_0_c_RNIDC571_LC_14_19_4  (
            .in0(N__78274),
            .in1(N__90247),
            .in2(_gnd_net_),
            .in3(N__77848),
            .lcout(\pid_front.N_188 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_3_21_LC_14_19_5 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_3_21_LC_14_19_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_3_21_LC_14_19_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_3_21_LC_14_19_5  (
            .in0(N__73860),
            .in1(N__62947),
            .in2(_gnd_net_),
            .in3(N__62932),
            .lcout(),
            .ltout(\pid_front.N_478_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_1_21_LC_14_19_6 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_1_21_LC_14_19_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_1_21_LC_14_19_6 .LUT_INIT=16'b0000111100001101;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_1_21_LC_14_19_6  (
            .in0(N__76876),
            .in1(N__81441),
            .in2(N__61000),
            .in3(N__74270),
            .lcout(),
            .ltout(\pid_front.error_i_reg_9_N_5L8_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_0_21_LC_14_19_7 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_21_LC_14_19_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_21_LC_14_19_7 .LUT_INIT=16'b0000000010110000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_21_LC_14_19_7  (
            .in0(N__87790),
            .in1(N__66332),
            .in2(N__60997),
            .in3(N__80527),
            .lcout(\pid_front.error_i_reg_esr_RNO_0Z0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_0_c_RNI85F82_LC_14_20_0 .C_ON=1'b0;
    defparam \pid_front.error_cry_0_0_c_RNI85F82_LC_14_20_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_0_c_RNI85F82_LC_14_20_0 .LUT_INIT=16'b0000001011110010;
    LogicCell40 \pid_front.error_cry_0_0_c_RNI85F82_LC_14_20_0  (
            .in0(N__83029),
            .in1(N__77959),
            .in2(N__90676),
            .in3(N__63177),
            .lcout(),
            .ltout(\pid_front.N_45_i_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_1_0_c_RNINF5A3_LC_14_20_1 .C_ON=1'b0;
    defparam \pid_front.error_cry_1_0_c_RNINF5A3_LC_14_20_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_1_0_c_RNINF5A3_LC_14_20_1 .LUT_INIT=16'b0000111100000011;
    LogicCell40 \pid_front.error_cry_1_0_c_RNINF5A3_LC_14_20_1  (
            .in0(_gnd_net_),
            .in1(N__81322),
            .in2(N__61132),
            .in3(N__77856),
            .lcout(\pid_front.error_cry_1_0_c_RNINF5AZ0Z3 ),
            .ltout(\pid_front.error_cry_1_0_c_RNINF5AZ0Z3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_1_18_LC_14_20_2 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_1_18_LC_14_20_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_1_18_LC_14_20_2 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_1_18_LC_14_20_2  (
            .in0(_gnd_net_),
            .in1(N__84192),
            .in2(N__61129),
            .in3(N__66264),
            .lcout(\pid_front.m6_2_01 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_4_18_LC_14_20_3 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_4_18_LC_14_20_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_4_18_LC_14_20_3 .LUT_INIT=16'b0010000000101111;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_4_18_LC_14_20_3  (
            .in0(N__76877),
            .in1(N__77089),
            .in2(N__89376),
            .in3(N__80677),
            .lcout(),
            .ltout(\pid_front.un4_error_i_reg_28_ns_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_2_18_LC_14_20_4 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_2_18_LC_14_20_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_2_18_LC_14_20_4 .LUT_INIT=16'b0000000000000111;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_2_18_LC_14_20_4  (
            .in0(N__81323),
            .in1(N__66333),
            .in2(N__61126),
            .in3(N__74530),
            .lcout(),
            .ltout(\pid_front.un4_error_i_reg_28_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_18_LC_14_20_5 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_18_LC_14_20_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_18_LC_14_20_5 .LUT_INIT=16'b1001100000010000;
    LogicCell40 \pid_front.error_i_reg_esr_18_LC_14_20_5  (
            .in0(N__84550),
            .in1(N__61123),
            .in2(N__61111),
            .in3(N__61108),
            .lcout(\pid_front.error_i_regZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94262),
            .ce(N__78135),
            .sr(N__86373));
    defparam \pid_front.error_d_reg_prev_esr_RNIIUAC3_20_LC_14_21_0 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIIUAC3_20_LC_14_21_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIIUAC3_20_LC_14_21_0 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIIUAC3_20_LC_14_21_0  (
            .in0(N__64174),
            .in1(N__66622),
            .in2(_gnd_net_),
            .in3(N__71390),
            .lcout(\pid_front.un1_pid_prereg_0_12 ),
            .ltout(\pid_front.un1_pid_prereg_0_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIV42AC_21_LC_14_21_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIV42AC_21_LC_14_21_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIV42AC_21_LC_14_21_1 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIV42AC_21_LC_14_21_1  (
            .in0(N__61102),
            .in1(N__61214),
            .in2(N__61078),
            .in3(N__61075),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIV42ACZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIU58I5_21_LC_14_21_2 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIU58I5_21_LC_14_21_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIU58I5_21_LC_14_21_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIU58I5_21_LC_14_21_2  (
            .in0(N__61215),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61242),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIU58I5Z0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIC7T52_21_LC_14_21_3 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIC7T52_21_LC_14_21_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIC7T52_21_LC_14_21_3 .LUT_INIT=16'b1110111100001000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIC7T52_21_LC_14_21_3  (
            .in0(N__91718),
            .in1(N__66708),
            .in2(N__67093),
            .in3(N__69909),
            .lcout(\pid_front.un1_pid_prereg_0_14 ),
            .ltout(\pid_front.un1_pid_prereg_0_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNION3U9_21_LC_14_21_4 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNION3U9_21_LC_14_21_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNION3U9_21_LC_14_21_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNION3U9_21_LC_14_21_4  (
            .in0(N__61216),
            .in1(N__61243),
            .in2(N__61234),
            .in3(N__61557),
            .lcout(\pid_front.error_d_reg_prev_esr_RNION3U9Z0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIC7T52_0_21_LC_14_21_5 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIC7T52_0_21_LC_14_21_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIC7T52_0_21_LC_14_21_5 .LUT_INIT=16'b0001100011100111;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIC7T52_0_21_LC_14_21_5  (
            .in0(N__91717),
            .in1(N__66707),
            .in2(N__67092),
            .in3(N__69908),
            .lcout(\pid_front.un1_pid_prereg_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIEAU52_0_21_LC_14_21_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIEAU52_0_21_LC_14_21_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIEAU52_0_21_LC_14_21_6 .LUT_INIT=16'b0001111010000111;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIEAU52_0_21_LC_14_21_6  (
            .in0(N__66709),
            .in1(N__91719),
            .in2(N__72131),
            .in3(N__67078),
            .lcout(\pid_front.un1_pid_prereg_0_15 ),
            .ltout(\pid_front.un1_pid_prereg_0_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIQHRB4_21_LC_14_21_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIQHRB4_21_LC_14_21_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIQHRB4_21_LC_14_21_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIQHRB4_21_LC_14_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__61204),
            .in3(N__61578),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIQHRB4Z0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNID8DF2_3_LC_14_22_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNID8DF2_3_LC_14_22_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNID8DF2_3_LC_14_22_0 .LUT_INIT=16'b1110100011101000;
    LogicCell40 \pid_front.error_p_reg_esr_RNID8DF2_3_LC_14_22_0  (
            .in0(N__75510),
            .in1(N__61141),
            .in2(N__61177),
            .in3(N__61632),
            .lcout(\pid_front.error_p_reg_esr_RNID8DF2Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIR7E8_3_LC_14_22_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIR7E8_3_LC_14_22_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIR7E8_3_LC_14_22_1 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \pid_front.error_p_reg_esr_RNIR7E8_3_LC_14_22_1  (
            .in0(N__78768),
            .in1(_gnd_net_),
            .in2(N__61408),
            .in3(N__61429),
            .lcout(\pid_front.error_p_reg_esr_RNIR7E8Z0Z_3 ),
            .ltout(\pid_front.error_p_reg_esr_RNIR7E8Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIRJAF2_3_LC_14_22_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIRJAF2_3_LC_14_22_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIRJAF2_3_LC_14_22_2 .LUT_INIT=16'b1001011010010110;
    LogicCell40 \pid_front.error_p_reg_esr_RNIRJAF2_3_LC_14_22_2  (
            .in0(N__75509),
            .in1(N__61140),
            .in2(N__61168),
            .in3(N__61443),
            .lcout(\pid_front.error_p_reg_esr_RNIRJAF2Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIUAE8_0_4_LC_14_22_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIUAE8_0_4_LC_14_22_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIUAE8_0_4_LC_14_22_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_p_reg_esr_RNIUAE8_0_4_LC_14_22_3  (
            .in0(N__61159),
            .in1(N__66960),
            .in2(_gnd_net_),
            .in3(N__66990),
            .lcout(\pid_front.error_p_reg_esr_RNIUAE8_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_3_LC_14_22_4 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_3_LC_14_22_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_3_LC_14_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_3_LC_14_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78769),
            .lcout(\pid_front.error_d_reg_prevZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94296),
            .ce(N__71747),
            .sr(N__71628));
    defparam \pid_front.error_p_reg_esr_RNIPKK71_2_LC_14_22_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIPKK71_2_LC_14_22_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIPKK71_2_LC_14_22_5 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIPKK71_2_LC_14_22_5  (
            .in0(N__61396),
            .in1(N__63574),
            .in2(_gnd_net_),
            .in3(N__74589),
            .lcout(\pid_front.error_p_reg_esr_RNIPKK71Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIR7E8_0_3_LC_14_22_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIR7E8_0_3_LC_14_22_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIR7E8_0_3_LC_14_22_6 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_p_reg_esr_RNIR7E8_0_3_LC_14_22_6  (
            .in0(N__61428),
            .in1(N__61404),
            .in2(_gnd_net_),
            .in3(N__78767),
            .lcout(\pid_front.error_p_reg_esr_RNIR7E8_0Z0Z_3 ),
            .ltout(\pid_front.error_p_reg_esr_RNIR7E8_0Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIQ7CF2_2_LC_14_22_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIQ7CF2_2_LC_14_22_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIQ7CF2_2_LC_14_22_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_p_reg_esr_RNIQ7CF2_2_LC_14_22_7  (
            .in0(N__61291),
            .in1(N__63573),
            .in2(N__61390),
            .in3(N__74588),
            .lcout(\pid_front.error_p_reg_esr_RNIQ7CF2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNI1JN71_1_LC_14_23_0 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNI1JN71_1_LC_14_23_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNI1JN71_1_LC_14_23_0 .LUT_INIT=16'b1111110111010000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNI1JN71_1_LC_14_23_0  (
            .in0(N__61378),
            .in1(N__61345),
            .in2(N__63615),
            .in3(N__61312),
            .lcout(\pid_front.error_d_reg_prev_esr_RNI1JN71Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.state_RNIR49E_0_LC_14_23_1 .C_ON=1'b0;
    defparam \pid_alt.state_RNIR49E_0_LC_14_23_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.state_RNIR49E_0_LC_14_23_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pid_alt.state_RNIR49E_0_LC_14_23_1  (
            .in0(_gnd_net_),
            .in1(N__69077),
            .in2(_gnd_net_),
            .in3(N__86580),
            .lcout(\pid_alt.state_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNI1K4E5_0_10_LC_14_23_2 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNI1K4E5_0_10_LC_14_23_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNI1K4E5_0_10_LC_14_23_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNI1K4E5_0_10_LC_14_23_2  (
            .in0(N__75136),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63761),
            .lcout(\pid_front.error_d_reg_prev_esr_RNI1K4E5_0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNI1K4E5_10_LC_14_23_3 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNI1K4E5_10_LC_14_23_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNI1K4E5_10_LC_14_23_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNI1K4E5_10_LC_14_23_3  (
            .in0(N__63762),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75137),
            .lcout(\pid_front.error_d_reg_prev_esr_RNI1K4E5Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNI80O6_8_LC_14_23_4 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNI80O6_8_LC_14_23_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNI80O6_8_LC_14_23_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNI80O6_8_LC_14_23_4  (
            .in0(_gnd_net_),
            .in1(N__71338),
            .in2(_gnd_net_),
            .in3(N__78805),
            .lcout(\pid_front.N_2370_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIUO6U_1_12_LC_14_23_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIUO6U_1_12_LC_14_23_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIUO6U_1_12_LC_14_23_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIUO6U_1_12_LC_14_23_6  (
            .in0(_gnd_net_),
            .in1(N__78703),
            .in2(_gnd_net_),
            .in3(N__81833),
            .lcout(\pid_front.g1_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIB9N71_5_LC_14_23_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIB9N71_5_LC_14_23_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIB9N71_5_LC_14_23_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIB9N71_5_LC_14_23_7  (
            .in0(_gnd_net_),
            .in1(N__61651),
            .in2(_gnd_net_),
            .in3(N__75282),
            .lcout(\pid_front.error_p_reg_esr_RNIB9N71Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIJS6B3_0_15_LC_14_24_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIJS6B3_0_15_LC_14_24_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIJS6B3_0_15_LC_14_24_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_p_reg_esr_RNIJS6B3_0_15_LC_14_24_0  (
            .in0(N__63789),
            .in1(N__67134),
            .in2(_gnd_net_),
            .in3(N__71255),
            .lcout(\pid_front.un1_pid_prereg_0_1 ),
            .ltout(\pid_front.un1_pid_prereg_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIUFCM6_14_LC_14_24_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIUFCM6_14_LC_14_24_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIUFCM6_14_LC_14_24_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIUFCM6_14_LC_14_24_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__61498),
            .in3(N__61476),
            .lcout(\pid_front.error_p_reg_esr_RNIUFCM6Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIJS6B3_15_LC_14_24_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIJS6B3_15_LC_14_24_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIJS6B3_15_LC_14_24_2 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIJS6B3_15_LC_14_24_2  (
            .in0(N__63790),
            .in1(N__67135),
            .in2(_gnd_net_),
            .in3(N__71256),
            .lcout(\pid_front.un1_pid_prereg_0_2 ),
            .ltout(\pid_front.un1_pid_prereg_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNICIRCD_14_LC_14_24_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNICIRCD_14_LC_14_24_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNICIRCD_14_LC_14_24_3 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_front.error_p_reg_esr_RNICIRCD_14_LC_14_24_3  (
            .in0(N__61468),
            .in1(N__61477),
            .in2(N__61486),
            .in3(N__63836),
            .lcout(\pid_front.error_p_reg_esr_RNICIRCDZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIR58B3_0_16_LC_14_24_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIR58B3_0_16_LC_14_24_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIR58B3_0_16_LC_14_24_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_p_reg_esr_RNIR58B3_0_16_LC_14_24_4  (
            .in0(N__63870),
            .in1(N__63882),
            .in2(_gnd_net_),
            .in3(N__71219),
            .lcout(\pid_front.un1_pid_prereg_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIBJ5B3_14_LC_14_24_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIBJ5B3_14_LC_14_24_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIBJ5B3_14_LC_14_24_5 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIBJ5B3_14_LC_14_24_5  (
            .in0(N__71116),
            .in1(N__71146),
            .in2(_gnd_net_),
            .in3(N__71131),
            .lcout(\pid_front.un1_pid_prereg_0_0 ),
            .ltout(\pid_front.un1_pid_prereg_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIA6C3N_14_LC_14_24_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIA6C3N_14_LC_14_24_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIA6C3N_14_LC_14_24_6 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pid_front.error_p_reg_esr_RNIA6C3N_14_LC_14_24_6  (
            .in0(N__71092),
            .in1(N__61467),
            .in2(N__61459),
            .in3(N__71562),
            .lcout(\pid_front.error_p_reg_esr_RNIA6C3NZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIQ9AED_10_LC_14_24_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIQ9AED_10_LC_14_24_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIQ9AED_10_LC_14_24_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIQ9AED_10_LC_14_24_7  (
            .in0(N__63763),
            .in1(N__63718),
            .in2(N__75151),
            .in3(N__63742),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIQ9AEDZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIGDV52_0_21_LC_14_25_0 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIGDV52_0_21_LC_14_25_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIGDV52_0_21_LC_14_25_0 .LUT_INIT=16'b0001100011100111;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIGDV52_0_21_LC_14_25_0  (
            .in0(N__91758),
            .in1(N__66704),
            .in2(N__67097),
            .in3(N__71183),
            .lcout(\pid_front.un1_pid_prereg_0_17 ),
            .ltout(\pid_front.un1_pid_prereg_0_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIUNTB4_21_LC_14_25_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIUNTB4_21_LC_14_25_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIUNTB4_21_LC_14_25_1 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIUNTB4_21_LC_14_25_1  (
            .in0(N__63735),
            .in1(_gnd_net_),
            .in2(N__61606),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIUNTB4Z0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIGDV52_21_LC_14_25_2 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIGDV52_21_LC_14_25_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIGDV52_21_LC_14_25_2 .LUT_INIT=16'b1110111100001000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIGDV52_21_LC_14_25_2  (
            .in0(N__91759),
            .in1(N__66705),
            .in2(N__67098),
            .in3(N__71184),
            .lcout(\pid_front.un1_pid_prereg_0_18 ),
            .ltout(\pid_front.un1_pid_prereg_0_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNI0MTN8_21_LC_14_25_3 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNI0MTN8_21_LC_14_25_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNI0MTN8_21_LC_14_25_3 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNI0MTN8_21_LC_14_25_3  (
            .in0(N__63736),
            .in1(N__61546),
            .in2(N__61594),
            .in3(N__61836),
            .lcout(\pid_front.error_d_reg_prev_esr_RNI0MTN8Z0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIO9PN8_21_LC_14_25_4 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIO9PN8_21_LC_14_25_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIO9PN8_21_LC_14_25_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIO9PN8_21_LC_14_25_4  (
            .in0(N__61585),
            .in1(N__63734),
            .in2(N__61567),
            .in3(N__61545),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIO9PN8Z0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIE2FM6_15_LC_14_25_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIE2FM6_15_LC_14_25_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIE2FM6_15_LC_14_25_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIE2FM6_15_LC_14_25_5  (
            .in0(_gnd_net_),
            .in1(N__63849),
            .in2(_gnd_net_),
            .in3(N__63837),
            .lcout(\pid_front.error_p_reg_esr_RNIE2FM6Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIIG062_0_21_LC_14_25_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIIG062_0_21_LC_14_25_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIIG062_0_21_LC_14_25_6 .LUT_INIT=16'b0110010101011001;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIIG062_0_21_LC_14_25_6  (
            .in0(N__64086),
            .in1(N__67088),
            .in2(N__91773),
            .in3(N__66706),
            .lcout(\pid_front.un1_pid_prereg_0_19 ),
            .ltout(\pid_front.un1_pid_prereg_0_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNI2UVB4_21_LC_14_25_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNI2UVB4_21_LC_14_25_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNI2UVB4_21_LC_14_25_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNI2UVB4_21_LC_14_25_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__61519),
            .in3(N__61854),
            .lcout(\pid_front.error_d_reg_prev_esr_RNI2UVB4Z0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIMVC9_0_6_LC_14_26_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIMVC9_0_6_LC_14_26_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIMVC9_0_6_LC_14_26_0 .LUT_INIT=16'b0011100111000110;
    LogicCell40 \pid_front.error_p_reg_esr_RNIMVC9_0_6_LC_14_26_0  (
            .in0(N__61704),
            .in1(N__81725),
            .in2(N__94681),
            .in3(N__61783),
            .lcout(\pid_front.error_p_reg_esr_RNIMVC9_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_5_LC_14_26_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_5_LC_14_26_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_5_LC_14_26_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_5_LC_14_26_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__94678),
            .lcout(\pid_front.error_d_reg_prevZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94356),
            .ce(N__71809),
            .sr(N__71705));
    defparam \pid_front.error_p_reg_esr_RNIJ26O1_5_LC_14_26_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIJ26O1_5_LC_14_26_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIJ26O1_5_LC_14_26_2 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIJ26O1_5_LC_14_26_2  (
            .in0(N__75226),
            .in1(_gnd_net_),
            .in2(N__61741),
            .in3(N__61717),
            .lcout(\pid_front.error_p_reg_esr_RNIJ26O1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIK9971_6_LC_14_26_3 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIK9971_6_LC_14_26_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIK9971_6_LC_14_26_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIK9971_6_LC_14_26_3  (
            .in0(_gnd_net_),
            .in1(N__61737),
            .in2(_gnd_net_),
            .in3(N__75225),
            .lcout(),
            .ltout(\pid_front.un1_pid_prereg_66_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIUBTV2_5_LC_14_26_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIUBTV2_5_LC_14_26_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIUBTV2_5_LC_14_26_4 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pid_front.error_p_reg_esr_RNIUBTV2_5_LC_14_26_4  (
            .in0(N__75281),
            .in1(N__61716),
            .in2(N__61729),
            .in3(N__61650),
            .lcout(\pid_front.error_p_reg_esr_RNIUBTV2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIVOSG_5_LC_14_26_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIVOSG_5_LC_14_26_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIVOSG_5_LC_14_26_5 .LUT_INIT=16'b1101010011101000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIVOSG_5_LC_14_26_5  (
            .in0(N__94680),
            .in1(N__61668),
            .in2(N__61684),
            .in3(N__61706),
            .lcout(\pid_front.error_p_reg_esr_RNIVOSGZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIVOSG_0_5_LC_14_26_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIVOSG_0_5_LC_14_26_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIVOSG_0_5_LC_14_26_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \pid_front.error_p_reg_esr_RNIVOSG_0_5_LC_14_26_6  (
            .in0(N__61705),
            .in1(N__61680),
            .in2(N__61669),
            .in3(N__94679),
            .lcout(\pid_front.error_p_reg_esr_RNIVOSG_0Z0Z_5 ),
            .ltout(\pid_front.error_p_reg_esr_RNIVOSG_0Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIB9N71_0_5_LC_14_26_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIB9N71_0_5_LC_14_26_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIB9N71_0_5_LC_14_26_7 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIB9N71_0_5_LC_14_26_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__61636),
            .in3(N__75280),
            .lcout(\pid_front.error_p_reg_esr_RNIB9N71_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIIG062_21_LC_14_27_0 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIIG062_21_LC_14_27_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIIG062_21_LC_14_27_0 .LUT_INIT=16'b1010100011101010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIIG062_21_LC_14_27_0  (
            .in0(N__64085),
            .in1(N__66668),
            .in2(N__91780),
            .in3(N__67091),
            .lcout(\pid_front.un1_pid_prereg_0_20 ),
            .ltout(\pid_front.un1_pid_prereg_0_20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNI642C4_21_LC_14_27_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNI642C4_21_LC_14_27_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNI642C4_21_LC_14_27_1 .LUT_INIT=16'b1100000011000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNI642C4_21_LC_14_27_1  (
            .in0(_gnd_net_),
            .in1(N__61794),
            .in2(N__61882),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prev_esr_RNI642C4Z0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_esr_RNIETB61_3_13_LC_14_27_2 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_RNIETB61_3_13_LC_14_27_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_esr_RNIETB61_3_13_LC_14_27_2 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_d_reg_esr_RNIETB61_3_13_LC_14_27_2  (
            .in0(N__64352),
            .in1(N__67687),
            .in2(_gnd_net_),
            .in3(N__67639),
            .lcout(\pid_front.error_d_reg_esr_RNIETB61_3Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIKJ162_21_LC_14_27_3 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIKJ162_21_LC_14_27_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIKJ162_21_LC_14_27_3 .LUT_INIT=16'b1111110101000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIKJ162_21_LC_14_27_3  (
            .in0(N__67089),
            .in1(N__91779),
            .in2(N__66691),
            .in3(N__64053),
            .lcout(\pid_front.un1_pid_prereg_0_22 ),
            .ltout(\pid_front.un1_pid_prereg_0_22_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIGE6O8_21_LC_14_27_4 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIGE6O8_21_LC_14_27_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIGE6O8_21_LC_14_27_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIGE6O8_21_LC_14_27_4  (
            .in0(N__61795),
            .in1(N__61825),
            .in2(N__61870),
            .in3(N__66777),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIGE6O8Z0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNI822O8_21_LC_14_27_5 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNI822O8_21_LC_14_27_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNI822O8_21_LC_14_27_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNI822O8_21_LC_14_27_5  (
            .in0(N__61861),
            .in1(N__61793),
            .in2(N__61843),
            .in3(N__61824),
            .lcout(\pid_front.error_d_reg_prev_esr_RNI822O8Z0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIMM262_0_21_LC_14_27_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIMM262_0_21_LC_14_27_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIMM262_0_21_LC_14_27_6 .LUT_INIT=16'b0001111010000111;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIMM262_0_21_LC_14_27_6  (
            .in0(N__91775),
            .in1(N__66667),
            .in2(N__69883),
            .in3(N__67090),
            .lcout(\pid_front.un1_pid_prereg_0_23 ),
            .ltout(\pid_front.un1_pid_prereg_0_23_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIAA4C4_21_LC_14_27_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIAA4C4_21_LC_14_27_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIAA4C4_21_LC_14_27_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIAA4C4_21_LC_14_27_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__61807),
            .in3(N__66756),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIAA4C4Z0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIKJ162_0_21_LC_14_28_0 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIKJ162_0_21_LC_14_28_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIKJ162_0_21_LC_14_28_0 .LUT_INIT=16'b0001100011100111;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIKJ162_0_21_LC_14_28_0  (
            .in0(N__91774),
            .in1(N__66663),
            .in2(N__67099),
            .in3(N__64052),
            .lcout(\pid_front.un1_pid_prereg_0_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_esr_RNIETB61_2_13_LC_14_28_3 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_RNIETB61_2_13_LC_14_28_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_esr_RNIETB61_2_13_LC_14_28_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_d_reg_esr_RNIETB61_2_13_LC_14_28_3  (
            .in0(N__64353),
            .in1(N__67686),
            .in2(_gnd_net_),
            .in3(N__67641),
            .lcout(\pid_front.N_4_1_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_14_LC_15_3_0 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_14_LC_15_3_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_14_LC_15_3_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_14_LC_15_3_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76551),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94088),
            .ce(N__65070),
            .sr(N__86475));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIQGO21_0_14_LC_15_3_1 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIQGO21_0_14_LC_15_3_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIQGO21_0_14_LC_15_3_1 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIQGO21_0_14_LC_15_3_1  (
            .in0(N__61917),
            .in1(N__61932),
            .in2(_gnd_net_),
            .in3(N__62013),
            .lcout(\pid_side.error_i_acumm_13_i_o2_0_7_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIKIBE1_0_19_LC_15_3_2 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIKIBE1_0_19_LC_15_3_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIKIBE1_0_19_LC_15_3_2 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIKIBE1_0_19_LC_15_3_2  (
            .in0(N__62181),
            .in1(N__61893),
            .in2(N__62169),
            .in3(N__62193),
            .lcout(\pid_side.error_i_acumm_13_i_o2_0_8_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIRN9E1_0_15_LC_15_3_3 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIRN9E1_0_15_LC_15_3_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIRN9E1_0_15_LC_15_3_3 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIRN9E1_0_15_LC_15_3_3  (
            .in0(N__62119),
            .in1(N__62151),
            .in2(N__62677),
            .in3(N__62107),
            .lcout(),
            .ltout(\pid_side.error_i_acumm_13_i_o2_0_9_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNI5LOD5_13_LC_15_3_4 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNI5LOD5_13_LC_15_3_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNI5LOD5_13_LC_15_3_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNI5LOD5_13_LC_15_3_4  (
            .in0(N__62002),
            .in1(N__61987),
            .in2(N__61981),
            .in3(N__61978),
            .lcout(\pid_side.N_203 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_22_LC_15_3_6 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_22_LC_15_3_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_22_LC_15_3_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_22_LC_15_3_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67990),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94088),
            .ce(N__65070),
            .sr(N__86475));
    defparam \pid_side.error_i_acumm_prereg_esr_27_LC_15_3_7 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_27_LC_15_3_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_27_LC_15_3_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_27_LC_15_3_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67890),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94088),
            .ce(N__65070),
            .sr(N__86475));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIKIBE1_19_LC_15_4_0 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIKIBE1_19_LC_15_4_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIKIBE1_19_LC_15_4_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIKIBE1_19_LC_15_4_0  (
            .in0(N__62182),
            .in1(N__61894),
            .in2(N__62170),
            .in3(N__62194),
            .lcout(\pid_side.error_i_acumm_13_i_o2_0_8_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_19_LC_15_4_1 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_19_LC_15_4_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_19_LC_15_4_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_19_LC_15_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65407),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94094),
            .ce(N__65071),
            .sr(N__86466));
    defparam \pid_side.error_i_acumm_prereg_esr_20_LC_15_4_2 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_20_LC_15_4_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_20_LC_15_4_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_20_LC_15_4_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65278),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94094),
            .ce(N__65071),
            .sr(N__86466));
    defparam \pid_side.error_i_acumm_prereg_esr_21_LC_15_4_3 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_21_LC_15_4_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_21_LC_15_4_3 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_21_LC_15_4_3  (
            .in0(_gnd_net_),
            .in1(N__65308),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94094),
            .ce(N__65071),
            .sr(N__86466));
    defparam \pid_side.error_i_acumm_prereg_esr_23_LC_15_4_4 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_23_LC_15_4_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_23_LC_15_4_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_23_LC_15_4_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68254),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94094),
            .ce(N__65071),
            .sr(N__86466));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIRN9E1_15_LC_15_4_5 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIRN9E1_15_LC_15_4_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIRN9E1_15_LC_15_4_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIRN9E1_15_LC_15_4_5  (
            .in0(N__62152),
            .in1(N__62106),
            .in2(N__62676),
            .in3(N__62118),
            .lcout(\pid_side.error_i_acumm_13_i_o2_0_9_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_15_LC_15_4_6 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_15_LC_15_4_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_15_LC_15_4_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_15_LC_15_4_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62491),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94094),
            .ce(N__65071),
            .sr(N__86466));
    defparam \pid_side.error_i_acumm_prereg_esr_16_LC_15_4_7 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_16_LC_15_4_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_16_LC_15_4_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_16_LC_15_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62632),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94094),
            .ce(N__65071),
            .sr(N__86466));
    defparam \pid_side.pid_prereg_esr_RNI2L63_24_LC_15_5_0 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNI2L63_24_LC_15_5_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNI2L63_24_LC_15_5_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_side.pid_prereg_esr_RNI2L63_24_LC_15_5_0  (
            .in0(N__64906),
            .in1(N__64930),
            .in2(N__65197),
            .in3(N__64942),
            .lcout(\pid_side.un11lto30_i_a2_5_and ),
            .ltout(\pid_side.un11lto30_i_a2_5_and_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNI5HTB_16_LC_15_5_1 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNI5HTB_16_LC_15_5_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNI5HTB_16_LC_15_5_1 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \pid_side.pid_prereg_esr_RNI5HTB_16_LC_15_5_1  (
            .in0(N__62244),
            .in1(N__62217),
            .in2(N__62086),
            .in3(N__62232),
            .lcout(\pid_side.N_175 ),
            .ltout(\pid_side.N_175_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNI9ACR_15_LC_15_5_2 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNI9ACR_15_LC_15_5_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNI9ACR_15_LC_15_5_2 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \pid_side.pid_prereg_esr_RNI9ACR_15_LC_15_5_2  (
            .in0(_gnd_net_),
            .in1(N__64743),
            .in2(N__62068),
            .in3(N__62064),
            .lcout(\pid_side.N_277 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNIB2E2_28_LC_15_5_3 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNIB2E2_28_LC_15_5_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNIB2E2_28_LC_15_5_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \pid_side.pid_prereg_esr_RNIB2E2_28_LC_15_5_3  (
            .in0(N__65164),
            .in1(N__65108),
            .in2(_gnd_net_),
            .in3(N__65152),
            .lcout(\pid_side.un11lto30_i_a2_6_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNI6L23_16_LC_15_5_4 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNI6L23_16_LC_15_5_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNI6L23_16_LC_15_5_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_side.pid_prereg_esr_RNI6L23_16_LC_15_5_4  (
            .in0(N__64693),
            .in1(N__64669),
            .in2(N__64996),
            .in3(N__64717),
            .lcout(\pid_side.un11lto30_i_a2_3_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNII463_20_LC_15_5_5 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNII463_20_LC_15_5_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNII463_20_LC_15_5_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_side.pid_prereg_esr_RNII463_20_LC_15_5_5  (
            .in0(N__64975),
            .in1(N__64966),
            .in2(N__64957),
            .in3(N__64984),
            .lcout(\pid_side.un11lto30_i_a2_4_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIFCVC2_0_15_LC_15_6_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIFCVC2_0_15_LC_15_6_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIFCVC2_0_15_LC_15_6_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIFCVC2_0_15_LC_15_6_0  (
            .in0(N__62271),
            .in1(N__67782),
            .in2(_gnd_net_),
            .in3(N__62630),
            .lcout(\pid_side.un1_pid_prereg_0_1 ),
            .ltout(\pid_side.un1_pid_prereg_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIMFTP4_14_LC_15_6_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIMFTP4_14_LC_15_6_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIMFTP4_14_LC_15_6_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIMFTP4_14_LC_15_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__62203),
            .in3(N__62343),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIMFTP4Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIFCVC2_15_LC_15_6_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIFCVC2_15_LC_15_6_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIFCVC2_15_LC_15_6_2 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIFCVC2_15_LC_15_6_2  (
            .in0(N__62272),
            .in1(N__67783),
            .in2(_gnd_net_),
            .in3(N__62631),
            .lcout(\pid_side.un1_pid_prereg_0_2 ),
            .ltout(\pid_side.un1_pid_prereg_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNISHTJ9_14_LC_15_6_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNISHTJ9_14_LC_15_6_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNISHTJ9_14_LC_15_6_3 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNISHTJ9_14_LC_15_6_3  (
            .in0(N__62344),
            .in1(N__62329),
            .in2(N__62200),
            .in3(N__62295),
            .lcout(\pid_side.error_d_reg_prev_esr_RNISHTJ9Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNINL0D2_0_16_LC_15_6_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNINL0D2_0_16_LC_15_6_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNINL0D2_0_16_LC_15_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNINL0D2_0_16_LC_15_6_4  (
            .in0(N__62259),
            .in1(N__62320),
            .in2(_gnd_net_),
            .in3(N__62606),
            .lcout(\pid_side.un1_pid_prereg_0_3 ),
            .ltout(\pid_side.un1_pid_prereg_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI620Q4_15_LC_15_6_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI620Q4_15_LC_15_6_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI620Q4_15_LC_15_6_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI620Q4_15_LC_15_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__62197),
            .in3(N__62307),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI620Q4Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI73UC2_14_LC_15_6_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI73UC2_14_LC_15_6_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI73UC2_14_LC_15_6_6 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI73UC2_14_LC_15_6_6  (
            .in0(N__62356),
            .in1(N__67809),
            .in2(_gnd_net_),
            .in3(N__62487),
            .lcout(\pid_side.un1_pid_prereg_0_0 ),
            .ltout(\pid_side.un1_pid_prereg_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI2SL2G_12_LC_15_6_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI2SL2G_12_LC_15_6_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI2SL2G_12_LC_15_6_7 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI2SL2G_12_LC_15_6_7  (
            .in0(N__68040),
            .in1(N__68593),
            .in2(N__62332),
            .in3(N__62328),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI2SL2GZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIB1JO_16_LC_15_7_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIB1JO_16_LC_15_7_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIB1JO_16_LC_15_7_0 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIB1JO_16_LC_15_7_0  (
            .in0(N__90046),
            .in1(N__62281),
            .in2(_gnd_net_),
            .in3(N__92709),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIB1JOZ0Z_16 ),
            .ltout(\pid_side.error_d_reg_prev_esr_RNIB1JOZ0Z_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNINL0D2_16_LC_15_7_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNINL0D2_16_LC_15_7_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNINL0D2_16_LC_15_7_1 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNINL0D2_16_LC_15_7_1  (
            .in0(_gnd_net_),
            .in1(N__62260),
            .in2(N__62311),
            .in3(N__62607),
            .lcout(\pid_side.un1_pid_prereg_0_4 ),
            .ltout(\pid_side.un1_pid_prereg_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNISM2K9_15_LC_15_7_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNISM2K9_15_LC_15_7_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNISM2K9_15_LC_15_7_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNISM2K9_15_LC_15_7_2  (
            .in0(N__62308),
            .in1(N__62296),
            .in2(N__62284),
            .in3(N__68196),
            .lcout(\pid_side.error_d_reg_prev_esr_RNISM2K9Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_16_LC_15_7_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_16_LC_15_7_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_16_LC_15_7_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_16_LC_15_7_3  (
            .in0(N__92710),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94112),
            .ce(N__88090),
            .sr(N__87941));
    defparam \pid_side.error_d_reg_prev_esr_RNIB1JO_0_16_LC_15_7_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIB1JO_0_16_LC_15_7_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIB1JO_0_16_LC_15_7_4 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIB1JO_0_16_LC_15_7_4  (
            .in0(N__90045),
            .in1(N__62280),
            .in2(_gnd_net_),
            .in3(N__92708),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIB1JO_0Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIE4JO_0_17_LC_15_7_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIE4JO_0_17_LC_15_7_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIE4JO_0_17_LC_15_7_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIE4JO_0_17_LC_15_7_5  (
            .in0(N__90789),
            .in1(N__67753),
            .in2(_gnd_net_),
            .in3(N__91174),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIE4JO_0Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIVU1D2_0_17_LC_15_7_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIVU1D2_0_17_LC_15_7_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIVU1D2_0_17_LC_15_7_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIVU1D2_0_17_LC_15_7_6  (
            .in0(N__87853),
            .in1(N__67771),
            .in2(_gnd_net_),
            .in3(N__65235),
            .lcout(\pid_side.un1_pid_prereg_0_5 ),
            .ltout(\pid_side.un1_pid_prereg_0_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIMK2Q4_16_LC_15_7_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIMK2Q4_16_LC_15_7_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIMK2Q4_16_LC_15_7_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIMK2Q4_16_LC_15_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__62464),
            .in3(N__68217),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIMK2Q4Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_RNI115E_0_LC_15_8_0 .C_ON=1'b1;
    defparam \pid_side.error_i_acumm_RNI115E_0_LC_15_8_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_RNI115E_0_LC_15_8_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pid_side.error_i_acumm_RNI115E_0_LC_15_8_0  (
            .in0(_gnd_net_),
            .in1(N__62451),
            .in2(N__63015),
            .in3(_gnd_net_),
            .lcout(\pid_side.un1_pid_prereg_0 ),
            .ltout(),
            .carryin(bfn_15_8_0_),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_0_c_RNITGKN_LC_15_8_1 .C_ON=1'b1;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_0_c_RNITGKN_LC_15_8_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_0_c_RNITGKN_LC_15_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_0_c_RNITGKN_LC_15_8_1  (
            .in0(_gnd_net_),
            .in1(N__62440),
            .in2(N__62653),
            .in3(N__62434),
            .lcout(\pid_side.un1_error_i_acumm_prereg_cry_0_c_RNITGKN ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_0 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_1_c_RNI0LLN_LC_15_8_2 .C_ON=1'b1;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_1_c_RNI0LLN_LC_15_8_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_1_c_RNI0LLN_LC_15_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_1_c_RNI0LLN_LC_15_8_2  (
            .in0(_gnd_net_),
            .in1(N__62431),
            .in2(N__79504),
            .in3(N__62425),
            .lcout(\pid_side.un1_error_i_acumm_prereg_cry_1_c_RNI0LLN ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_1 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_2_c_RNIQUGJ_LC_15_8_3 .C_ON=1'b1;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_2_c_RNIQUGJ_LC_15_8_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_2_c_RNIQUGJ_LC_15_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_2_c_RNIQUGJ_LC_15_8_3  (
            .in0(_gnd_net_),
            .in1(N__62421),
            .in2(N__62401),
            .in3(N__62389),
            .lcout(\pid_side.un1_error_i_acumm_prereg_cry_2_c_RNIQUGJ ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_2 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_3_c_RNI6TNN_LC_15_8_4 .C_ON=1'b1;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_3_c_RNI6TNN_LC_15_8_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_3_c_RNI6TNN_LC_15_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_3_c_RNI6TNN_LC_15_8_4  (
            .in0(_gnd_net_),
            .in1(N__62386),
            .in2(N__83203),
            .in3(N__62377),
            .lcout(\pid_side.un1_error_i_acumm_prereg_cry_3_c_RNI6TNN ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_3 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_4_c_RNI91PN_LC_15_8_5 .C_ON=1'b1;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_4_c_RNI91PN_LC_15_8_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_4_c_RNI91PN_LC_15_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_4_c_RNI91PN_LC_15_8_5  (
            .in0(_gnd_net_),
            .in1(N__62374),
            .in2(N__79681),
            .in3(N__62368),
            .lcout(\pid_side.un1_error_i_acumm_prereg_cry_4_c_RNI91PN ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_4 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_5_c_RNIC5QN_LC_15_8_6 .C_ON=1'b1;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_5_c_RNIC5QN_LC_15_8_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_5_c_RNIC5QN_LC_15_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_5_c_RNIC5QN_LC_15_8_6  (
            .in0(_gnd_net_),
            .in1(N__62365),
            .in2(N__68815),
            .in3(N__62359),
            .lcout(\pid_side.un1_error_i_acumm_prereg_cry_5_c_RNIC5QN ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_5 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_6_c_RNI6FLJ_LC_15_8_7 .C_ON=1'b1;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_6_c_RNI6FLJ_LC_15_8_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_6_c_RNI6FLJ_LC_15_8_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_6_c_RNI6FLJ_LC_15_8_7  (
            .in0(_gnd_net_),
            .in1(N__65442),
            .in2(N__62560),
            .in3(N__62551),
            .lcout(\pid_side.un1_error_i_acumm_prereg_cry_6_c_RNI6FLJ ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_6 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_7_c_RNIIDSN_LC_15_9_0 .C_ON=1'b1;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_7_c_RNIIDSN_LC_15_9_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_7_c_RNIIDSN_LC_15_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_7_c_RNIIDSN_LC_15_9_0  (
            .in0(_gnd_net_),
            .in1(N__62548),
            .in2(N__72151),
            .in3(N__62539),
            .lcout(\pid_side.un1_error_i_acumm_prereg_cry_7_c_RNIIDSN ),
            .ltout(),
            .carryin(bfn_15_9_0_),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_8_c_RNICNNJ_LC_15_9_1 .C_ON=1'b1;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_8_c_RNICNNJ_LC_15_9_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_8_c_RNICNNJ_LC_15_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_8_c_RNICNNJ_LC_15_9_1  (
            .in0(_gnd_net_),
            .in1(N__62536),
            .in2(N__65503),
            .in3(N__62527),
            .lcout(\pid_side.un1_error_i_acumm_prereg_cry_8_c_RNICNNJ ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_8 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNI6OOI_10_LC_15_9_2 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNI6OOI_10_LC_15_9_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNI6OOI_10_LC_15_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNI6OOI_10_LC_15_9_2  (
            .in0(_gnd_net_),
            .in1(N__62524),
            .in2(N__73528),
            .in3(N__62518),
            .lcout(\pid_side.error_i_reg_esr_RNI6OOIZ0Z_10 ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_9 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNIGRJR_11_LC_15_9_3 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNIGRJR_11_LC_15_9_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNIGRJR_11_LC_15_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNIGRJR_11_LC_15_9_3  (
            .in0(_gnd_net_),
            .in1(N__62515),
            .in2(N__68788),
            .in3(N__62509),
            .lcout(\pid_side.error_i_reg_esr_RNIGRJRZ0Z_11 ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_10 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNIJVKR_12_LC_15_9_4 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNIJVKR_12_LC_15_9_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNIJVKR_12_LC_15_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNIJVKR_12_LC_15_9_4  (
            .in0(_gnd_net_),
            .in1(N__62506),
            .in2(N__68851),
            .in3(N__62500),
            .lcout(\pid_side.error_i_reg_esr_RNIJVKRZ0Z_12 ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_11 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNIM3MR_13_LC_15_9_5 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNIM3MR_13_LC_15_9_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNIM3MR_13_LC_15_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNIM3MR_13_LC_15_9_5  (
            .in0(_gnd_net_),
            .in1(N__62876),
            .in2(N__68728),
            .in3(N__62497),
            .lcout(\pid_side.error_i_reg_esr_RNIM3MRZ0Z_13 ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_12 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNIO6NR_14_LC_15_9_6 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNIO6NR_14_LC_15_9_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNIO6NR_14_LC_15_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNIO6NR_14_LC_15_9_6  (
            .in0(_gnd_net_),
            .in1(N__62956),
            .in2(N__62894),
            .in3(N__62494),
            .lcout(\pid_side.error_i_reg_esr_RNIO6NRZ0Z_14 ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_13 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNIQ9OR_15_LC_15_9_7 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNIQ9OR_15_LC_15_9_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNIQ9OR_15_LC_15_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNIQ9OR_15_LC_15_9_7  (
            .in0(_gnd_net_),
            .in1(N__62880),
            .in2(N__76588),
            .in3(N__62467),
            .lcout(\pid_side.error_i_reg_esr_RNIQ9ORZ0Z_15 ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_14 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNISCPR_16_LC_15_10_0 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNISCPR_16_LC_15_10_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNISCPR_16_LC_15_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNISCPR_16_LC_15_10_0  (
            .in0(_gnd_net_),
            .in1(N__62849),
            .in2(N__66118),
            .in3(N__62614),
            .lcout(\pid_side.error_i_reg_esr_RNISCPRZ0Z_16 ),
            .ltout(),
            .carryin(bfn_15_10_0_),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNIUFQR_17_LC_15_10_1 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNIUFQR_17_LC_15_10_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNIUFQR_17_LC_15_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNIUFQR_17_LC_15_10_1  (
            .in0(_gnd_net_),
            .in1(N__68872),
            .in2(N__62881),
            .in3(N__62584),
            .lcout(\pid_side.error_i_reg_esr_RNIUFQRZ0Z_17 ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_16 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNI0JRR_18_LC_15_10_2 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNI0JRR_18_LC_15_10_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNI0JRR_18_LC_15_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNI0JRR_18_LC_15_10_2  (
            .in0(_gnd_net_),
            .in1(N__62853),
            .in2(N__79552),
            .in3(N__62581),
            .lcout(\pid_side.error_i_reg_esr_RNI0JRRZ0Z_18 ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_17 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNI2MSR_19_LC_15_10_3 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNI2MSR_19_LC_15_10_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNI2MSR_19_LC_15_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNI2MSR_19_LC_15_10_3  (
            .in0(_gnd_net_),
            .in1(N__86797),
            .in2(N__62882),
            .in3(N__62578),
            .lcout(\pid_side.error_i_reg_esr_RNI2MSRZ0Z_19 ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_18 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNIRGUR_20_LC_15_10_4 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNIRGUR_20_LC_15_10_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNIRGUR_20_LC_15_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNIRGUR_20_LC_15_10_4  (
            .in0(_gnd_net_),
            .in1(N__62857),
            .in2(N__83698),
            .in3(N__62575),
            .lcout(\pid_side.error_i_reg_esr_RNIRGURZ0Z_20 ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_19 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNIK2OS_21_LC_15_10_5 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNIK2OS_21_LC_15_10_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNIK2OS_21_LC_15_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNIK2OS_21_LC_15_10_5  (
            .in0(_gnd_net_),
            .in1(N__81355),
            .in2(N__62883),
            .in3(N__62572),
            .lcout(\pid_side.error_i_reg_esr_RNIK2OSZ0Z_21 ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_20 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNIM5PS_22_LC_15_10_6 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNIM5PS_22_LC_15_10_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNIM5PS_22_LC_15_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNIM5PS_22_LC_15_10_6  (
            .in0(_gnd_net_),
            .in1(N__62861),
            .in2(N__73501),
            .in3(N__62569),
            .lcout(\pid_side.error_i_reg_esr_RNIM5PSZ0Z_22 ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_21 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNIO8QS_23_LC_15_10_7 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNIO8QS_23_LC_15_10_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNIO8QS_23_LC_15_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNIO8QS_23_LC_15_10_7  (
            .in0(_gnd_net_),
            .in1(N__73252),
            .in2(N__62884),
            .in3(N__62566),
            .lcout(\pid_side.error_i_reg_esr_RNIO8QSZ0Z_23 ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_22 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNIQBRS_24_LC_15_11_0 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNIQBRS_24_LC_15_11_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNIQBRS_24_LC_15_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNIQBRS_24_LC_15_11_0  (
            .in0(_gnd_net_),
            .in1(N__62885),
            .in2(N__73333),
            .in3(N__62563),
            .lcout(\pid_side.error_i_reg_esr_RNIQBRSZ0Z_24 ),
            .ltout(),
            .carryin(bfn_15_11_0_),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNISESS_25_LC_15_11_1 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNISESS_25_LC_15_11_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNISESS_25_LC_15_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNISESS_25_LC_15_11_1  (
            .in0(_gnd_net_),
            .in1(N__62638),
            .in2(N__62895),
            .in3(N__62920),
            .lcout(\pid_side.error_i_reg_esr_RNISESSZ0Z_25 ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_24 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNIUHTS_26_LC_15_11_2 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNIUHTS_26_LC_15_11_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNIUHTS_26_LC_15_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNIUHTS_26_LC_15_11_2  (
            .in0(_gnd_net_),
            .in1(N__62889),
            .in2(N__73567),
            .in3(N__62902),
            .lcout(\pid_side.error_i_reg_esr_RNIUHTSZ0Z_26 ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_25 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_26_c_RNI0LUS_LC_15_11_3 .C_ON=1'b1;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_26_c_RNI0LUS_LC_15_11_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_26_c_RNI0LUS_LC_15_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_26_c_RNI0LUS_LC_15_11_3  (
            .in0(_gnd_net_),
            .in1(N__62964),
            .in2(N__62896),
            .in3(N__62899),
            .lcout(\pid_side.un1_error_i_acumm_prereg_cry_26_c_RNI0LUS ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_26 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_27_c_RNI1NVS_LC_15_11_4 .C_ON=1'b0;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_27_c_RNI1NVS_LC_15_11_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_27_c_RNI1NVS_LC_15_11_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_27_c_RNI1NVS_LC_15_11_4  (
            .in0(N__62965),
            .in1(N__62893),
            .in2(_gnd_net_),
            .in3(N__62800),
            .lcout(\pid_side.un1_error_i_acumm_prereg_cry_27_c_RNI1NVS ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_28_LC_15_11_5 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_28_LC_15_11_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_28_LC_15_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_28_LC_15_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72603),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94145),
            .ce(N__65079),
            .sr(N__86440));
    defparam \pid_side.error_i_acumm_prereg_esr_24_LC_15_11_6 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_24_LC_15_11_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_24_LC_15_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_24_LC_15_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68169),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94145),
            .ce(N__65079),
            .sr(N__86440));
    defparam \pid_side.error_i_reg_esr_1_LC_15_12_0 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_1_LC_15_12_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_1_LC_15_12_0 .LUT_INIT=16'b1100010000000100;
    LogicCell40 \pid_side.error_i_reg_esr_1_LC_15_12_0  (
            .in0(N__66133),
            .in1(N__82082),
            .in2(N__84118),
            .in3(N__77622),
            .lcout(\pid_side.error_i_regZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94157),
            .ce(N__86744),
            .sr(N__86436));
    defparam \pid_side.error_i_reg_esr_RNO_0_25_LC_15_12_1 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_25_LC_15_12_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_25_LC_15_12_1 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_25_LC_15_12_1  (
            .in0(N__81653),
            .in1(_gnd_net_),
            .in2(N__73387),
            .in3(N__85934),
            .lcout(),
            .ltout(\pid_side.N_302_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_25_LC_15_12_2 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_25_LC_15_12_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_25_LC_15_12_2 .LUT_INIT=16'b1000100011000000;
    LogicCell40 \pid_side.error_i_reg_esr_25_LC_15_12_2  (
            .in0(N__65512),
            .in1(N__87034),
            .in2(N__62641),
            .in3(N__84575),
            .lcout(\pid_side.error_i_regZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94157),
            .ce(N__86744),
            .sr(N__86436));
    defparam \pid_side.m78_0_a2_0_0_LC_15_12_3 .C_ON=1'b0;
    defparam \pid_side.m78_0_a2_0_0_LC_15_12_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.m78_0_a2_0_0_LC_15_12_3 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \pid_side.m78_0_a2_0_0_LC_15_12_3  (
            .in0(N__87032),
            .in1(N__84063),
            .in2(_gnd_net_),
            .in3(N__84435),
            .lcout(pid_side_m78_0_a2_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_2_27_LC_15_12_4 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_2_27_LC_15_12_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_2_27_LC_15_12_4 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_2_27_LC_15_12_4  (
            .in0(N__85935),
            .in1(N__84576),
            .in2(_gnd_net_),
            .in3(N__87033),
            .lcout(),
            .ltout(\pid_side.error_i_reg_9_rn_0_27_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_27_LC_15_12_5 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_27_LC_15_12_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_27_LC_15_12_5 .LUT_INIT=16'b0101000001110010;
    LogicCell40 \pid_side.error_i_reg_esr_27_LC_15_12_5  (
            .in0(N__65413),
            .in1(N__80032),
            .in2(N__62974),
            .in3(N__62971),
            .lcout(\pid_side.error_i_regZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94157),
            .ce(N__86744),
            .sr(N__86436));
    defparam \pid_side.error_i_reg_esr_RNO_6_15_LC_15_12_6 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_6_15_LC_15_12_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_6_15_LC_15_12_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_6_15_LC_15_12_6  (
            .in0(N__84434),
            .in1(N__87408),
            .in2(N__84117),
            .in3(N__87031),
            .lcout(\pid_side.error_i_reg_9_sn_sn_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_14_LC_15_12_7 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_14_LC_15_12_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_14_LC_15_12_7 .LUT_INIT=16'b0001110000010000;
    LogicCell40 \pid_side.error_i_reg_esr_14_LC_15_12_7  (
            .in0(N__63061),
            .in1(N__66232),
            .in2(N__84577),
            .in3(N__66085),
            .lcout(\pid_side.error_i_regZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94157),
            .ce(N__86744),
            .sr(N__86436));
    defparam \pid_front.error_i_reg_esr_RNO_5_21_LC_15_13_0 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_5_21_LC_15_13_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_5_21_LC_15_13_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_5_21_LC_15_13_0  (
            .in0(N__82637),
            .in1(N__81403),
            .in2(N__89099),
            .in3(N__74504),
            .lcout(\pid_front.error_i_reg_esr_RNO_5Z0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.m24_2_03_0_o2_LC_15_13_1 .C_ON=1'b0;
    defparam \pid_side.m24_2_03_0_o2_LC_15_13_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.m24_2_03_0_o2_LC_15_13_1 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \pid_side.m24_2_03_0_o2_LC_15_13_1  (
            .in0(_gnd_net_),
            .in1(N__73404),
            .in2(_gnd_net_),
            .in3(N__80119),
            .lcout(pid_side_N_174),
            .ltout(pid_side_N_174_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_4_21_LC_15_13_2 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_4_21_LC_15_13_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_4_21_LC_15_13_2 .LUT_INIT=16'b0000000100000011;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_4_21_LC_15_13_2  (
            .in0(N__89073),
            .in1(N__82639),
            .in2(N__62935),
            .in3(N__74503),
            .lcout(\pid_front.error_i_reg_esr_RNO_4Z0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_ki_fast_fast_esr_3_LC_15_13_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_fast_fast_esr_3_LC_15_13_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_fast_fast_esr_3_LC_15_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_fast_fast_esr_3_LC_15_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__92329),
            .lcout(xy_ki_fast_fast_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94168),
            .ce(N__83900),
            .sr(N__86427));
    defparam \Commands_frame_decoder.source_xy_ki_fast_esr_2_LC_15_13_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_fast_esr_2_LC_15_13_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_fast_esr_2_LC_15_13_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_fast_esr_2_LC_15_13_4  (
            .in0(N__92514),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(xy_ki_fast_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94168),
            .ce(N__83900),
            .sr(N__86427));
    defparam \Commands_frame_decoder.source_xy_ki_fast_esr_3_LC_15_13_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_fast_esr_3_LC_15_13_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_fast_esr_3_LC_15_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_fast_esr_3_LC_15_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__92328),
            .lcout(xy_ki_fast_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94168),
            .ce(N__83900),
            .sr(N__86427));
    defparam \pid_side.m78_0_a2_5_LC_15_13_6 .C_ON=1'b0;
    defparam \pid_side.m78_0_a2_5_LC_15_13_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.m78_0_a2_5_LC_15_13_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \pid_side.m78_0_a2_5_LC_15_13_6  (
            .in0(N__80120),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78439),
            .lcout(pid_side_N_495),
            .ltout(pid_side_N_495_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_0_0_c_RNITALU1_LC_15_13_7 .C_ON=1'b0;
    defparam \pid_side.error_cry_0_0_c_RNITALU1_LC_15_13_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_0_c_RNITALU1_LC_15_13_7 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \pid_side.error_cry_0_0_c_RNITALU1_LC_15_13_7  (
            .in0(N__89077),
            .in1(N__82638),
            .in2(N__63022),
            .in3(N__80311),
            .lcout(\pid_side.N_543 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_0_c_RNI7VTI3_LC_15_14_0 .C_ON=1'b0;
    defparam \pid_side.error_cry_0_c_RNI7VTI3_LC_15_14_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_c_RNI7VTI3_LC_15_14_0 .LUT_INIT=16'b0100111101000010;
    LogicCell40 \pid_side.error_cry_0_c_RNI7VTI3_LC_15_14_0  (
            .in0(N__89068),
            .in1(N__62986),
            .in2(N__84134),
            .in3(N__83538),
            .lcout(\pid_side.m4_2_01 ),
            .ltout(\pid_side.m4_2_01_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_0_LC_15_14_1 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_0_LC_15_14_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_0_LC_15_14_1 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \pid_side.error_i_reg_0_LC_15_14_1  (
            .in0(N__65468),
            .in1(N__82078),
            .in2(N__63019),
            .in3(N__63005),
            .lcout(\pid_side.error_i_regZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94183),
            .ce(),
            .sr(N__86417));
    defparam \pid_side.error_cry_0_c_RNIMI671_LC_15_14_2 .C_ON=1'b0;
    defparam \pid_side.error_cry_0_c_RNIMI671_LC_15_14_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_c_RNIMI671_LC_15_14_2 .LUT_INIT=16'b0101010011110100;
    LogicCell40 \pid_side.error_cry_0_c_RNIMI671_LC_15_14_2  (
            .in0(N__82737),
            .in1(N__80940),
            .in2(N__90647),
            .in3(N__81023),
            .lcout(\pid_side.m4_2_01_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_0_c_RNINMCR_LC_15_14_3 .C_ON=1'b0;
    defparam \pid_side.error_cry_0_c_RNINMCR_LC_15_14_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_c_RNINMCR_LC_15_14_3 .LUT_INIT=16'b0101110100001100;
    LogicCell40 \pid_side.error_cry_0_c_RNINMCR_LC_15_14_3  (
            .in0(N__81024),
            .in1(N__89067),
            .in2(N__80949),
            .in3(N__82739),
            .lcout(),
            .ltout(\pid_side.m64_i_o2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_1_c_RNI6K4B1_LC_15_14_4 .C_ON=1'b0;
    defparam \pid_side.error_cry_1_c_RNI6K4B1_LC_15_14_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_1_c_RNI6K4B1_LC_15_14_4 .LUT_INIT=16'b1111100011111001;
    LogicCell40 \pid_side.error_cry_1_c_RNI6K4B1_LC_15_14_4  (
            .in0(N__87389),
            .in1(N__89819),
            .in2(N__62980),
            .in3(N__81111),
            .lcout(\pid_side.error_cry_1_c_RNI6K4BZ0Z1 ),
            .ltout(\pid_side.error_cry_1_c_RNI6K4BZ0Z1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_14_LC_15_14_5 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_14_LC_15_14_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_14_LC_15_14_5 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_14_LC_15_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__62977),
            .in3(N__84838),
            .lcout(\pid_side.N_111 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.m13_2_03_4_i_0_a2_3_0_LC_15_14_7 .C_ON=1'b0;
    defparam \pid_side.m13_2_03_4_i_0_a2_3_0_LC_15_14_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.m13_2_03_4_i_0_a2_3_0_LC_15_14_7 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \pid_side.m13_2_03_4_i_0_a2_3_0_LC_15_14_7  (
            .in0(N__89110),
            .in1(N__85158),
            .in2(_gnd_net_),
            .in3(N__82738),
            .lcout(pid_side_m13_2_03_4_i_0_a2_3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_0_11_LC_15_15_0 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_11_LC_15_15_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_11_LC_15_15_0 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_11_LC_15_15_0  (
            .in0(N__74935),
            .in1(N__83369),
            .in2(N__63034),
            .in3(N__63049),
            .lcout(\pid_front.m78_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_7_c_RNI8G5F1_LC_15_15_1 .C_ON=1'b0;
    defparam \pid_front.error_cry_7_c_RNI8G5F1_LC_15_15_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_7_c_RNI8G5F1_LC_15_15_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \pid_front.error_cry_7_c_RNI8G5F1_LC_15_15_1  (
            .in0(N__78468),
            .in1(N__74318),
            .in2(_gnd_net_),
            .in3(N__79883),
            .lcout(\pid_front.N_161 ),
            .ltout(\pid_front.N_161_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_2_11_LC_15_15_2 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_2_11_LC_15_15_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_2_11_LC_15_15_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_2_11_LC_15_15_2  (
            .in0(N__84119),
            .in1(N__87779),
            .in2(N__63052),
            .in3(N__83368),
            .lcout(\pid_front.N_398 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_1_11_LC_15_15_3 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_1_11_LC_15_15_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_1_11_LC_15_15_3 .LUT_INIT=16'b1100110011101100;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_1_11_LC_15_15_3  (
            .in0(N__83370),
            .in1(N__66007),
            .in2(N__85769),
            .in3(N__66193),
            .lcout(),
            .ltout(\pid_front.m78_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_11_LC_15_15_4 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_11_LC_15_15_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_11_LC_15_15_4 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \pid_front.error_i_reg_esr_11_LC_15_15_4  (
            .in0(N__68670),
            .in1(N__63043),
            .in2(N__63037),
            .in3(N__63241),
            .lcout(\pid_front.error_i_regZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94195),
            .ce(N__78014),
            .sr(N__86406));
    defparam \pid_front.error_cry_2_0_c_RNIVKQ02_LC_15_15_5 .C_ON=1'b0;
    defparam \pid_front.error_cry_2_0_c_RNIVKQ02_LC_15_15_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_2_0_c_RNIVKQ02_LC_15_15_5 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \pid_front.error_cry_2_0_c_RNIVKQ02_LC_15_15_5  (
            .in0(N__82756),
            .in1(N__77853),
            .in2(N__90657),
            .in3(N__77722),
            .lcout(\pid_front.N_626 ),
            .ltout(\pid_front.N_626_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_3_c_RNI2H9H3_LC_15_15_6 .C_ON=1'b0;
    defparam \pid_front.error_cry_3_c_RNI2H9H3_LC_15_15_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_3_c_RNI2H9H3_LC_15_15_6 .LUT_INIT=16'b1111001000000000;
    LogicCell40 \pid_front.error_cry_3_c_RNI2H9H3_LC_15_15_6  (
            .in0(N__79884),
            .in1(N__87778),
            .in2(N__63025),
            .in3(N__83506),
            .lcout(\pid_front.N_576 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_c_RNICF3L2_LC_15_16_1 .C_ON=1'b0;
    defparam \pid_front.error_cry_0_c_RNICF3L2_LC_15_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_c_RNICF3L2_LC_15_16_1 .LUT_INIT=16'b1111000010000000;
    LogicCell40 \pid_front.error_cry_0_c_RNICF3L2_LC_15_16_1  (
            .in0(N__74175),
            .in1(N__74964),
            .in2(N__76868),
            .in3(N__66071),
            .lcout(\pid_front.N_556 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_0_6_LC_15_16_3 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_6_LC_15_16_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_6_LC_15_16_3 .LUT_INIT=16'b1111100011111000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_6_LC_15_16_3  (
            .in0(N__81312),
            .in1(N__63156),
            .in2(N__63130),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\pid_front.error_i_reg_esr_RNO_0Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_6_LC_15_16_4 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_6_LC_15_16_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_6_LC_15_16_4 .LUT_INIT=16'b1100110011000000;
    LogicCell40 \pid_front.error_i_reg_esr_6_LC_15_16_4  (
            .in0(_gnd_net_),
            .in1(N__83355),
            .in2(N__63190),
            .in3(N__63166),
            .lcout(\pid_front.error_i_regZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94212),
            .ce(N__78106),
            .sr(N__86397));
    defparam \pid_front.error_cry_2_c_RNI8A755_LC_15_16_5 .C_ON=1'b0;
    defparam \pid_front.error_cry_2_c_RNI8A755_LC_15_16_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_2_c_RNI8A755_LC_15_16_5 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \pid_front.error_cry_2_c_RNI8A755_LC_15_16_5  (
            .in0(N__74638),
            .in1(N__63187),
            .in2(N__69508),
            .in3(N__73631),
            .lcout(\pid_front.m10_2_03_3_i_0_o2_0 ),
            .ltout(\pid_front.m10_2_03_3_i_0_o2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_1_22_LC_15_16_6 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_1_22_LC_15_16_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_1_22_LC_15_16_6 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_1_22_LC_15_16_6  (
            .in0(N__63155),
            .in1(N__63126),
            .in2(N__63118),
            .in3(N__81313),
            .lcout(),
            .ltout(\pid_front.m10_2_03_3_i_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_22_LC_15_16_7 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_22_LC_15_16_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_22_LC_15_16_7 .LUT_INIT=16'b1100010010000000;
    LogicCell40 \pid_front.error_i_reg_esr_22_LC_15_16_7  (
            .in0(N__84564),
            .in1(N__87047),
            .in2(N__63115),
            .in3(N__63112),
            .lcout(\pid_front.error_i_regZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94212),
            .ce(N__78106),
            .sr(N__86397));
    defparam \pid_front.error_cry_3_0_c_RNI50IA3_LC_15_17_0 .C_ON=1'b0;
    defparam \pid_front.error_cry_3_0_c_RNI50IA3_LC_15_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_3_0_c_RNI50IA3_LC_15_17_0 .LUT_INIT=16'b1110000011000000;
    LogicCell40 \pid_front.error_cry_3_0_c_RNI50IA3_LC_15_17_0  (
            .in0(N__76864),
            .in1(N__63103),
            .in2(N__83527),
            .in3(N__74849),
            .lcout(),
            .ltout(\pid_front.N_554_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_0_c_RNISRSC6_LC_15_17_1 .C_ON=1'b0;
    defparam \pid_front.error_cry_0_0_c_RNISRSC6_LC_15_17_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_0_c_RNISRSC6_LC_15_17_1 .LUT_INIT=16'b1111110111111100;
    LogicCell40 \pid_front.error_cry_0_0_c_RNISRSC6_LC_15_17_1  (
            .in0(N__81442),
            .in1(N__63088),
            .in2(N__63091),
            .in3(N__69580),
            .lcout(\pid_front.m13_2_03_4_i_0_o2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_0_c_RNI4QFK1_LC_15_17_2 .C_ON=1'b0;
    defparam \pid_front.error_cry_0_0_c_RNI4QFK1_LC_15_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_0_c_RNI4QFK1_LC_15_17_2 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \pid_front.error_cry_0_0_c_RNI4QFK1_LC_15_17_2  (
            .in0(N__74963),
            .in1(N__83026),
            .in2(N__90658),
            .in3(N__77973),
            .lcout(\pid_front.N_543 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_7_c_RNI07ND4_LC_15_17_3 .C_ON=1'b0;
    defparam \pid_front.error_cry_7_c_RNI07ND4_LC_15_17_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_7_c_RNI07ND4_LC_15_17_3 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \pid_front.error_cry_7_c_RNI07ND4_LC_15_17_3  (
            .in0(N__76865),
            .in1(N__74332),
            .in2(N__63082),
            .in3(N__77079),
            .lcout(\pid_front.m13_2_03_4_i_0_o2_2 ),
            .ltout(\pid_front.m13_2_03_4_i_0_o2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_0_9_LC_15_17_4 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_9_LC_15_17_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_9_LC_15_17_4 .LUT_INIT=16'b1111110011110000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_9_LC_15_17_4  (
            .in0(_gnd_net_),
            .in1(N__69491),
            .in2(N__63274),
            .in3(N__74717),
            .lcout(),
            .ltout(\pid_front.error_i_reg_esr_RNO_0Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_9_LC_15_17_5 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_9_LC_15_17_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_9_LC_15_17_5 .LUT_INIT=16'b1100110011000000;
    LogicCell40 \pid_front.error_i_reg_esr_9_LC_15_17_5  (
            .in0(_gnd_net_),
            .in1(N__83377),
            .in2(N__63271),
            .in3(N__63267),
            .lcout(\pid_front.error_i_regZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94228),
            .ce(N__78141),
            .sr(N__86387));
    defparam \pid_front.error_i_reg_esr_RNO_1_27_LC_15_18_0 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_1_27_LC_15_18_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_1_27_LC_15_18_0 .LUT_INIT=16'b0001010100010000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_1_27_LC_15_18_0  (
            .in0(N__87447),
            .in1(N__74716),
            .in2(N__84182),
            .in3(N__74677),
            .lcout(\pid_front.N_339 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_5_c_RNI9J5J2_LC_15_18_2 .C_ON=1'b0;
    defparam \pid_front.error_cry_5_c_RNI9J5J2_LC_15_18_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_5_c_RNI9J5J2_LC_15_18_2 .LUT_INIT=16'b0011111000110010;
    LogicCell40 \pid_front.error_cry_5_c_RNI9J5J2_LC_15_18_2  (
            .in0(N__78396),
            .in1(N__73291),
            .in2(N__85179),
            .in3(N__74506),
            .lcout(\pid_front.N_184 ),
            .ltout(\pid_front.N_184_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_3_0_c_RNIK8ST3_LC_15_18_3 .C_ON=1'b0;
    defparam \pid_front.error_cry_3_0_c_RNIK8ST3_LC_15_18_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_3_0_c_RNIK8ST3_LC_15_18_3 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \pid_front.error_cry_3_0_c_RNIK8ST3_LC_15_18_3  (
            .in0(N__89755),
            .in1(N__89112),
            .in2(N__63256),
            .in3(N__66216),
            .lcout(\pid_front.N_229 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_c_RNICF3L2_0_LC_15_18_4 .C_ON=1'b0;
    defparam \pid_front.error_cry_0_c_RNICF3L2_0_LC_15_18_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_c_RNICF3L2_0_LC_15_18_4 .LUT_INIT=16'b1110000011000000;
    LogicCell40 \pid_front.error_cry_0_c_RNICF3L2_0_LC_15_18_4  (
            .in0(N__74965),
            .in1(N__66064),
            .in2(N__85775),
            .in3(N__74164),
            .lcout(),
            .ltout(\pid_front.N_575_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_c_RNI86D9A_LC_15_18_5 .C_ON=1'b0;
    defparam \pid_front.error_cry_0_c_RNI86D9A_LC_15_18_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_c_RNI86D9A_LC_15_18_5 .LUT_INIT=16'b1111110111111100;
    LogicCell40 \pid_front.error_cry_0_c_RNI86D9A_LC_15_18_5  (
            .in0(N__84178),
            .in1(N__63253),
            .in2(N__63244),
            .in3(N__63237),
            .lcout(\pid_front.m11_2_03_3_i_3 ),
            .ltout(\pid_front.m11_2_03_3_i_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_7_LC_15_18_6 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_7_LC_15_18_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_7_LC_15_18_6 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \pid_front.error_i_reg_7_LC_15_18_6  (
            .in0(N__82129),
            .in1(N__83365),
            .in2(N__63220),
            .in3(N__63306),
            .lcout(\pid_front.error_i_regZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94244),
            .ce(),
            .sr(N__86379));
    defparam \pid_front.error_i_reg_esr_RNII1MD_0_LC_15_19_0 .C_ON=1'b1;
    defparam \pid_front.error_i_reg_esr_RNII1MD_0_LC_15_19_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNII1MD_0_LC_15_19_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNII1MD_0_LC_15_19_0  (
            .in0(_gnd_net_),
            .in1(N__66366),
            .in2(N__66282),
            .in3(_gnd_net_),
            .lcout(\pid_front.un1_pid_prereg_0 ),
            .ltout(),
            .carryin(bfn_15_19_0_),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_0_c_RNI9AGE_LC_15_19_1 .C_ON=1'b1;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_0_c_RNI9AGE_LC_15_19_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_0_c_RNI9AGE_LC_15_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_0_c_RNI9AGE_LC_15_19_1  (
            .in0(_gnd_net_),
            .in1(N__66517),
            .in2(N__66424),
            .in3(N__63352),
            .lcout(\pid_front.un1_error_i_acumm_prereg_cry_0_c_RNI9AGE ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_0 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_1_c_RNICEHE_LC_15_19_2 .C_ON=1'b1;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_1_c_RNICEHE_LC_15_19_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_1_c_RNICEHE_LC_15_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_1_c_RNICEHE_LC_15_19_2  (
            .in0(_gnd_net_),
            .in1(N__66502),
            .in2(N__66433),
            .in3(N__63349),
            .lcout(\pid_front.un1_error_i_acumm_prereg_cry_1_c_RNICEHE ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_1 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_2_c_RNI68OM_LC_15_19_3 .C_ON=1'b1;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_2_c_RNI68OM_LC_15_19_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_2_c_RNI68OM_LC_15_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_2_c_RNI68OM_LC_15_19_3  (
            .in0(_gnd_net_),
            .in1(N__81991),
            .in2(N__66583),
            .in3(N__63346),
            .lcout(\pid_front.un1_error_i_acumm_prereg_cry_2_c_RNI68OM ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_2 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_3_c_RNI9CPM_LC_15_19_4 .C_ON=1'b1;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_3_c_RNI9CPM_LC_15_19_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_3_c_RNI9CPM_LC_15_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_3_c_RNI9CPM_LC_15_19_4  (
            .in0(_gnd_net_),
            .in1(N__73597),
            .in2(N__66460),
            .in3(N__63343),
            .lcout(\pid_front.un1_error_i_acumm_prereg_cry_3_c_RNI9CPM ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_3 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_4_c_RNICGQM_LC_15_19_5 .C_ON=1'b1;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_4_c_RNICGQM_LC_15_19_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_4_c_RNICGQM_LC_15_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_4_c_RNICGQM_LC_15_19_5  (
            .in0(_gnd_net_),
            .in1(N__66487),
            .in2(N__63340),
            .in3(N__63322),
            .lcout(\pid_front.un1_error_i_acumm_prereg_cry_4_c_RNICGQM ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_4 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_5_c_RNIOULE_LC_15_19_6 .C_ON=1'b1;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_5_c_RNIOULE_LC_15_19_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_5_c_RNIOULE_LC_15_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_5_c_RNIOULE_LC_15_19_6  (
            .in0(_gnd_net_),
            .in1(N__63319),
            .in2(N__66496),
            .in3(N__63310),
            .lcout(\pid_front.un1_error_i_acumm_prereg_cry_5_c_RNIOULE ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_5 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_6_c_RNIIOSM_LC_15_19_7 .C_ON=1'b1;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_6_c_RNIIOSM_LC_15_19_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_6_c_RNIIOSM_LC_15_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_6_c_RNIIOSM_LC_15_19_7  (
            .in0(_gnd_net_),
            .in1(N__66598),
            .in2(N__63307),
            .in3(N__63292),
            .lcout(\pid_front.un1_error_i_acumm_prereg_cry_6_c_RNIIOSM ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_6 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_7_c_RNIU6OE_LC_15_20_0 .C_ON=1'b1;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_7_c_RNIU6OE_LC_15_20_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_7_c_RNIU6OE_LC_15_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_7_c_RNIU6OE_LC_15_20_0  (
            .in0(_gnd_net_),
            .in1(N__66592),
            .in2(N__63289),
            .in3(N__63277),
            .lcout(\pid_front.un1_error_i_acumm_prereg_cry_7_c_RNIU6OE ),
            .ltout(),
            .carryin(bfn_15_20_0_),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_8_c_RNI1BPE_LC_15_20_1 .C_ON=1'b1;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_8_c_RNI1BPE_LC_15_20_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_8_c_RNI1BPE_LC_15_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_8_c_RNI1BPE_LC_15_20_1  (
            .in0(_gnd_net_),
            .in1(N__70129),
            .in2(N__63421),
            .in3(N__63409),
            .lcout(\pid_front.un1_error_i_acumm_prereg_cry_8_c_RNI1BPE ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_8 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_9_c_RNIIPQK_LC_15_20_2 .C_ON=1'b1;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_9_c_RNIIPQK_LC_15_20_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_9_c_RNIIPQK_LC_15_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_9_c_RNIIPQK_LC_15_20_2  (
            .in0(_gnd_net_),
            .in1(N__75070),
            .in2(N__63406),
            .in3(N__63391),
            .lcout(\pid_front.un1_error_i_acumm_prereg_cry_9_c_RNIIPQK ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_9 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNIS09U_11_LC_15_20_3 .C_ON=1'b1;
    defparam \pid_front.error_i_reg_esr_RNIS09U_11_LC_15_20_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNIS09U_11_LC_15_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNIS09U_11_LC_15_20_3  (
            .in0(_gnd_net_),
            .in1(N__74980),
            .in2(N__63388),
            .in3(N__63373),
            .lcout(\pid_front.error_i_reg_esr_RNIS09UZ0Z_11 ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_10 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNIV4AU_12_LC_15_20_4 .C_ON=1'b1;
    defparam \pid_front.error_i_reg_esr_RNIV4AU_12_LC_15_20_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNIV4AU_12_LC_15_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNIV4AU_12_LC_15_20_4  (
            .in0(_gnd_net_),
            .in1(N__75781),
            .in2(N__69739),
            .in3(N__63370),
            .lcout(\pid_front.error_i_reg_esr_RNIV4AUZ0Z_12 ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_11 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNI29BU_13_LC_15_20_5 .C_ON=1'b1;
    defparam \pid_front.error_i_reg_esr_RNI29BU_13_LC_15_20_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNI29BU_13_LC_15_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNI29BU_13_LC_15_20_5  (
            .in0(_gnd_net_),
            .in1(N__63673),
            .in2(N__74737),
            .in3(N__63367),
            .lcout(\pid_front.error_i_reg_esr_RNI29BUZ0Z_13 ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_12 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNI4CCU_14_LC_15_20_6 .C_ON=1'b1;
    defparam \pid_front.error_i_reg_esr_RNI4CCU_14_LC_15_20_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNI4CCU_14_LC_15_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNI4CCU_14_LC_15_20_6  (
            .in0(_gnd_net_),
            .in1(N__69721),
            .in2(N__63703),
            .in3(N__63364),
            .lcout(\pid_front.error_i_reg_esr_RNI4CCUZ0Z_14 ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_13 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNI6FDU_15_LC_15_20_7 .C_ON=1'b1;
    defparam \pid_front.error_i_reg_esr_RNI6FDU_15_LC_15_20_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNI6FDU_15_LC_15_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNI6FDU_15_LC_15_20_7  (
            .in0(_gnd_net_),
            .in1(N__63677),
            .in2(N__73942),
            .in3(N__63361),
            .lcout(\pid_front.error_i_reg_esr_RNI6FDUZ0Z_15 ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_14 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNI8IEU_16_LC_15_21_0 .C_ON=1'b1;
    defparam \pid_front.error_i_reg_esr_RNI8IEU_16_LC_15_21_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNI8IEU_16_LC_15_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNI8IEU_16_LC_15_21_0  (
            .in0(_gnd_net_),
            .in1(N__63678),
            .in2(N__69826),
            .in3(N__63358),
            .lcout(\pid_front.error_i_reg_esr_RNI8IEUZ0Z_16 ),
            .ltout(),
            .carryin(bfn_15_21_0_),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNIALFU_17_LC_15_21_1 .C_ON=1'b1;
    defparam \pid_front.error_i_reg_esr_RNIALFU_17_LC_15_21_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNIALFU_17_LC_15_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNIALFU_17_LC_15_21_1  (
            .in0(_gnd_net_),
            .in1(N__69619),
            .in2(N__63704),
            .in3(N__63355),
            .lcout(\pid_front.error_i_reg_esr_RNIALFUZ0Z_17 ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_16 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNICOGU_18_LC_15_21_2 .C_ON=1'b1;
    defparam \pid_front.error_i_reg_esr_RNICOGU_18_LC_15_21_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNICOGU_18_LC_15_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNICOGU_18_LC_15_21_2  (
            .in0(_gnd_net_),
            .in1(N__63682),
            .in2(N__63535),
            .in3(N__63526),
            .lcout(\pid_front.error_i_reg_esr_RNICOGUZ0Z_18 ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_17 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNIERHU_19_LC_15_21_3 .C_ON=1'b1;
    defparam \pid_front.error_i_reg_esr_RNIERHU_19_LC_15_21_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNIERHU_19_LC_15_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNIERHU_19_LC_15_21_3  (
            .in0(_gnd_net_),
            .in1(N__78163),
            .in2(N__63705),
            .in3(N__63523),
            .lcout(\pid_front.error_i_reg_esr_RNIERHUZ0Z_19 ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_18 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNI7MJU_20_LC_15_21_4 .C_ON=1'b1;
    defparam \pid_front.error_i_reg_esr_RNI7MJU_20_LC_15_21_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNI7MJU_20_LC_15_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNI7MJU_20_LC_15_21_4  (
            .in0(_gnd_net_),
            .in1(N__63686),
            .in2(N__66304),
            .in3(N__63520),
            .lcout(\pid_front.error_i_reg_esr_RNI7MJUZ0Z_20 ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_19 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNI08DV_21_LC_15_21_5 .C_ON=1'b1;
    defparam \pid_front.error_i_reg_esr_RNI08DV_21_LC_15_21_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNI08DV_21_LC_15_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNI08DV_21_LC_15_21_5  (
            .in0(_gnd_net_),
            .in1(N__63517),
            .in2(N__63706),
            .in3(N__63505),
            .lcout(\pid_front.error_i_reg_esr_RNI08DVZ0Z_21 ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_20 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNI2BEV_22_LC_15_21_6 .C_ON=1'b1;
    defparam \pid_front.error_i_reg_esr_RNI2BEV_22_LC_15_21_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNI2BEV_22_LC_15_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNI2BEV_22_LC_15_21_6  (
            .in0(_gnd_net_),
            .in1(N__63690),
            .in2(N__63502),
            .in3(N__63487),
            .lcout(\pid_front.error_i_reg_esr_RNI2BEVZ0Z_22 ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_21 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNI4EFV_23_LC_15_21_7 .C_ON=1'b1;
    defparam \pid_front.error_i_reg_esr_RNI4EFV_23_LC_15_21_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNI4EFV_23_LC_15_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNI4EFV_23_LC_15_21_7  (
            .in0(_gnd_net_),
            .in1(N__63484),
            .in2(N__63707),
            .in3(N__63475),
            .lcout(\pid_front.error_i_reg_esr_RNI4EFVZ0Z_23 ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_22 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNI6HGV_24_LC_15_22_0 .C_ON=1'b1;
    defparam \pid_front.error_i_reg_esr_RNI6HGV_24_LC_15_22_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNI6HGV_24_LC_15_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNI6HGV_24_LC_15_22_0  (
            .in0(_gnd_net_),
            .in1(N__63694),
            .in2(N__63472),
            .in3(N__63457),
            .lcout(\pid_front.error_i_reg_esr_RNI6HGVZ0Z_24 ),
            .ltout(),
            .carryin(bfn_15_22_0_),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNI8KHV_25_LC_15_22_1 .C_ON=1'b1;
    defparam \pid_front.error_i_reg_esr_RNI8KHV_25_LC_15_22_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNI8KHV_25_LC_15_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNI8KHV_25_LC_15_22_1  (
            .in0(_gnd_net_),
            .in1(N__63454),
            .in2(N__63708),
            .in3(N__63442),
            .lcout(\pid_front.error_i_reg_esr_RNI8KHVZ0Z_25 ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_24 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNIANIV_26_LC_15_22_2 .C_ON=1'b1;
    defparam \pid_front.error_i_reg_esr_RNIANIV_26_LC_15_22_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNIANIV_26_LC_15_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNIANIV_26_LC_15_22_2  (
            .in0(_gnd_net_),
            .in1(N__63698),
            .in2(N__63439),
            .in3(N__63424),
            .lcout(\pid_front.error_i_reg_esr_RNIANIVZ0Z_26 ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_25 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_26_c_RNICQJV_LC_15_22_3 .C_ON=1'b1;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_26_c_RNICQJV_LC_15_22_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_26_c_RNICQJV_LC_15_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_26_c_RNICQJV_LC_15_22_3  (
            .in0(_gnd_net_),
            .in1(N__66156),
            .in2(N__63709),
            .in3(N__63712),
            .lcout(\pid_front.un1_error_i_acumm_prereg_cry_26_c_RNICQJV ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_26 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_27_c_RNIDSKV_LC_15_22_4 .C_ON=1'b0;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_27_c_RNIDSKV_LC_15_22_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_27_c_RNIDSKV_LC_15_22_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_27_c_RNIDSKV_LC_15_22_4  (
            .in0(N__66157),
            .in1(N__63702),
            .in2(_gnd_net_),
            .in3(N__63619),
            .lcout(\pid_front.un1_error_i_acumm_prereg_cry_27_c_RNIDSKV ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_28_LC_15_22_5 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_28_LC_15_22_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_28_LC_15_22_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_28_LC_15_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66835),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94311),
            .ce(N__75324),
            .sr(N__86362));
    defparam \pid_front.error_p_reg_esr_RNIO4E8_0_2_LC_15_23_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIO4E8_0_2_LC_15_23_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIO4E8_0_2_LC_15_23_0 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_p_reg_esr_RNIO4E8_0_2_LC_15_23_0  (
            .in0(N__63594),
            .in1(N__63582),
            .in2(_gnd_net_),
            .in3(N__81923),
            .lcout(\pid_front.error_p_reg_esr_RNIO4E8_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_2_LC_15_23_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_2_LC_15_23_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_2_LC_15_23_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_2_LC_15_23_1  (
            .in0(N__81925),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prevZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94328),
            .ce(N__71794),
            .sr(N__71699));
    defparam \pid_front.error_p_reg_esr_RNIO4E8_2_LC_15_23_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIO4E8_2_LC_15_23_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIO4E8_2_LC_15_23_2 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_front.error_p_reg_esr_RNIO4E8_2_LC_15_23_2  (
            .in0(N__63595),
            .in1(N__63583),
            .in2(_gnd_net_),
            .in3(N__81924),
            .lcout(\pid_front.error_p_reg_esr_RNIO4E8Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIQ9C61_0_17_LC_15_23_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIQ9C61_0_17_LC_15_23_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIQ9C61_0_17_LC_15_23_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_p_reg_esr_RNIQ9C61_0_17_LC_15_23_3  (
            .in0(N__63564),
            .in1(N__63543),
            .in2(_gnd_net_),
            .in3(N__94433),
            .lcout(\pid_front.error_p_reg_esr_RNIQ9C61_0Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_17_LC_15_23_4 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_17_LC_15_23_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_17_LC_15_23_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_17_LC_15_23_4  (
            .in0(N__94435),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prevZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94328),
            .ce(N__71794),
            .sr(N__71699));
    defparam \pid_front.error_p_reg_esr_RNIQ9C61_17_LC_15_23_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIQ9C61_17_LC_15_23_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIQ9C61_17_LC_15_23_5 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_front.error_p_reg_esr_RNIQ9C61_17_LC_15_23_5  (
            .in0(N__63565),
            .in1(N__63544),
            .in2(_gnd_net_),
            .in3(N__94434),
            .lcout(\pid_front.error_p_reg_esr_RNIQ9C61Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNITCC61_0_18_LC_15_23_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNITCC61_0_18_LC_15_23_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNITCC61_0_18_LC_15_23_6 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_p_reg_esr_RNITCC61_0_18_LC_15_23_6  (
            .in0(N__76188),
            .in1(N__81956),
            .in2(_gnd_net_),
            .in3(N__76158),
            .lcout(\pid_front.error_p_reg_esr_RNITCC61_0Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_18_LC_15_23_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_18_LC_15_23_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_18_LC_15_23_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_18_LC_15_23_7  (
            .in0(N__81957),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prevZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94328),
            .ce(N__71794),
            .sr(N__71699));
    defparam \pid_front.error_p_reg_esr_RNIKG5U_0_10_LC_15_24_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIKG5U_0_10_LC_15_24_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIKG5U_0_10_LC_15_24_0 .LUT_INIT=16'b1000111010101111;
    LogicCell40 \pid_front.error_p_reg_esr_RNIKG5U_0_10_LC_15_24_0  (
            .in0(N__70395),
            .in1(N__78727),
            .in2(N__81898),
            .in3(N__71360),
            .lcout(),
            .ltout(\pid_front.error_p_reg_esr_RNIKG5U_0Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNI379B2_10_LC_15_24_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNI379B2_10_LC_15_24_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNI379B2_10_LC_15_24_1 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNI379B2_10_LC_15_24_1  (
            .in0(_gnd_net_),
            .in1(N__70277),
            .in2(N__63769),
            .in3(N__63748),
            .lcout(\pid_front.error_d_reg_prev_esr_RNI379B2Z0Z_10 ),
            .ltout(\pid_front.error_d_reg_prev_esr_RNI379B2Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNI5JRF4_0_10_LC_15_24_2 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNI5JRF4_0_10_LC_15_24_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNI5JRF4_0_10_LC_15_24_2 .LUT_INIT=16'b1011010001001011;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNI5JRF4_0_10_LC_15_24_2  (
            .in0(N__81894),
            .in1(N__70281),
            .in2(N__63766),
            .in3(N__67155),
            .lcout(\pid_front.error_d_reg_prev_esr_RNI5JRF4_0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIKG5U_10_LC_15_24_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIKG5U_10_LC_15_24_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIKG5U_10_LC_15_24_3 .LUT_INIT=16'b1111110111000100;
    LogicCell40 \pid_front.error_p_reg_esr_RNIKG5U_10_LC_15_24_3  (
            .in0(N__71359),
            .in1(N__81890),
            .in2(N__78736),
            .in3(N__70394),
            .lcout(\pid_front.error_p_reg_esr_RNIKG5UZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIK2AG3_12_LC_15_24_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIK2AG3_12_LC_15_24_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIK2AG3_12_LC_15_24_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_front.error_p_reg_esr_RNIK2AG3_12_LC_15_24_4  (
            .in0(_gnd_net_),
            .in1(N__67209),
            .in2(_gnd_net_),
            .in3(N__75695),
            .lcout(\pid_front.un1_pid_prereg_153_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIEAU52_21_LC_15_24_5 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIEAU52_21_LC_15_24_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIEAU52_21_LC_15_24_5 .LUT_INIT=16'b1110111100001000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIEAU52_21_LC_15_24_5  (
            .in0(N__91757),
            .in1(N__66703),
            .in2(N__67070),
            .in3(N__72132),
            .lcout(\pid_front.un1_pid_prereg_0_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNI5JRF4_10_LC_15_24_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNI5JRF4_10_LC_15_24_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNI5JRF4_10_LC_15_24_6 .LUT_INIT=16'b1110111110001100;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNI5JRF4_10_LC_15_24_6  (
            .in0(N__81895),
            .in1(N__67156),
            .in2(N__70282),
            .in3(N__63724),
            .lcout(\pid_front.error_d_reg_prev_esr_RNI5JRF4Z0Z_10 ),
            .ltout(\pid_front.error_d_reg_prev_esr_RNI5JRF4Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIEU1SD_12_LC_15_24_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIEU1SD_12_LC_15_24_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIEU1SD_12_LC_15_24_7 .LUT_INIT=16'b1110100011101000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIEU1SD_12_LC_15_24_7  (
            .in0(N__75696),
            .in1(N__67210),
            .in2(N__63931),
            .in3(N__64014),
            .lcout(\pid_front.error_p_reg_esr_RNIEU1SDZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIN6C61_16_LC_15_25_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIN6C61_16_LC_15_25_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIN6C61_16_LC_15_25_0 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_front.error_p_reg_esr_RNIN6C61_16_LC_15_25_0  (
            .in0(N__63808),
            .in1(N__63778),
            .in2(_gnd_net_),
            .in3(N__94464),
            .lcout(\pid_front.error_p_reg_esr_RNIN6C61Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIUKHM6_16_LC_15_25_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIUKHM6_16_LC_15_25_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIUKHM6_16_LC_15_25_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIUKHM6_16_LC_15_25_1  (
            .in0(N__63858),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63942),
            .lcout(\pid_front.error_p_reg_esr_RNIUKHM6Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI3F9B3_17_LC_15_25_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI3F9B3_17_LC_15_25_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI3F9B3_17_LC_15_25_2 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_front.error_p_reg_esr_RNI3F9B3_17_LC_15_25_2  (
            .in0(N__63976),
            .in1(N__63994),
            .in2(_gnd_net_),
            .in3(N__63961),
            .lcout(\pid_front.un1_pid_prereg_0_6 ),
            .ltout(\pid_front.un1_pid_prereg_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNICS5DD_16_LC_15_25_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNICS5DD_16_LC_15_25_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNICS5DD_16_LC_15_25_3 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pid_front.error_p_reg_esr_RNICS5DD_16_LC_15_25_3  (
            .in0(N__63859),
            .in1(N__72033),
            .in2(N__63901),
            .in3(N__63943),
            .lcout(\pid_front.error_p_reg_esr_RNICS5DDZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIR58B3_16_LC_15_25_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIR58B3_16_LC_15_25_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIR58B3_16_LC_15_25_4 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIR58B3_16_LC_15_25_4  (
            .in0(N__63889),
            .in1(N__63871),
            .in2(_gnd_net_),
            .in3(N__71224),
            .lcout(\pid_front.un1_pid_prereg_0_4 ),
            .ltout(\pid_front.un1_pid_prereg_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNICN0DD_15_LC_15_25_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNICN0DD_15_LC_15_25_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNICN0DD_15_LC_15_25_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_front.error_p_reg_esr_RNICN0DD_15_LC_15_25_5  (
            .in0(N__63850),
            .in1(N__63838),
            .in2(N__63820),
            .in3(N__63941),
            .lcout(\pid_front.error_p_reg_esr_RNICN0DDZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIN6C61_0_16_LC_15_25_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIN6C61_0_16_LC_15_25_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIN6C61_0_16_LC_15_25_6 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_p_reg_esr_RNIN6C61_0_16_LC_15_25_6  (
            .in0(N__63807),
            .in1(N__63777),
            .in2(_gnd_net_),
            .in3(N__94463),
            .lcout(\pid_front.error_p_reg_esr_RNIN6C61_0Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_16_LC_15_25_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_16_LC_15_25_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_16_LC_15_25_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_16_LC_15_25_7  (
            .in0(N__94465),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prevZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94357),
            .ce(N__71804),
            .sr(N__71700));
    defparam \pid_front.error_i_acumm_prereg_esr_RNICMI41_0_13_LC_15_26_0 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNICMI41_0_13_LC_15_26_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNICMI41_0_13_LC_15_26_0 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNICMI41_0_13_LC_15_26_0  (
            .in0(N__64062),
            .in1(N__64095),
            .in2(N__64029),
            .in3(N__64104),
            .lcout(\pid_front.error_i_acumm_13_i_o2_0_10_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_13_LC_15_26_1 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_13_LC_15_26_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_13_LC_15_26_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_13_LC_15_26_1  (
            .in0(N__64397),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94367),
            .ce(N__75319),
            .sr(N__86353));
    defparam \pid_front.error_i_acumm_prereg_esr_RNICMI41_13_LC_15_26_2 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNICMI41_13_LC_15_26_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNICMI41_13_LC_15_26_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNICMI41_13_LC_15_26_2  (
            .in0(N__64063),
            .in1(N__64096),
            .in2(N__64030),
            .in3(N__64105),
            .lcout(\pid_front.error_i_acumm_13_i_o2_0_10_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_18_LC_15_26_3 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_18_LC_15_26_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_18_LC_15_26_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_18_LC_15_26_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63960),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94367),
            .ce(N__75319),
            .sr(N__86353));
    defparam \pid_front.error_i_acumm_prereg_esr_25_LC_15_26_4 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_25_LC_15_26_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_25_LC_15_26_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_25_LC_15_26_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64087),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94367),
            .ce(N__75319),
            .sr(N__86353));
    defparam \pid_front.error_i_acumm_prereg_esr_26_LC_15_26_5 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_26_LC_15_26_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_26_LC_15_26_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_26_LC_15_26_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64054),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94367),
            .ce(N__75319),
            .sr(N__86353));
    defparam \pid_front.error_d_reg_prev_esr_RNIL8SR5_12_LC_15_26_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIL8SR5_12_LC_15_26_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIL8SR5_12_LC_15_26_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIL8SR5_12_LC_15_26_6  (
            .in0(_gnd_net_),
            .in1(N__64396),
            .in2(_gnd_net_),
            .in3(N__67221),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIL8SR5Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI3F9B3_0_17_LC_15_26_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI3F9B3_0_17_LC_15_26_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI3F9B3_0_17_LC_15_26_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_p_reg_esr_RNI3F9B3_0_17_LC_15_26_7  (
            .in0(N__63993),
            .in1(N__63975),
            .in2(_gnd_net_),
            .in3(N__63959),
            .lcout(\pid_front.un1_pid_prereg_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_fast_esr_RNIR9PO_0_13_LC_15_27_0 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_fast_esr_RNIR9PO_0_13_LC_15_27_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_fast_esr_RNIR9PO_0_13_LC_15_27_0 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_d_reg_fast_esr_RNIR9PO_0_13_LC_15_27_0  (
            .in0(N__67692),
            .in1(N__67633),
            .in2(_gnd_net_),
            .in3(N__67599),
            .lcout(\pid_front.error_d_reg_fast_esr_RNIR9PO_0Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_fast_esr_13_LC_15_27_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_fast_esr_13_LC_15_27_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_fast_esr_13_LC_15_27_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_fast_esr_13_LC_15_27_1  (
            .in0(N__64231),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_fastZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94374),
            .ce(N__93370),
            .sr(N__93005));
    defparam \pid_front.error_d_reg_esr_13_LC_15_27_2 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_13_LC_15_27_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_13_LC_15_27_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_13_LC_15_27_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64230),
            .lcout(\pid_front.error_d_regZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94374),
            .ce(N__93370),
            .sr(N__93005));
    defparam \pid_front.error_p_reg_esr_13_LC_15_27_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_13_LC_15_27_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_13_LC_15_27_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_13_LC_15_27_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64210),
            .lcout(\pid_front.error_p_regZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94374),
            .ce(N__93370),
            .sr(N__93005));
    defparam \pid_front.error_d_reg_prev_esr_RNI8QE61_0_20_LC_15_27_4 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNI8QE61_0_20_LC_15_27_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNI8QE61_0_20_LC_15_27_4 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNI8QE61_0_20_LC_15_27_4  (
            .in0(N__66662),
            .in1(N__67113),
            .in2(_gnd_net_),
            .in3(N__91856),
            .lcout(\pid_front.error_d_reg_prev_esr_RNI8QE61_0Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNI8QE61_20_LC_15_27_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNI8QE61_20_LC_15_27_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNI8QE61_20_LC_15_27_6 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNI8QE61_20_LC_15_27_6  (
            .in0(N__66661),
            .in1(N__67114),
            .in2(_gnd_net_),
            .in3(N__91857),
            .lcout(\pid_front.error_d_reg_prev_esr_RNI8QE61Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_20_LC_15_27_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_20_LC_15_27_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_20_LC_15_27_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_20_LC_15_27_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64150),
            .lcout(\pid_front.error_p_regZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94374),
            .ce(N__93370),
            .sr(N__93005));
    defparam \pid_front.error_d_reg_fast_esr_RNISQ181_12_LC_15_28_0 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_fast_esr_RNISQ181_12_LC_15_28_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_fast_esr_RNISQ181_12_LC_15_28_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \pid_front.error_d_reg_fast_esr_RNISQ181_12_LC_15_28_0  (
            .in0(N__64347),
            .in1(N__67635),
            .in2(N__71980),
            .in3(N__67685),
            .lcout(),
            .ltout(\pid_front.error_d_reg_fast_esr_RNISQ181Z0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_fast_esr_RNIKO3P2_12_LC_15_28_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_fast_esr_RNIKO3P2_12_LC_15_28_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_fast_esr_RNIKO3P2_12_LC_15_28_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \pid_front.error_d_reg_prev_fast_esr_RNIKO3P2_12_LC_15_28_1  (
            .in0(N__67432),
            .in1(_gnd_net_),
            .in2(N__64129),
            .in3(N__64126),
            .lcout(),
            .ltout(\pid_front.g0_3_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI7AR55_12_LC_15_28_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI7AR55_12_LC_15_28_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI7AR55_12_LC_15_28_2 .LUT_INIT=16'b1110000110000111;
    LogicCell40 \pid_front.error_p_reg_esr_RNI7AR55_12_LC_15_28_2  (
            .in0(N__64120),
            .in1(N__67168),
            .in2(N__64108),
            .in3(N__71904),
            .lcout(),
            .ltout(\pid_front.g1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIOH2JD_12_LC_15_28_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIOH2JD_12_LC_15_28_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIOH2JD_12_LC_15_28_3 .LUT_INIT=16'b1000000011101010;
    LogicCell40 \pid_front.error_p_reg_esr_RNIOH2JD_12_LC_15_28_3  (
            .in0(N__69961),
            .in1(N__64404),
            .in2(N__64366),
            .in3(N__67516),
            .lcout(\pid_front.error_p_reg_esr_RNIOH2JDZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_13_LC_15_28_5 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_13_LC_15_28_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_13_LC_15_28_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_13_LC_15_28_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64348),
            .lcout(\pid_front.error_d_reg_prevZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94382),
            .ce(N__71824),
            .sr(N__71714));
    defparam \pid_front.error_d_reg_esr_RNIETB61_0_13_LC_15_28_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_RNIETB61_0_13_LC_15_28_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_esr_RNIETB61_0_13_LC_15_28_6 .LUT_INIT=16'b1000100011101110;
    LogicCell40 \pid_front.error_d_reg_esr_RNIETB61_0_13_LC_15_28_6  (
            .in0(N__64346),
            .in1(N__67684),
            .in2(_gnd_net_),
            .in3(N__67634),
            .lcout(),
            .ltout(\pid_front.N_2401_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIVTNC2_14_LC_15_28_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIVTNC2_14_LC_15_28_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIVTNC2_14_LC_15_28_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \pid_front.error_p_reg_esr_RNIVTNC2_14_LC_15_28_7  (
            .in0(N__67579),
            .in1(N__67557),
            .in2(N__64321),
            .in3(N__94536),
            .lcout(\pid_front.g0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un11lto30_i_a2_0_c_RNO_LC_16_3_5 .C_ON=1'b0;
    defparam \pid_side.un11lto30_i_a2_0_c_RNO_LC_16_3_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.un11lto30_i_a2_0_c_RNO_LC_16_3_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_side.un11lto30_i_a2_0_c_RNO_LC_16_3_5  (
            .in0(N__64245),
            .in1(N__64266),
            .in2(N__64658),
            .in3(N__64289),
            .lcout(\pid_side.source_pid10lt4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_16_4_0 .C_ON=1'b1;
    defparam \pid_side.un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_16_4_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_16_4_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_side.un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_16_4_0  (
            .in0(_gnd_net_),
            .in1(N__89874),
            .in2(N__89878),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_16_4_0_),
            .carryout(\pid_side.un1_pid_prereg_0_cry_0_c_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_0_LC_16_4_1 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_0_LC_16_4_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_0_LC_16_4_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_0_LC_16_4_1  (
            .in0(_gnd_net_),
            .in1(N__72679),
            .in2(N__72702),
            .in3(N__64276),
            .lcout(\pid_side.pid_preregZ0Z_0 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_0_c_THRU_CO ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_0 ),
            .clk(N__94100),
            .ce(N__65074),
            .sr(N__86462));
    defparam \pid_side.pid_prereg_esr_1_LC_16_4_2 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_1_LC_16_4_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_1_LC_16_4_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_1_LC_16_4_2  (
            .in0(_gnd_net_),
            .in1(N__72307),
            .in2(N__72336),
            .in3(N__64255),
            .lcout(\pid_side.pid_preregZ0Z_1 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_0 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_1 ),
            .clk(N__94100),
            .ce(N__65074),
            .sr(N__86462));
    defparam \pid_side.pid_prereg_esr_2_LC_16_4_3 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_2_LC_16_4_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_2_LC_16_4_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_2_LC_16_4_3  (
            .in0(_gnd_net_),
            .in1(N__76414),
            .in2(N__76449),
            .in3(N__64234),
            .lcout(\pid_side.pid_preregZ0Z_2 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_1 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_2 ),
            .clk(N__94100),
            .ce(N__65074),
            .sr(N__86462));
    defparam \pid_side.pid_prereg_esr_3_LC_16_4_4 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_3_LC_16_4_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_3_LC_16_4_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_3_LC_16_4_4  (
            .in0(_gnd_net_),
            .in1(N__79015),
            .in2(N__78988),
            .in3(N__64639),
            .lcout(\pid_side.pid_preregZ0Z_3 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_2 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_3 ),
            .clk(N__94100),
            .ce(N__65074),
            .sr(N__86462));
    defparam \pid_side.pid_prereg_esr_4_LC_16_4_5 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_4_LC_16_4_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_4_LC_16_4_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_4_LC_16_4_5  (
            .in0(_gnd_net_),
            .in1(N__76333),
            .in2(N__78937),
            .in3(N__64603),
            .lcout(\pid_side.pid_preregZ0Z_4 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_3 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_4 ),
            .clk(N__94100),
            .ce(N__65074),
            .sr(N__86462));
    defparam \pid_side.pid_prereg_esr_5_LC_16_4_6 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_5_LC_16_4_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_5_LC_16_4_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_5_LC_16_4_6  (
            .in0(_gnd_net_),
            .in1(N__76027),
            .in2(N__76387),
            .in3(N__64567),
            .lcout(\pid_side.pid_preregZ0Z_5 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_4 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_5 ),
            .clk(N__94100),
            .ce(N__65074),
            .sr(N__86462));
    defparam \pid_side.pid_prereg_esr_6_LC_16_4_7 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_6_LC_16_4_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_6_LC_16_4_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_6_LC_16_4_7  (
            .in0(_gnd_net_),
            .in1(N__67858),
            .in2(N__76093),
            .in3(N__64528),
            .lcout(\pid_side.pid_preregZ0Z_6 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_5 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_6 ),
            .clk(N__94100),
            .ce(N__65074),
            .sr(N__86462));
    defparam \pid_side.pid_prereg_esr_7_LC_16_5_0 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_7_LC_16_5_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_7_LC_16_5_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_7_LC_16_5_0  (
            .in0(_gnd_net_),
            .in1(N__72253),
            .in2(N__67819),
            .in3(N__64489),
            .lcout(\pid_side.pid_preregZ0Z_7 ),
            .ltout(),
            .carryin(bfn_16_5_0_),
            .carryout(\pid_side.un1_pid_prereg_0_cry_7 ),
            .clk(N__94106),
            .ce(N__65075),
            .sr(N__86457));
    defparam \pid_side.pid_prereg_esr_8_LC_16_5_1 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_8_LC_16_5_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_8_LC_16_5_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_8_LC_16_5_1  (
            .in0(_gnd_net_),
            .in1(N__72217),
            .in2(N__72163),
            .in3(N__64459),
            .lcout(\pid_side.pid_preregZ0Z_8 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_7 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_8 ),
            .clk(N__94106),
            .ce(N__65075),
            .sr(N__86457));
    defparam \pid_side.pid_prereg_esr_9_LC_16_5_2 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_9_LC_16_5_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_9_LC_16_5_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_9_LC_16_5_2  (
            .in0(_gnd_net_),
            .in1(N__72421),
            .in2(N__72441),
            .in3(N__64435),
            .lcout(\pid_side.pid_preregZ0Z_9 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_8 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_9 ),
            .clk(N__94106),
            .ce(N__65075),
            .sr(N__86457));
    defparam \pid_side.pid_prereg_esr_10_LC_16_5_3 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_10_LC_16_5_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_10_LC_16_5_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_10_LC_16_5_3  (
            .in0(_gnd_net_),
            .in1(N__72787),
            .in2(N__72814),
            .in3(N__64408),
            .lcout(\pid_side.pid_preregZ0Z_10 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_9 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_10 ),
            .clk(N__94106),
            .ce(N__65075),
            .sr(N__86457));
    defparam \pid_side.pid_prereg_esr_11_LC_16_5_4 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_11_LC_16_5_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_11_LC_16_5_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_11_LC_16_5_4  (
            .in0(_gnd_net_),
            .in1(N__73152),
            .in2(N__73114),
            .in3(N__64846),
            .lcout(\pid_side.pid_preregZ0Z_11 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_10 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_11 ),
            .clk(N__94106),
            .ce(N__65075),
            .sr(N__86457));
    defparam \pid_side.pid_prereg_esr_12_LC_16_5_5 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_12_LC_16_5_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_12_LC_16_5_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_12_LC_16_5_5  (
            .in0(_gnd_net_),
            .in1(N__68398),
            .in2(N__72505),
            .in3(N__64807),
            .lcout(\pid_side.pid_preregZ0Z_12 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_11 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_12 ),
            .clk(N__94106),
            .ce(N__65075),
            .sr(N__86457));
    defparam \pid_side.pid_prereg_esr_13_LC_16_5_6 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_13_LC_16_5_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_13_LC_16_5_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_13_LC_16_5_6  (
            .in0(_gnd_net_),
            .in1(N__68650),
            .in2(N__68611),
            .in3(N__64771),
            .lcout(\pid_side.pid_preregZ0Z_13 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_12 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_13 ),
            .clk(N__94106),
            .ce(N__65075),
            .sr(N__86457));
    defparam \pid_side.un1_pid_prereg_0_cry_13_THRU_LUT4_0_LC_16_5_7 .C_ON=1'b1;
    defparam \pid_side.un1_pid_prereg_0_cry_13_THRU_LUT4_0_LC_16_5_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_pid_prereg_0_cry_13_THRU_LUT4_0_LC_16_5_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.un1_pid_prereg_0_cry_13_THRU_LUT4_0_LC_16_5_7  (
            .in0(_gnd_net_),
            .in1(N__65343),
            .in2(_gnd_net_),
            .in3(N__64759),
            .lcout(\pid_side.un1_pid_prereg_0_cry_13_THRU_CO ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_13 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_15_LC_16_6_0 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_15_LC_16_6_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_15_LC_16_6_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_15_LC_16_6_0  (
            .in0(_gnd_net_),
            .in1(N__68047),
            .in2(N__76486),
            .in3(N__64729),
            .lcout(\pid_side.pid_preregZ0Z_15 ),
            .ltout(),
            .carryin(bfn_16_6_0_),
            .carryout(\pid_side.un1_pid_prereg_0_cry_15 ),
            .clk(N__94113),
            .ce(N__65076),
            .sr(N__86452));
    defparam \pid_side.pid_prereg_esr_16_LC_16_6_1 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_16_LC_16_6_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_16_LC_16_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_16_LC_16_6_1  (
            .in0(_gnd_net_),
            .in1(N__68011),
            .in2(N__64726),
            .in3(N__64711),
            .lcout(\pid_side.pid_preregZ0Z_16 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_15 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_16 ),
            .clk(N__94113),
            .ce(N__65076),
            .sr(N__86452));
    defparam \pid_side.pid_prereg_esr_17_LC_16_6_2 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_17_LC_16_6_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_17_LC_16_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_17_LC_16_6_2  (
            .in0(_gnd_net_),
            .in1(N__64708),
            .in2(N__64702),
            .in3(N__64687),
            .lcout(\pid_side.pid_preregZ0Z_17 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_16 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_17 ),
            .clk(N__94113),
            .ce(N__65076),
            .sr(N__86452));
    defparam \pid_side.pid_prereg_esr_18_LC_16_6_3 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_18_LC_16_6_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_18_LC_16_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_18_LC_16_6_3  (
            .in0(_gnd_net_),
            .in1(N__64684),
            .in2(N__64678),
            .in3(N__64663),
            .lcout(\pid_side.pid_preregZ0Z_18 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_17 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_18 ),
            .clk(N__94113),
            .ce(N__65076),
            .sr(N__86452));
    defparam \pid_side.pid_prereg_esr_19_LC_16_6_4 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_19_LC_16_6_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_19_LC_16_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_19_LC_16_6_4  (
            .in0(_gnd_net_),
            .in1(N__68185),
            .in2(N__65005),
            .in3(N__64987),
            .lcout(\pid_side.pid_preregZ0Z_19 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_18 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_19 ),
            .clk(N__94113),
            .ce(N__65076),
            .sr(N__86452));
    defparam \pid_side.pid_prereg_esr_20_LC_16_6_5 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_20_LC_16_6_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_20_LC_16_6_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_20_LC_16_6_5  (
            .in0(_gnd_net_),
            .in1(N__68452),
            .in2(N__65386),
            .in3(N__64978),
            .lcout(\pid_side.pid_preregZ0Z_20 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_19 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_20 ),
            .clk(N__94113),
            .ce(N__65076),
            .sr(N__86452));
    defparam \pid_side.pid_prereg_esr_21_LC_16_6_6 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_21_LC_16_6_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_21_LC_16_6_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_21_LC_16_6_6  (
            .in0(_gnd_net_),
            .in1(N__68005),
            .in2(N__65251),
            .in3(N__64969),
            .lcout(\pid_side.pid_preregZ0Z_21 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_20 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_21 ),
            .clk(N__94113),
            .ce(N__65076),
            .sr(N__86452));
    defparam \pid_side.pid_prereg_esr_22_LC_16_6_7 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_22_LC_16_6_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_22_LC_16_6_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_22_LC_16_6_7  (
            .in0(_gnd_net_),
            .in1(N__67903),
            .in2(N__65026),
            .in3(N__64960),
            .lcout(\pid_side.pid_preregZ0Z_22 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_21 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_22 ),
            .clk(N__94113),
            .ce(N__65076),
            .sr(N__86452));
    defparam \pid_side.pid_prereg_esr_23_LC_16_7_0 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_23_LC_16_7_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_23_LC_16_7_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_23_LC_16_7_0  (
            .in0(_gnd_net_),
            .in1(N__67999),
            .in2(N__65041),
            .in3(N__64945),
            .lcout(\pid_side.pid_preregZ0Z_23 ),
            .ltout(),
            .carryin(bfn_16_7_0_),
            .carryout(\pid_side.un1_pid_prereg_0_cry_23 ),
            .clk(N__94120),
            .ce(N__65077),
            .sr(N__86449));
    defparam \pid_side.pid_prereg_esr_24_LC_16_7_1 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_24_LC_16_7_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_24_LC_16_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_24_LC_16_7_1  (
            .in0(_gnd_net_),
            .in1(N__65314),
            .in2(N__68263),
            .in3(N__64933),
            .lcout(\pid_side.pid_preregZ0Z_24 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_23 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_24 ),
            .clk(N__94120),
            .ce(N__65077),
            .sr(N__86449));
    defparam \pid_side.pid_prereg_esr_25_LC_16_7_2 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_25_LC_16_7_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_25_LC_16_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_25_LC_16_7_2  (
            .in0(_gnd_net_),
            .in1(N__68125),
            .in2(N__65014),
            .in3(N__64921),
            .lcout(\pid_side.pid_preregZ0Z_25 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_24 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_25 ),
            .clk(N__94120),
            .ce(N__65077),
            .sr(N__86449));
    defparam \pid_side.pid_prereg_esr_26_LC_16_7_3 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_26_LC_16_7_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_26_LC_16_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_26_LC_16_7_3  (
            .in0(_gnd_net_),
            .in1(N__64918),
            .in2(N__68425),
            .in3(N__64897),
            .lcout(\pid_side.pid_preregZ0Z_26 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_25 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_26 ),
            .clk(N__94120),
            .ce(N__65077),
            .sr(N__86449));
    defparam \pid_side.pid_prereg_esr_27_LC_16_7_4 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_27_LC_16_7_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_27_LC_16_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_27_LC_16_7_4  (
            .in0(_gnd_net_),
            .in1(N__64894),
            .in2(N__65212),
            .in3(N__65185),
            .lcout(\pid_side.pid_preregZ0Z_27 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_26 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_27 ),
            .clk(N__94120),
            .ce(N__65077),
            .sr(N__86449));
    defparam \pid_side.pid_prereg_esr_28_LC_16_7_5 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_28_LC_16_7_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_28_LC_16_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_28_LC_16_7_5  (
            .in0(_gnd_net_),
            .in1(N__68305),
            .in2(N__65182),
            .in3(N__65155),
            .lcout(\pid_side.pid_preregZ0Z_28 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_27 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_28 ),
            .clk(N__94120),
            .ce(N__65077),
            .sr(N__86449));
    defparam \pid_side.pid_prereg_esr_29_LC_16_7_6 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_29_LC_16_7_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_29_LC_16_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_29_LC_16_7_6  (
            .in0(_gnd_net_),
            .in1(N__68299),
            .in2(N__72715),
            .in3(N__65140),
            .lcout(\pid_side.pid_preregZ0Z_29 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_28 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_29 ),
            .clk(N__94120),
            .ce(N__65077),
            .sr(N__86449));
    defparam \pid_side.pid_prereg_esr_30_LC_16_7_7 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_30_LC_16_7_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_30_LC_16_7_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_side.pid_prereg_esr_30_LC_16_7_7  (
            .in0(_gnd_net_),
            .in1(N__67897),
            .in2(_gnd_net_),
            .in3(N__65137),
            .lcout(\pid_side.pid_preregZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94120),
            .ce(N__65077),
            .sr(N__86449));
    defparam \pid_side.error_d_reg_prev_esr_RNIC7HE7_21_LC_16_8_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIC7HE7_21_LC_16_8_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIC7HE7_21_LC_16_8_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIC7HE7_21_LC_16_8_0  (
            .in0(N__67918),
            .in1(N__68292),
            .in2(N__67960),
            .in3(N__68279),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIC7HE7Z0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIEE3E2_0_20_LC_16_8_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIEE3E2_0_20_LC_16_8_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIEE3E2_0_20_LC_16_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIEE3E2_0_20_LC_16_8_1  (
            .in0(N__65287),
            .in1(N__67483),
            .in2(_gnd_net_),
            .in3(N__65304),
            .lcout(\pid_side.un1_pid_prereg_0_11 ),
            .ltout(\pid_side.un1_pid_prereg_0_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIPUAR4_19_LC_16_8_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIPUAR4_19_LC_16_8_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIPUAR4_19_LC_16_8_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIPUAR4_19_LC_16_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__65029),
            .in3(N__67945),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIPUAR4Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIBG7D2_19_LC_16_8_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIBG7D2_19_LC_16_8_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIBG7D2_19_LC_16_8_3 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIBG7D2_19_LC_16_8_3  (
            .in0(N__67509),
            .in1(N__76317),
            .in2(_gnd_net_),
            .in3(N__65277),
            .lcout(\pid_side.un1_pid_prereg_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIE21B3_21_LC_16_8_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIE21B3_21_LC_16_8_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIE21B3_21_LC_16_8_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIE21B3_21_LC_16_8_4  (
            .in0(_gnd_net_),
            .in1(N__68143),
            .in2(_gnd_net_),
            .in3(N__68154),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIE21B3Z0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIMVFL1_0_21_LC_16_8_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIMVFL1_0_21_LC_16_8_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIMVFL1_0_21_LC_16_8_5 .LUT_INIT=16'b0001100011100111;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIMVFL1_0_21_LC_16_8_5  (
            .in0(N__91374),
            .in1(N__91646),
            .in2(N__72930),
            .in3(N__68253),
            .lcout(\pid_side.un1_pid_prereg_0_15 ),
            .ltout(\pid_side.un1_pid_prereg_0_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIASUA3_21_LC_16_8_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIASUA3_21_LC_16_8_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIASUA3_21_LC_16_8_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIASUA3_21_LC_16_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__65317),
            .in3(N__68280),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIASUA3Z0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIEE3E2_20_LC_16_8_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIEE3E2_20_LC_16_8_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIEE3E2_20_LC_16_8_7 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIEE3E2_20_LC_16_8_7  (
            .in0(N__65286),
            .in1(N__67482),
            .in2(_gnd_net_),
            .in3(N__65303),
            .lcout(\pid_side.un1_pid_prereg_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIUMLO_21_LC_16_9_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIUMLO_21_LC_16_9_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIUMLO_21_LC_16_9_0 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIUMLO_21_LC_16_9_0  (
            .in0(N__72928),
            .in1(N__91370),
            .in2(_gnd_net_),
            .in3(N__91625),
            .lcout(\pid_side.un1_pid_prereg_370_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIBG7D2_0_19_LC_16_9_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIBG7D2_0_19_LC_16_9_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIBG7D2_0_19_LC_16_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIBG7D2_0_19_LC_16_9_1  (
            .in0(N__67510),
            .in1(N__76318),
            .in2(_gnd_net_),
            .in3(N__65273),
            .lcout(\pid_side.un1_pid_prereg_0_9 ),
            .ltout(\pid_side.un1_pid_prereg_0_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIIOAQ4_18_LC_16_9_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIIOAQ4_18_LC_16_9_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIIOAQ4_18_LC_16_9_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIIOAQ4_18_LC_16_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__65254),
            .in3(N__68063),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIIOAQ4Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI783D2_18_LC_16_9_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI783D2_18_LC_16_9_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI783D2_18_LC_16_9_3 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI783D2_18_LC_16_9_3  (
            .in0(N__76296),
            .in1(N__82440),
            .in2(_gnd_net_),
            .in3(N__65402),
            .lcout(\pid_side.un1_pid_prereg_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIVU1D2_17_LC_16_9_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIVU1D2_17_LC_16_9_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIVU1D2_17_LC_16_9_4 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIVU1D2_17_LC_16_9_4  (
            .in0(N__87849),
            .in1(N__67770),
            .in2(_gnd_net_),
            .in3(N__65228),
            .lcout(\pid_side.un1_pid_prereg_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIKSEL1_21_LC_16_9_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIKSEL1_21_LC_16_9_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIKSEL1_21_LC_16_9_5 .LUT_INIT=16'b1111101100100000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIKSEL1_21_LC_16_9_5  (
            .in0(N__91626),
            .in1(N__72929),
            .in2(N__91384),
            .in3(N__67979),
            .lcout(\pid_side.un1_pid_prereg_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI783D2_0_18_LC_16_9_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI783D2_0_18_LC_16_9_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI783D2_0_18_LC_16_9_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI783D2_0_18_LC_16_9_6  (
            .in0(N__65403),
            .in1(_gnd_net_),
            .in2(N__82444),
            .in3(N__76297),
            .lcout(\pid_side.un1_pid_prereg_0_7 ),
            .ltout(\pid_side.un1_pid_prereg_0_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI675Q4_17_LC_16_9_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI675Q4_17_LC_16_9_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI675Q4_17_LC_16_9_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI675Q4_17_LC_16_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__65389),
            .in3(N__68084),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI675Q4Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIMERG_2_12_LC_16_10_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIMERG_2_12_LC_16_10_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIMERG_2_12_LC_16_10_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIMERG_2_12_LC_16_10_0  (
            .in0(_gnd_net_),
            .in1(N__79445),
            .in2(_gnd_net_),
            .in3(N__91244),
            .lcout(),
            .ltout(\pid_side.N_3_i_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIR3TQ1_12_LC_16_10_1 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIR3TQ1_12_LC_16_10_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIR3TQ1_12_LC_16_10_1 .LUT_INIT=16'b0000010100010111;
    LogicCell40 \pid_side.error_p_reg_esr_RNIR3TQ1_12_LC_16_10_1  (
            .in0(N__90982),
            .in1(N__82405),
            .in2(N__65371),
            .in3(N__68563),
            .lcout(),
            .ltout(\pid_side.N_3_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIQTGL4_12_LC_16_10_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIQTGL4_12_LC_16_10_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIQTGL4_12_LC_16_10_2 .LUT_INIT=16'b0010101111010100;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIQTGL4_12_LC_16_10_2  (
            .in0(N__65326),
            .in1(N__65368),
            .in2(N__65356),
            .in3(N__76462),
            .lcout(),
            .ltout(\pid_side.error_d_reg_prev_esr_RNIQTGL4Z0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIRPTT9_12_LC_16_10_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIRPTT9_12_LC_16_10_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIRPTT9_12_LC_16_10_3 .LUT_INIT=16'b1001011001011010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIRPTT9_12_LC_16_10_3  (
            .in0(N__76535),
            .in1(N__76512),
            .in2(N__65353),
            .in3(N__68538),
            .lcout(\pid_side.un1_pid_prereg_0_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIMERG_12_LC_16_10_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIMERG_12_LC_16_10_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIMERG_12_LC_16_10_4 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIMERG_12_LC_16_10_4  (
            .in0(_gnd_net_),
            .in1(N__79446),
            .in2(_gnd_net_),
            .in3(N__91245),
            .lcout(\pid_side.N_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_12_LC_16_10_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_12_LC_16_10_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_12_LC_16_10_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_12_LC_16_10_5  (
            .in0(N__91246),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94146),
            .ce(N__88107),
            .sr(N__87940));
    defparam \pid_side.error_d_reg_prev_esr_RNI0TN9_11_LC_16_10_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI0TN9_11_LC_16_10_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI0TN9_11_LC_16_10_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI0TN9_11_LC_16_10_6  (
            .in0(_gnd_net_),
            .in1(N__91026),
            .in2(_gnd_net_),
            .in3(N__82372),
            .lcout(\pid_side.un1_pid_prereg_79 ),
            .ltout(\pid_side.un1_pid_prereg_79_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIL0VP1_12_LC_16_10_7 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIL0VP1_12_LC_16_10_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIL0VP1_12_LC_16_10_7 .LUT_INIT=16'b0110011001101001;
    LogicCell40 \pid_side.error_p_reg_esr_RNIL0VP1_12_LC_16_10_7  (
            .in0(N__69658),
            .in1(N__90973),
            .in2(N__65320),
            .in3(N__82404),
            .lcout(\pid_side.error_p_reg_esr_RNIL0VP1Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_0_0_c_RNI6CR94_LC_16_11_0 .C_ON=1'b0;
    defparam \pid_side.error_cry_0_0_c_RNI6CR94_LC_16_11_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_0_c_RNI6CR94_LC_16_11_0 .LUT_INIT=16'b0101010100010101;
    LogicCell40 \pid_side.error_cry_0_0_c_RNI6CR94_LC_16_11_0  (
            .in0(N__65965),
            .in1(N__81332),
            .in2(N__65428),
            .in3(N__89373),
            .lcout(),
            .ltout(\pid_side.m13_2_03_4_i_0_o2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_3_0_c_RNIK741H_LC_16_11_1 .C_ON=1'b0;
    defparam \pid_side.error_cry_3_0_c_RNIK741H_LC_16_11_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_3_0_c_RNIK741H_LC_16_11_1 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \pid_side.error_cry_3_0_c_RNIK741H_LC_16_11_1  (
            .in0(N__65868),
            .in1(_gnd_net_),
            .in2(N__65515),
            .in3(N__65974),
            .lcout(\pid_side.m13_2_03_4_i_3 ),
            .ltout(\pid_side.m13_2_03_4_i_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_9_LC_16_11_2 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_9_LC_16_11_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_9_LC_16_11_2 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \pid_side.error_i_reg_9_LC_16_11_2  (
            .in0(N__83267),
            .in1(N__65483),
            .in2(N__65506),
            .in3(N__65499),
            .lcout(\pid_side.error_i_regZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94158),
            .ce(),
            .sr(N__86437));
    defparam \pid_side.error_i_reg_7_LC_16_11_3 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_7_LC_16_11_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_7_LC_16_11_3 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \pid_side.error_i_reg_7_LC_16_11_3  (
            .in0(N__65482),
            .in1(N__83268),
            .in2(N__65446),
            .in3(N__73234),
            .lcout(\pid_side.error_i_regZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94158),
            .ce(),
            .sr(N__86437));
    defparam \pid_side.error_i_reg_esr_RNO_1_11_LC_16_11_4 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_1_11_LC_16_11_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_1_11_LC_16_11_4 .LUT_INIT=16'b1100110011101100;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_1_11_LC_16_11_4  (
            .in0(N__85738),
            .in1(N__68677),
            .in2(N__83311),
            .in3(N__73428),
            .lcout(\pid_side.m78_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_4_c_RNIEP6K1_LC_16_11_5 .C_ON=1'b0;
    defparam \pid_side.error_cry_4_c_RNIEP6K1_LC_16_11_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_4_c_RNIEP6K1_LC_16_11_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \pid_side.error_cry_4_c_RNIEP6K1_LC_16_11_5  (
            .in0(N__90427),
            .in1(N__80489),
            .in2(_gnd_net_),
            .in3(N__80417),
            .lcout(\pid_side.N_163 ),
            .ltout(\pid_side.N_163_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_0_c_RNIR8943_LC_16_11_6 .C_ON=1'b0;
    defparam \pid_side.error_cry_0_c_RNIR8943_LC_16_11_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_c_RNIR8943_LC_16_11_6 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \pid_side.error_cry_0_c_RNIR8943_LC_16_11_6  (
            .in0(_gnd_net_),
            .in1(N__89372),
            .in2(N__65419),
            .in3(N__82885),
            .lcout(\pid_side.N_186 ),
            .ltout(\pid_side.N_186_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_3_27_LC_16_11_7 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_3_27_LC_16_11_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_3_27_LC_16_11_7 .LUT_INIT=16'b0010101000000000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_3_27_LC_16_11_7  (
            .in0(N__87035),
            .in1(N__85737),
            .in2(N__65416),
            .in3(N__84322),
            .lcout(\pid_side.error_i_reg_9_sn_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_3_11_LC_16_12_0 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_3_11_LC_16_12_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_3_11_LC_16_12_0 .LUT_INIT=16'b0000111000000100;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_3_11_LC_16_12_0  (
            .in0(N__82640),
            .in1(N__80699),
            .in2(N__73675),
            .in3(N__78325),
            .lcout(\pid_front.N_394 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_0_26_LC_16_12_1 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_26_LC_16_12_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_26_LC_16_12_1 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_26_LC_16_12_1  (
            .in0(N__80700),
            .in1(N__86970),
            .in2(_gnd_net_),
            .in3(N__84321),
            .lcout(\pid_front.error_i_reg_9_rn_1_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_ki_0_rep2_esr_LC_16_12_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_0_rep2_esr_LC_16_12_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_0_rep2_esr_LC_16_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_0_rep2_esr_LC_16_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88305),
            .lcout(xy_ki_0_rep2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94169),
            .ce(N__83894),
            .sr(N__86428));
    defparam \pid_side.error_cry_3_c_RNIMCQD2_LC_16_12_3 .C_ON=1'b0;
    defparam \pid_side.error_cry_3_c_RNIMCQD2_LC_16_12_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_3_c_RNIMCQD2_LC_16_12_3 .LUT_INIT=16'b0010000001110000;
    LogicCell40 \pid_side.error_cry_3_c_RNIMCQD2_LC_16_12_3  (
            .in0(N__82635),
            .in1(N__77231),
            .in2(N__90545),
            .in3(N__80310),
            .lcout(\pid_side.N_27_0_i_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_ki_1_rep1_esr_LC_16_12_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_1_rep1_esr_LC_16_12_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_1_rep1_esr_LC_16_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_1_rep1_esr_LC_16_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85528),
            .lcout(xy_ki_1_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94169),
            .ce(N__83894),
            .sr(N__86428));
    defparam \pid_front.m10_2_03_3_i_0_a2_1_0_LC_16_12_5 .C_ON=1'b0;
    defparam \pid_front.m10_2_03_3_i_0_a2_1_0_LC_16_12_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.m10_2_03_3_i_0_a2_1_0_LC_16_12_5 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \pid_front.m10_2_03_3_i_0_a2_1_0_LC_16_12_5  (
            .in0(N__90498),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__90343),
            .lcout(pid_side_m10_2_03_3_i_0_a2_1_0),
            .ltout(pid_side_m10_2_03_3_i_0_a2_1_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_5_c_RNIA9135_LC_16_12_6 .C_ON=1'b0;
    defparam \pid_side.error_cry_5_c_RNIA9135_LC_16_12_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_5_c_RNIA9135_LC_16_12_6 .LUT_INIT=16'b0000101110111011;
    LogicCell40 \pid_side.error_cry_5_c_RNIA9135_LC_16_12_6  (
            .in0(N__81404),
            .in1(N__77605),
            .in2(N__65980),
            .in3(N__80056),
            .lcout(),
            .ltout(\pid_side.m13_2_03_4_i_0_o2_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_3_0_c_RNIER8NC_LC_16_12_7 .C_ON=1'b0;
    defparam \pid_side.error_cry_3_0_c_RNIER8NC_LC_16_12_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_3_0_c_RNIER8NC_LC_16_12_7 .LUT_INIT=16'b1111111110001111;
    LogicCell40 \pid_side.error_cry_3_0_c_RNIER8NC_LC_16_12_7  (
            .in0(N__83496),
            .in1(N__79738),
            .in2(N__65977),
            .in3(N__68755),
            .lcout(\pid_side.error_cry_3_0_c_RNIER8NCZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_6_c_RNINJQB2_LC_16_13_0 .C_ON=1'b0;
    defparam \pid_side.error_cry_6_c_RNINJQB2_LC_16_13_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_6_c_RNINJQB2_LC_16_13_0 .LUT_INIT=16'b1000110010011100;
    LogicCell40 \pid_side.error_cry_6_c_RNINJQB2_LC_16_13_0  (
            .in0(N__90211),
            .in1(N__66079),
            .in2(N__90408),
            .in3(N__87554),
            .lcout(),
            .ltout(\pid_side.m18_2_03_4_o3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_6_c_RNII55P7_LC_16_13_1 .C_ON=1'b0;
    defparam \pid_side.error_cry_6_c_RNII55P7_LC_16_13_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_6_c_RNII55P7_LC_16_13_1 .LUT_INIT=16'b1110110011101101;
    LogicCell40 \pid_side.error_cry_6_c_RNII55P7_LC_16_13_1  (
            .in0(N__89842),
            .in1(N__69526),
            .in2(N__65968),
            .in3(N__76647),
            .lcout(\pid_side.N_263 ),
            .ltout(\pid_side.N_263_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_1_14_LC_16_13_2 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_1_14_LC_16_13_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_1_14_LC_16_13_2 .LUT_INIT=16'b0000000000010011;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_1_14_LC_16_13_2  (
            .in0(N__87376),
            .in1(N__73219),
            .in2(N__66088),
            .in3(N__76762),
            .lcout(\pid_side.error_i_reg_esr_RNO_1Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_2_c_RNIKQQ01_LC_16_13_3 .C_ON=1'b0;
    defparam \pid_side.error_cry_2_c_RNIKQQ01_LC_16_13_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_2_c_RNIKQQ01_LC_16_13_3 .LUT_INIT=16'b0001010110010101;
    LogicCell40 \pid_side.error_cry_2_c_RNIKQQ01_LC_16_13_3  (
            .in0(N__82636),
            .in1(N__90207),
            .in2(N__90347),
            .in3(N__80863),
            .lcout(\pid_side.m18_2_03_4_o3_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_4_c_RNIMV991_0_LC_16_13_4 .C_ON=1'b0;
    defparam \pid_front.error_cry_4_c_RNIMV991_0_LC_16_13_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_4_c_RNIMV991_0_LC_16_13_4 .LUT_INIT=16'b0000111000000010;
    LogicCell40 \pid_front.error_cry_4_c_RNIMV991_0_LC_16_13_4  (
            .in0(N__73794),
            .in1(N__90302),
            .in2(N__90239),
            .in3(N__77972),
            .lcout(\pid_front.N_629 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_2_12_LC_16_13_5 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_2_12_LC_16_13_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_2_12_LC_16_13_5 .LUT_INIT=16'b1010001000000010;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_2_12_LC_16_13_5  (
            .in0(N__89109),
            .in1(N__66031),
            .in2(N__89850),
            .in3(N__80512),
            .lcout(),
            .ltout(\pid_side.m16_2_03_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_1_12_LC_16_13_6 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_1_12_LC_16_13_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_1_12_LC_16_13_6 .LUT_INIT=16'b1111010111110100;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_1_12_LC_16_13_6  (
            .in0(N__87375),
            .in1(N__68745),
            .in2(N__66016),
            .in3(N__66013),
            .lcout(\pid_side.m16_2_03_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_ki_2_rep1_esr_LC_16_13_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_2_rep1_esr_LC_16_13_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_2_rep1_esr_LC_16_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_2_rep1_esr_LC_16_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__92513),
            .lcout(xy_ki_2_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94184),
            .ce(N__83889),
            .sr(N__86418));
    defparam \pid_front.m28_2_03_0_a2_1_1_LC_16_14_0 .C_ON=1'b0;
    defparam \pid_front.m28_2_03_0_a2_1_1_LC_16_14_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.m28_2_03_0_a2_1_1_LC_16_14_0 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \pid_front.m28_2_03_0_a2_1_1_LC_16_14_0  (
            .in0(N__83084),
            .in1(N__82259),
            .in2(N__79650),
            .in3(N__80135),
            .lcout(pid_front_N_474_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_ki_fast_esr_1_LC_16_14_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_fast_esr_1_LC_16_14_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_fast_esr_1_LC_16_14_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_fast_esr_1_LC_16_14_1  (
            .in0(N__85513),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(xy_ki_fast_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94196),
            .ce(N__83888),
            .sr(N__86407));
    defparam \pid_side.N_45_i_i_a2_2_LC_16_14_2 .C_ON=1'b0;
    defparam \pid_side.N_45_i_i_a2_2_LC_16_14_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.N_45_i_i_a2_2_LC_16_14_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \pid_side.N_45_i_i_a2_2_LC_16_14_2  (
            .in0(N__83083),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82258),
            .lcout(pid_side_N_492),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_2_c_RNI72F32_LC_16_14_3 .C_ON=1'b0;
    defparam \pid_side.error_cry_2_c_RNI72F32_LC_16_14_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_2_c_RNI72F32_LC_16_14_3 .LUT_INIT=16'b0010001001110010;
    LogicCell40 \pid_side.error_cry_2_c_RNI72F32_LC_16_14_3  (
            .in0(N__82741),
            .in1(N__77574),
            .in2(N__90613),
            .in3(N__80865),
            .lcout(\pid_side.m5_0_03_4_i_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_3_c_RNIPBV01_LC_16_14_4 .C_ON=1'b0;
    defparam \pid_side.error_cry_3_c_RNIPBV01_LC_16_14_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_3_c_RNIPBV01_LC_16_14_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \pid_side.error_cry_3_c_RNIPBV01_LC_16_14_4  (
            .in0(N__83085),
            .in1(N__77218),
            .in2(_gnd_net_),
            .in3(N__81103),
            .lcout(\pid_side.N_189 ),
            .ltout(\pid_side.N_189_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_2_c_RNI72F32_0_LC_16_14_5 .C_ON=1'b0;
    defparam \pid_side.error_cry_2_c_RNI72F32_0_LC_16_14_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_2_c_RNI72F32_0_LC_16_14_5 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \pid_side.error_cry_2_c_RNI72F32_0_LC_16_14_5  (
            .in0(N__82740),
            .in1(N__90544),
            .in2(N__66142),
            .in3(N__80864),
            .lcout(\pid_side.N_230 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_0_0_c_RNIAFOI3_LC_16_14_6 .C_ON=1'b0;
    defparam \pid_side.error_cry_0_0_c_RNIAFOI3_LC_16_14_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_0_c_RNIAFOI3_LC_16_14_6 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \pid_side.error_cry_0_0_c_RNIAFOI3_LC_16_14_6  (
            .in0(N__81318),
            .in1(N__66139),
            .in2(_gnd_net_),
            .in3(N__80312),
            .lcout(\pid_side.N_6 ),
            .ltout(\pid_side.N_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_1_17_LC_16_14_7 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_1_17_LC_16_14_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_1_17_LC_16_14_7 .LUT_INIT=16'b0100010100000001;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_1_17_LC_16_14_7  (
            .in0(N__89351),
            .in1(N__84188),
            .in2(N__66124),
            .in3(N__77612),
            .lcout(\pid_side.error_i_reg_esr_RNO_1_0_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_2_17_LC_16_15_0 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_2_17_LC_16_15_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_2_17_LC_16_15_0 .LUT_INIT=16'b1010000011100100;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_2_17_LC_16_15_0  (
            .in0(N__89572),
            .in1(N__89353),
            .in2(N__74692),
            .in3(N__73983),
            .lcout(\pid_front.N_262 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_5_c_RNI4NT91_LC_16_15_1 .C_ON=1'b0;
    defparam \pid_front.error_cry_5_c_RNI4NT91_LC_16_15_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_5_c_RNI4NT91_LC_16_15_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \pid_front.error_cry_5_c_RNI4NT91_LC_16_15_1  (
            .in0(N__83019),
            .in1(N__78413),
            .in2(_gnd_net_),
            .in3(N__74505),
            .lcout(\pid_front.N_245 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_2_16_LC_16_15_2 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_2_16_LC_16_15_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_2_16_LC_16_15_2 .LUT_INIT=16'b0000000100010001;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_2_16_LC_16_15_2  (
            .in0(N__68749),
            .in1(N__81145),
            .in2(N__85768),
            .in3(N__66241),
            .lcout(),
            .ltout(\pid_side.error_i_reg_esr_RNO_2Z0Z_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_16_LC_16_15_3 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_16_LC_16_15_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_16_LC_16_15_3 .LUT_INIT=16'b0110001001000000;
    LogicCell40 \pid_side.error_i_reg_esr_16_LC_16_15_3  (
            .in0(N__84509),
            .in1(N__66397),
            .in2(N__66121),
            .in3(N__66094),
            .lcout(\pid_side.error_i_regZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94213),
            .ce(N__86783),
            .sr(N__86398));
    defparam \pid_side.error_i_reg_esr_RNO_1_16_LC_16_15_4 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_1_16_LC_16_15_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_1_16_LC_16_15_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_1_16_LC_16_15_4  (
            .in0(_gnd_net_),
            .in1(N__89354),
            .in2(_gnd_net_),
            .in3(N__66100),
            .lcout(\pid_side.error_i_reg_esr_RNO_1Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_5_c_RNISBHI3_LC_16_15_5 .C_ON=1'b0;
    defparam \pid_side.error_cry_5_c_RNISBHI3_LC_16_15_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_5_c_RNISBHI3_LC_16_15_5 .LUT_INIT=16'b0011000000111010;
    LogicCell40 \pid_side.error_cry_5_c_RNISBHI3_LC_16_15_5  (
            .in0(N__89352),
            .in1(N__80089),
            .in2(N__84158),
            .in3(N__81526),
            .lcout(\pid_side.N_259 ),
            .ltout(\pid_side.N_259_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_2_14_LC_16_15_6 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_2_14_LC_16_15_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_2_14_LC_16_15_6 .LUT_INIT=16'b0101010100101010;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_2_14_LC_16_15_6  (
            .in0(N__86971),
            .in1(N__81314),
            .in2(N__66235),
            .in3(N__84508),
            .lcout(\pid_side.error_i_reg_esr_RNO_2Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_4_27_LC_16_16_0 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_4_27_LC_16_16_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_4_27_LC_16_16_0 .LUT_INIT=16'b0000000101010001;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_4_27_LC_16_16_0  (
            .in0(N__87800),
            .in1(N__72963),
            .in2(N__89601),
            .in3(N__66220),
            .lcout(\pid_front.N_338 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_4_c_RNIIEF61_LC_16_16_1 .C_ON=1'b0;
    defparam \pid_front.error_cry_4_c_RNIIEF61_LC_16_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_4_c_RNIIEF61_LC_16_16_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \pid_front.error_cry_4_c_RNIIEF61_LC_16_16_1  (
            .in0(N__80198),
            .in1(_gnd_net_),
            .in2(N__73793),
            .in3(N__73887),
            .lcout(\pid_front.N_163 ),
            .ltout(\pid_front.N_163_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_0_c_RNIFQ6J2_LC_16_16_2 .C_ON=1'b0;
    defparam \pid_front.error_cry_0_0_c_RNIFQ6J2_LC_16_16_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_0_c_RNIFQ6J2_LC_16_16_2 .LUT_INIT=16'b1000101110001011;
    LogicCell40 \pid_front.error_cry_0_0_c_RNIFQ6J2_LC_16_16_2  (
            .in0(N__74214),
            .in1(N__85165),
            .in2(N__66196),
            .in3(_gnd_net_),
            .lcout(\pid_front.N_186 ),
            .ltout(\pid_front.N_186_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_3_27_LC_16_16_3 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_3_27_LC_16_16_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_3_27_LC_16_16_3 .LUT_INIT=16'b0010101000000000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_3_27_LC_16_16_3  (
            .in0(N__87073),
            .in1(N__85716),
            .in2(N__66184),
            .in3(N__84477),
            .lcout(\pid_front.error_i_reg_9_sn_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_0_27_LC_16_16_4 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_27_LC_16_16_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_27_LC_16_16_4 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_27_LC_16_16_4  (
            .in0(N__81286),
            .in1(N__74374),
            .in2(_gnd_net_),
            .in3(N__66181),
            .lcout(),
            .ltout(\pid_front.N_42_i_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_27_LC_16_16_5 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_27_LC_16_16_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_27_LC_16_16_5 .LUT_INIT=16'b0000001110101010;
    LogicCell40 \pid_front.error_i_reg_esr_27_LC_16_16_5  (
            .in0(N__66355),
            .in1(N__66175),
            .in2(N__66166),
            .in3(N__66163),
            .lcout(\pid_front.error_i_regZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94229),
            .ce(N__78136),
            .sr(N__86388));
    defparam \pid_front.error_i_reg_esr_RNO_2_27_LC_16_16_6 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_2_27_LC_16_16_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_2_27_LC_16_16_6 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_2_27_LC_16_16_6  (
            .in0(N__84476),
            .in1(N__87072),
            .in2(_gnd_net_),
            .in3(N__80695),
            .lcout(\pid_front.error_i_reg_9_rn_0_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_2_20_LC_16_17_0 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_2_20_LC_16_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_2_20_LC_16_17_0 .LUT_INIT=16'b0011001100100011;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_2_20_LC_16_17_0  (
            .in0(N__87801),
            .in1(N__66349),
            .in2(N__89334),
            .in3(N__77083),
            .lcout(\pid_front.m24_2_03_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_4_20_LC_16_17_1 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_4_20_LC_16_17_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_4_20_LC_16_17_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_4_20_LC_16_17_1  (
            .in0(N__90671),
            .in1(N__90419),
            .in2(_gnd_net_),
            .in3(N__80648),
            .lcout(\pid_front.N_458 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_3_20_LC_16_17_2 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_3_20_LC_16_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_3_20_LC_16_17_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_3_20_LC_16_17_2  (
            .in0(N__83027),
            .in1(N__74319),
            .in2(_gnd_net_),
            .in3(N__74507),
            .lcout(),
            .ltout(\pid_front.N_314_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_1_20_LC_16_17_3 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_1_20_LC_16_17_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_1_20_LC_16_17_3 .LUT_INIT=16'b0000101000111011;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_1_20_LC_16_17_3  (
            .in0(N__90082),
            .in1(N__89291),
            .in2(N__66343),
            .in3(N__80649),
            .lcout(),
            .ltout(\pid_front.m24_2_03_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_0_20_LC_16_17_4 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_20_LC_16_17_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_20_LC_16_17_4 .LUT_INIT=16'b1111100011111111;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_20_LC_16_17_4  (
            .in0(N__66340),
            .in1(N__85739),
            .in2(N__66316),
            .in3(N__66313),
            .lcout(),
            .ltout(\pid_front.m24_2_03_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_20_LC_16_17_5 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_20_LC_16_17_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_20_LC_16_17_5 .LUT_INIT=16'b1000101000000010;
    LogicCell40 \pid_front.error_i_reg_esr_20_LC_16_17_5  (
            .in0(N__86935),
            .in1(N__84542),
            .in2(N__66307),
            .in3(N__73609),
            .lcout(\pid_front.error_i_regZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94245),
            .ce(N__78070),
            .sr(N__86380));
    defparam \pid_front.error_i_reg_esr_0_LC_16_18_0 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_0_LC_16_18_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_0_LC_16_18_0 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \pid_front.error_i_reg_esr_0_LC_16_18_0  (
            .in0(N__84180),
            .in1(N__82297),
            .in2(N__82064),
            .in3(N__69667),
            .lcout(\pid_front.error_i_regZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94263),
            .ce(N__78129),
            .sr(N__86374));
    defparam \pid_front.m80_0_a2_0_LC_16_18_1 .C_ON=1'b0;
    defparam \pid_front.m80_0_a2_0_LC_16_18_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.m80_0_a2_0_LC_16_18_1 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \pid_front.m80_0_a2_0_LC_16_18_1  (
            .in0(N__86902),
            .in1(N__89300),
            .in2(_gnd_net_),
            .in3(N__84473),
            .lcout(pid_side_N_607),
            .ltout(pid_side_N_607_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_2_LC_16_18_2 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_2_LC_16_18_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_2_LC_16_18_2 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \pid_front.error_i_reg_esr_2_LC_16_18_2  (
            .in0(N__84179),
            .in1(N__66265),
            .in2(N__66451),
            .in3(N__66448),
            .lcout(\pid_front.error_i_regZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94263),
            .ce(N__78129),
            .sr(N__86374));
    defparam \pid_front.error_i_reg_esr_1_LC_16_18_3 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_1_LC_16_18_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_1_LC_16_18_3 .LUT_INIT=16'b1011000000010000;
    LogicCell40 \pid_front.error_i_reg_esr_1_LC_16_18_3  (
            .in0(N__84133),
            .in1(N__69601),
            .in2(N__82051),
            .in3(N__69582),
            .lcout(\pid_front.error_i_regZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94263),
            .ce(N__78129),
            .sr(N__86374));
    defparam \pid_front.OVER_0_a3_LC_16_18_4 .C_ON=1'b0;
    defparam \pid_front.OVER_0_a3_LC_16_18_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.OVER_0_a3_LC_16_18_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \pid_front.OVER_0_a3_LC_16_18_4  (
            .in0(N__68712),
            .in1(N__70065),
            .in2(_gnd_net_),
            .in3(N__70023),
            .lcout(pid_front_N_335),
            .ltout(pid_front_N_335_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_6_16_LC_16_18_5 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_6_16_LC_16_18_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_6_16_LC_16_18_5 .LUT_INIT=16'b0011110000101100;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_6_16_LC_16_18_5  (
            .in0(N__89111),
            .in1(N__84474),
            .in2(N__66415),
            .in3(N__85157),
            .lcout(),
            .ltout(\pid_side.error_i_reg_9_1_rn_sx_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_3_16_LC_16_18_6 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_3_16_LC_16_18_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_3_16_LC_16_18_6 .LUT_INIT=16'b1111010011110000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_3_16_LC_16_18_6  (
            .in0(N__84475),
            .in1(N__86903),
            .in2(N__66412),
            .in3(N__85925),
            .lcout(),
            .ltout(\pid_side.error_i_reg_9_1_rn_0_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_16_LC_16_18_7 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_16_LC_16_18_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_16_LC_16_18_7 .LUT_INIT=16'b0101000011111010;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_16_LC_16_18_7  (
            .in0(N__66409),
            .in1(_gnd_net_),
            .in2(N__66400),
            .in3(N__77368),
            .lcout(\pid_side.error_i_reg_9_1_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.state_RNIRT3N4_1_LC_16_19_1 .C_ON=1'b0;
    defparam \pid_front.state_RNIRT3N4_1_LC_16_19_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.state_RNIRT3N4_1_LC_16_19_1 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \pid_front.state_RNIRT3N4_1_LC_16_19_1  (
            .in0(N__70496),
            .in1(N__71030),
            .in2(_gnd_net_),
            .in3(N__76010),
            .lcout(),
            .ltout(\pid_front.N_600_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNILUUMB_3_LC_16_19_2 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNILUUMB_3_LC_16_19_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNILUUMB_3_LC_16_19_2 .LUT_INIT=16'b1101010111000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNILUUMB_3_LC_16_19_2  (
            .in0(N__70116),
            .in1(N__74605),
            .in2(N__66388),
            .in3(N__66559),
            .lcout(\pid_front.error_i_acumm_13_0_tz_1_0 ),
            .ltout(\pid_front.error_i_acumm_13_0_tz_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_0_LC_16_19_3 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_0_LC_16_19_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_0_LC_16_19_3 .LUT_INIT=16'b1010101010101000;
    LogicCell40 \pid_front.error_i_acumm_0_LC_16_19_3  (
            .in0(N__66385),
            .in1(N__70091),
            .in2(N__66376),
            .in3(N__66896),
            .lcout(\pid_front.error_i_acummZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94281),
            .ce(N__75767),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_1_LC_16_19_4 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_1_LC_16_19_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_1_LC_16_19_4 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \pid_front.error_i_acumm_1_LC_16_19_4  (
            .in0(N__66897),
            .in1(N__75580),
            .in2(N__70096),
            .in3(N__66510),
            .lcout(\pid_front.error_i_acummZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94281),
            .ce(N__75767),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_2_LC_16_19_5 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_2_LC_16_19_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_2_LC_16_19_5 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \pid_front.error_i_acumm_2_LC_16_19_5  (
            .in0(N__66511),
            .in1(N__70095),
            .in2(N__75529),
            .in3(N__66898),
            .lcout(\pid_front.error_i_acummZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94281),
            .ce(N__75767),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNI6EER_14_LC_16_19_6 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI6EER_14_LC_16_19_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI6EER_14_LC_16_19_6 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNI6EER_14_LC_16_19_6  (
            .in0(N__69895),
            .in1(N__69850),
            .in2(_gnd_net_),
            .in3(N__69930),
            .lcout(\pid_front.error_i_acumm_13_i_o2_0_7_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNIRESC_12_LC_16_20_0 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIRESC_12_LC_16_20_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIRESC_12_LC_16_20_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNIRESC_12_LC_16_20_0  (
            .in0(_gnd_net_),
            .in1(N__75671),
            .in2(_gnd_net_),
            .in3(N__66571),
            .lcout(\pid_front.N_530 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_6_LC_16_20_1 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_6_LC_16_20_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_6_LC_16_20_1 .LUT_INIT=16'b0100010001010100;
    LogicCell40 \pid_front.error_i_acumm_6_LC_16_20_1  (
            .in0(N__66472),
            .in1(N__75196),
            .in2(N__75962),
            .in3(N__66558),
            .lcout(\pid_front.error_i_acummZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94297),
            .ce(N__75764),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_5_LC_16_20_2 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_5_LC_16_20_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_5_LC_16_20_2 .LUT_INIT=16'b0000000011011100;
    LogicCell40 \pid_front.error_i_acumm_5_LC_16_20_2  (
            .in0(N__66556),
            .in1(N__75250),
            .in2(N__75967),
            .in3(N__66471),
            .lcout(\pid_front.error_i_acummZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94297),
            .ce(N__75764),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNIR7I45_10_LC_16_20_3 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIR7I45_10_LC_16_20_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIR7I45_10_LC_16_20_3 .LUT_INIT=16'b0000000000011111;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNIR7I45_10_LC_16_20_3  (
            .in0(N__75031),
            .in1(N__75115),
            .in2(N__75676),
            .in3(N__76009),
            .lcout(\pid_front.N_633 ),
            .ltout(\pid_front.N_633_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNIMLH86_28_LC_16_20_4 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIMLH86_28_LC_16_20_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIMLH86_28_LC_16_20_4 .LUT_INIT=16'b1101110111001101;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNIMLH86_28_LC_16_20_4  (
            .in0(N__75958),
            .in1(N__75850),
            .in2(N__66481),
            .in3(N__66478),
            .lcout(\pid_front.N_251 ),
            .ltout(\pid_front.N_251_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_4_LC_16_20_5 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_4_LC_16_20_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_4_LC_16_20_5 .LUT_INIT=16'b0000110000001110;
    LogicCell40 \pid_front.error_i_acumm_4_LC_16_20_5  (
            .in0(N__75940),
            .in1(N__75484),
            .in2(N__66463),
            .in3(N__66557),
            .lcout(\pid_front.error_i_acummZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94297),
            .ce(N__75764),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_7_LC_16_20_6 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_7_LC_16_20_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_7_LC_16_20_6 .LUT_INIT=16'b0101000001010001;
    LogicCell40 \pid_front.error_i_acumm_7_LC_16_20_6  (
            .in0(N__70183),
            .in1(N__75942),
            .in2(N__75412),
            .in3(N__70149),
            .lcout(\pid_front.error_i_acummZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94297),
            .ce(N__75764),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_8_LC_16_20_7 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_8_LC_16_20_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_8_LC_16_20_7 .LUT_INIT=16'b0011001100000001;
    LogicCell40 \pid_front.error_i_acumm_8_LC_16_20_7  (
            .in0(N__75941),
            .in1(N__70182),
            .in2(N__70150),
            .in3(N__75355),
            .lcout(\pid_front.error_i_acummZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94297),
            .ce(N__75764),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_RNO_0_3_LC_16_21_0 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_RNO_0_3_LC_16_21_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_RNO_0_3_LC_16_21_0 .LUT_INIT=16'b0000101111111011;
    LogicCell40 \pid_front.error_i_acumm_RNO_0_3_LC_16_21_0  (
            .in0(N__76012),
            .in1(N__66532),
            .in2(N__75939),
            .in3(N__66555),
            .lcout(),
            .ltout(\pid_front.N_62_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_3_LC_16_21_1 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_3_LC_16_21_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_3_LC_16_21_1 .LUT_INIT=16'b0101010001010100;
    LogicCell40 \pid_front.error_i_acumm_3_LC_16_21_1  (
            .in0(N__75849),
            .in1(N__74569),
            .in2(N__66586),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_i_acummZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94312),
            .ce(N__75768),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNISDO3_0_7_LC_16_21_2 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNISDO3_0_7_LC_16_21_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNISDO3_0_7_LC_16_21_2 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNISDO3_0_7_LC_16_21_2  (
            .in0(N__70169),
            .in1(N__75353),
            .in2(_gnd_net_),
            .in3(N__75407),
            .lcout(\pid_front.N_177 ),
            .ltout(\pid_front.N_177_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNIMD4V_10_LC_16_21_3 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIMD4V_10_LC_16_21_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIMD4V_10_LC_16_21_3 .LUT_INIT=16'b0101010101110101;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNIMD4V_10_LC_16_21_3  (
            .in0(N__75669),
            .in1(N__75027),
            .in2(N__66565),
            .in3(N__75111),
            .lcout(\pid_front.N_181 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNISDO3_7_LC_16_21_4 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNISDO3_7_LC_16_21_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNISDO3_7_LC_16_21_4 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNISDO3_7_LC_16_21_4  (
            .in0(N__70170),
            .in1(N__75354),
            .in2(_gnd_net_),
            .in3(N__75408),
            .lcout(),
            .ltout(\pid_front.N_158_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNINLA85_12_LC_16_21_5 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNINLA85_12_LC_16_21_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNINLA85_12_LC_16_21_5 .LUT_INIT=16'b0000000011011100;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNINLA85_12_LC_16_21_5  (
            .in0(N__70410),
            .in1(N__75675),
            .in2(N__66562),
            .in3(N__75055),
            .lcout(\pid_front.N_601 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_RNO_1_3_LC_16_21_6 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_RNO_1_3_LC_16_21_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_RNO_1_3_LC_16_21_6 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \pid_front.error_i_acumm_RNO_1_3_LC_16_21_6  (
            .in0(N__75483),
            .in1(N__74617),
            .in2(_gnd_net_),
            .in3(N__66525),
            .lcout(\pid_front.N_208 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNINKDV5_28_LC_16_21_7 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNINKDV5_28_LC_16_21_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNINKDV5_28_LC_16_21_7 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNINKDV5_28_LC_16_21_7  (
            .in0(N__66526),
            .in1(N__75909),
            .in2(N__75861),
            .in3(N__76011),
            .lcout(\pid_front.N_483 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNINO362_0_21_LC_16_22_0 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNINO362_0_21_LC_16_22_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNINO362_0_21_LC_16_22_0 .LUT_INIT=16'b0010010011011011;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNINO362_0_21_LC_16_22_0  (
            .in0(N__66694),
            .in1(N__67043),
            .in2(N__91755),
            .in3(N__66834),
            .lcout(\pid_front.un1_pid_prereg_0_25 ),
            .ltout(\pid_front.un1_pid_prereg_0_25_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIDF6C4_21_LC_16_22_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIDF6C4_21_LC_16_22_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIDF6C4_21_LC_16_22_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIDF6C4_21_LC_16_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__66880),
            .in3(N__66798),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIDF6C4Z0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNO_0_30_LC_16_22_2 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNO_0_30_LC_16_22_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNO_0_30_LC_16_22_2 .LUT_INIT=16'b1000011101111000;
    LogicCell40 \pid_front.pid_prereg_esr_RNO_0_30_LC_16_22_2  (
            .in0(N__66815),
            .in1(N__66739),
            .in2(N__66820),
            .in3(N__66740),
            .lcout(\pid_front.un1_pid_prereg_0_axb_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIR0EO8_21_LC_16_22_3 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIR0EO8_21_LC_16_22_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIR0EO8_21_LC_16_22_3 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIR0EO8_21_LC_16_22_3  (
            .in0(N__66799),
            .in1(N__66742),
            .in2(N__66819),
            .in3(N__66741),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIR0EO8Z0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNINO362_21_LC_16_22_4 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNINO362_21_LC_16_22_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNINO362_21_LC_16_22_4 .LUT_INIT=16'b1111101100100000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNINO362_21_LC_16_22_4  (
            .in0(N__66695),
            .in1(N__67044),
            .in2(N__91756),
            .in3(N__66833),
            .lcout(\pid_front.un1_pid_prereg_0_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIMM262_21_LC_16_22_5 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIMM262_21_LC_16_22_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIMM262_21_LC_16_22_5 .LUT_INIT=16'b1110111100001000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIMM262_21_LC_16_22_5  (
            .in0(N__91740),
            .in1(N__66693),
            .in2(N__67071),
            .in3(N__69866),
            .lcout(\pid_front.un1_pid_prereg_0_24 ),
            .ltout(\pid_front.un1_pid_prereg_0_24_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNINPAO8_21_LC_16_22_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNINPAO8_21_LC_16_22_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNINPAO8_21_LC_16_22_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNINPAO8_21_LC_16_22_6  (
            .in0(N__66787),
            .in1(N__66766),
            .in2(N__66745),
            .in3(N__66738),
            .lcout(\pid_front.error_d_reg_prev_esr_RNINPAO8Z0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIASE61_21_LC_16_22_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIASE61_21_LC_16_22_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIASE61_21_LC_16_22_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIASE61_21_LC_16_22_7  (
            .in0(N__67039),
            .in1(N__91730),
            .in2(_gnd_net_),
            .in3(N__66692),
            .lcout(\pid_front.un1_pid_prereg_370_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_14_LC_16_23_0 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_14_LC_16_23_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_14_LC_16_23_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_14_LC_16_23_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__94540),
            .lcout(\pid_front.error_d_reg_prevZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94343),
            .ce(N__71795),
            .sr(N__71704));
    defparam \pid_front.error_d_reg_prev_esr_15_LC_16_23_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_15_LC_16_23_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_15_LC_16_23_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_15_LC_16_23_1  (
            .in0(N__94495),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prevZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94343),
            .ce(N__71795),
            .sr(N__71704));
    defparam \pid_front.error_d_reg_prev_esr_19_LC_16_23_2 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_19_LC_16_23_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_19_LC_16_23_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_19_LC_16_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__91816),
            .lcout(\pid_front.error_d_reg_prevZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94343),
            .ce(N__71795),
            .sr(N__71704));
    defparam \pid_front.error_d_reg_prev_esr_20_LC_16_23_3 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_20_LC_16_23_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_20_LC_16_23_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_20_LC_16_23_3  (
            .in0(N__91858),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prevZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94343),
            .ce(N__71795),
            .sr(N__71704));
    defparam \pid_front.error_d_reg_prev_esr_21_LC_16_23_4 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_21_LC_16_23_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_21_LC_16_23_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_21_LC_16_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__91754),
            .lcout(\pid_front.error_d_reg_prevZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94343),
            .ce(N__71795),
            .sr(N__71704));
    defparam \pid_front.error_d_reg_prev_esr_4_LC_16_23_5 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_4_LC_16_23_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_4_LC_16_23_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_4_LC_16_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66997),
            .lcout(\pid_front.error_d_reg_prevZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94343),
            .ce(N__71795),
            .sr(N__71704));
    defparam \pid_front.error_d_reg_prev_esr_8_LC_16_23_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_8_LC_16_23_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_8_LC_16_23_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_8_LC_16_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78806),
            .lcout(\pid_front.error_d_reg_prevZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94343),
            .ce(N__71795),
            .sr(N__71704));
    defparam \pid_front.error_d_reg_prev_esr_9_LC_16_23_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_9_LC_16_23_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_9_LC_16_23_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_9_LC_16_23_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78739),
            .lcout(\pid_front.error_d_reg_prevZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94343),
            .ce(N__71795),
            .sr(N__71704));
    defparam \pid_front.error_p_reg_esr_RNI6R6D1_8_LC_16_24_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI6R6D1_8_LC_16_24_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI6R6D1_8_LC_16_24_0 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_front.error_p_reg_esr_RNI6R6D1_8_LC_16_24_0  (
            .in0(N__66921),
            .in1(N__71286),
            .in2(_gnd_net_),
            .in3(N__66934),
            .lcout(\pid_front.error_p_reg_esr_RNI6R6D1Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_9_LC_16_24_1 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_9_LC_16_24_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_9_LC_16_24_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_9_LC_16_24_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66922),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94358),
            .ce(N__75322),
            .sr(N__86355));
    defparam \pid_front.error_p_reg_esr_RNI8NB61_11_LC_16_24_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI8NB61_11_LC_16_24_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI8NB61_11_LC_16_24_2 .LUT_INIT=16'b1111010101010000;
    LogicCell40 \pid_front.error_p_reg_esr_RNI8NB61_11_LC_16_24_2  (
            .in0(N__71854),
            .in1(_gnd_net_),
            .in2(N__71950),
            .in3(N__94591),
            .lcout(\pid_front.g0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI8NB61_1_11_LC_16_24_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI8NB61_1_11_LC_16_24_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI8NB61_1_11_LC_16_24_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_p_reg_esr_RNI8NB61_1_11_LC_16_24_3  (
            .in0(N__94590),
            .in1(N__71946),
            .in2(_gnd_net_),
            .in3(N__71853),
            .lcout(\pid_front.error_p_reg_esr_RNI8NB61_1Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIH0C61_0_14_LC_16_24_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIH0C61_0_14_LC_16_24_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIH0C61_0_14_LC_16_24_4 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_p_reg_esr_RNIH0C61_0_14_LC_16_24_4  (
            .in0(N__67544),
            .in1(N__67583),
            .in2(_gnd_net_),
            .in3(N__94519),
            .lcout(\pid_front.error_p_reg_esr_RNIH0C61_0Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIH0C61_14_LC_16_24_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIH0C61_14_LC_16_24_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIH0C61_14_LC_16_24_5 .LUT_INIT=16'b1011001010110010;
    LogicCell40 \pid_front.error_p_reg_esr_RNIH0C61_14_LC_16_24_5  (
            .in0(N__94520),
            .in1(N__67545),
            .in2(N__67588),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_p_reg_esr_RNIH0C61Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIK3C61_0_15_LC_16_24_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIK3C61_0_15_LC_16_24_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIK3C61_0_15_LC_16_24_6 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_p_reg_esr_RNIK3C61_0_15_LC_16_24_6  (
            .in0(N__67716),
            .in1(N__67143),
            .in2(_gnd_net_),
            .in3(N__94487),
            .lcout(\pid_front.error_p_reg_esr_RNIK3C61_0Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIK3C61_15_LC_16_24_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIK3C61_15_LC_16_24_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIK3C61_15_LC_16_24_7 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \pid_front.error_p_reg_esr_RNIK3C61_15_LC_16_24_7  (
            .in0(N__94488),
            .in1(_gnd_net_),
            .in2(N__67147),
            .in3(N__67717),
            .lcout(\pid_front.error_p_reg_esr_RNIK3C61Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_fast_esr_RNI5VGK_12_LC_16_25_0 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_fast_esr_RNI5VGK_12_LC_16_25_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_fast_esr_RNI5VGK_12_LC_16_25_0 .LUT_INIT=16'b1101110111101110;
    LogicCell40 \pid_front.error_d_reg_fast_esr_RNI5VGK_12_LC_16_25_0  (
            .in0(N__71969),
            .in1(N__71905),
            .in2(_gnd_net_),
            .in3(N__67427),
            .lcout(\pid_front.error_d_reg_fast_esr_RNI5VGKZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_fast_esr_RNID6KB1_12_LC_16_25_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_fast_esr_RNID6KB1_12_LC_16_25_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_fast_esr_RNID6KB1_12_LC_16_25_1 .LUT_INIT=16'b1111011001100000;
    LogicCell40 \pid_front.error_d_reg_fast_esr_RNID6KB1_12_LC_16_25_1  (
            .in0(N__67428),
            .in1(N__71970),
            .in2(N__71913),
            .in3(N__67465),
            .lcout(),
            .ltout(\pid_front.error_d_reg_fast_esr_RNID6KB1Z0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_fast_esr_RNIQSG63_12_LC_16_25_2 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_fast_esr_RNIQSG63_12_LC_16_25_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_fast_esr_RNIQSG63_12_LC_16_25_2 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \pid_front.error_d_reg_fast_esr_RNIQSG63_12_LC_16_25_2  (
            .in0(_gnd_net_),
            .in1(N__67123),
            .in2(N__67117),
            .in3(N__67448),
            .lcout(\pid_front.error_d_reg_fast_esr_RNIQSG63Z0Z_12 ),
            .ltout(\pid_front.error_d_reg_fast_esr_RNIQSG63Z0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIK42C6_14_LC_16_25_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIK42C6_14_LC_16_25_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIK42C6_14_LC_16_25_3 .LUT_INIT=16'b1110100010001000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIK42C6_14_LC_16_25_3  (
            .in0(N__67269),
            .in1(N__67284),
            .in2(N__67288),
            .in3(N__67248),
            .lcout(),
            .ltout(\pid_front.error_p_reg_esr_RNIK42C6Z0Z_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNI13Q1D_12_LC_16_25_4 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNI13Q1D_12_LC_16_25_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNI13Q1D_12_LC_16_25_4 .LUT_INIT=16'b1110111011110000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNI13Q1D_12_LC_16_25_4  (
            .in0(N__67285),
            .in1(N__67270),
            .in2(N__67261),
            .in3(N__67255),
            .lcout(\pid_front.error_d_reg_prev_esr_RNI13Q1DZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNILTVH2_0_12_LC_16_25_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNILTVH2_0_12_LC_16_25_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNILTVH2_0_12_LC_16_25_5 .LUT_INIT=16'b0000110001001101;
    LogicCell40 \pid_front.error_p_reg_esr_RNILTVH2_0_12_LC_16_25_5  (
            .in0(N__67447),
            .in1(N__67194),
            .in2(N__71914),
            .in3(N__67466),
            .lcout(),
            .ltout(\pid_front.un1_pid_prereg_167_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIE0094_12_LC_16_25_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIE0094_12_LC_16_25_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIE0094_12_LC_16_25_6 .LUT_INIT=16'b1010111100100011;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIE0094_12_LC_16_25_6  (
            .in0(N__67247),
            .in1(N__78682),
            .in2(N__67258),
            .in3(N__81834),
            .lcout(\pid_front.un1_pid_prereg_167_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIJVGT4_12_LC_16_25_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIJVGT4_12_LC_16_25_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIJVGT4_12_LC_16_25_7 .LUT_INIT=16'b1001110001100011;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIJVGT4_12_LC_16_25_7  (
            .in0(N__81835),
            .in1(N__67249),
            .in2(N__78695),
            .in3(N__67234),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIJVGT4Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNILTVH2_12_LC_16_26_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNILTVH2_12_LC_16_26_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNILTVH2_12_LC_16_26_0 .LUT_INIT=16'b0011110001101001;
    LogicCell40 \pid_front.error_p_reg_esr_RNILTVH2_12_LC_16_26_0  (
            .in0(N__67449),
            .in1(N__67195),
            .in2(N__71912),
            .in3(N__67467),
            .lcout(\pid_front.error_p_reg_esr_RNILTVH2Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_fast_esr_RNIOTBC_12_LC_16_26_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_fast_esr_RNIOTBC_12_LC_16_26_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_fast_esr_RNIOTBC_12_LC_16_26_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \pid_front.error_d_reg_fast_esr_RNIOTBC_12_LC_16_26_1  (
            .in0(_gnd_net_),
            .in1(N__67426),
            .in2(_gnd_net_),
            .in3(N__71968),
            .lcout(\pid_front.N_2394_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIUO6U_2_12_LC_16_26_2 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIUO6U_2_12_LC_16_26_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIUO6U_2_12_LC_16_26_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIUO6U_2_12_LC_16_26_2  (
            .in0(_gnd_net_),
            .in1(N__78689),
            .in2(_gnd_net_),
            .in3(N__81823),
            .lcout(),
            .ltout(\pid_front.N_3_i_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIROQ33_12_LC_16_26_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIROQ33_12_LC_16_26_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIROQ33_12_LC_16_26_3 .LUT_INIT=16'b0000001100010111;
    LogicCell40 \pid_front.error_p_reg_esr_RNIROQ33_12_LC_16_26_3  (
            .in0(N__67468),
            .in1(N__71902),
            .in2(N__67183),
            .in3(N__67450),
            .lcout(\pid_front.N_3_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI873N_11_LC_16_26_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI873N_11_LC_16_26_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI873N_11_LC_16_26_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \pid_front.error_p_reg_esr_RNI873N_11_LC_16_26_4  (
            .in0(_gnd_net_),
            .in1(N__71935),
            .in2(_gnd_net_),
            .in3(N__71842),
            .lcout(\pid_front.un1_pid_prereg_79 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI8NB61_0_11_LC_16_26_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI8NB61_0_11_LC_16_26_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI8NB61_0_11_LC_16_26_5 .LUT_INIT=16'b1111010100000000;
    LogicCell40 \pid_front.error_p_reg_esr_RNI8NB61_0_11_LC_16_26_5  (
            .in0(N__71843),
            .in1(_gnd_net_),
            .in2(N__71945),
            .in3(N__94587),
            .lcout(\pid_front.un1_pid_prereg_135_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_fast_esr_12_LC_16_26_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_fast_esr_12_LC_16_26_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_fast_esr_12_LC_16_26_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_prev_fast_esr_12_LC_16_26_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81825),
            .lcout(\pid_front.error_d_reg_prev_fastZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94375),
            .ce(N__71817),
            .sr(N__71715));
    defparam \pid_front.error_d_reg_prev_esr_12_LC_16_26_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_12_LC_16_26_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_12_LC_16_26_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_12_LC_16_26_7  (
            .in0(N__81824),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prevZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94375),
            .ce(N__71817),
            .sr(N__71715));
    defparam \pid_front.error_p_reg_esr_0_LC_16_27_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_0_LC_16_27_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_0_LC_16_27_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_0_LC_16_27_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67408),
            .lcout(\pid_front.error_p_regZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94383),
            .ce(N__93394),
            .sr(N__93006));
    defparam \pid_front.error_p_reg_esr_10_LC_16_27_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_10_LC_16_27_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_10_LC_16_27_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_10_LC_16_27_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67369),
            .lcout(\pid_front.error_p_regZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94383),
            .ce(N__93394),
            .sr(N__93006));
    defparam \pid_front.error_p_reg_esr_11_LC_16_27_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_11_LC_16_27_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_11_LC_16_27_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_11_LC_16_27_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67348),
            .lcout(\pid_front.error_p_regZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94383),
            .ce(N__93394),
            .sr(N__93006));
    defparam \pid_front.error_p_reg_esr_12_LC_16_27_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_12_LC_16_27_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_12_LC_16_27_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_12_LC_16_27_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67327),
            .lcout(\pid_front.error_p_regZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94383),
            .ce(N__93394),
            .sr(N__93006));
    defparam \pid_front.error_p_reg_esr_14_LC_16_27_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_14_LC_16_27_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_14_LC_16_27_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_14_LC_16_27_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67306),
            .lcout(\pid_front.error_p_regZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94383),
            .ce(N__93394),
            .sr(N__93006));
    defparam \pid_front.error_p_reg_esr_15_LC_16_27_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_15_LC_16_27_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_15_LC_16_27_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_p_reg_esr_15_LC_16_27_6  (
            .in0(N__67735),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_p_regZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94383),
            .ce(N__93394),
            .sr(N__93006));
    defparam \pid_front.error_d_reg_fast_esr_RNIR9PO_13_LC_16_28_2 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_fast_esr_RNIR9PO_13_LC_16_28_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_fast_esr_RNIR9PO_13_LC_16_28_2 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_front.error_d_reg_fast_esr_RNIR9PO_13_LC_16_28_2  (
            .in0(N__67688),
            .in1(N__67640),
            .in2(_gnd_net_),
            .in3(N__67600),
            .lcout(),
            .ltout(\pid_front.N_2401_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNICA5V1_14_LC_16_28_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNICA5V1_14_LC_16_28_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNICA5V1_14_LC_16_28_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \pid_front.error_p_reg_esr_RNICA5V1_14_LC_16_28_3  (
            .in0(N__67587),
            .in1(N__67558),
            .in2(N__67531),
            .in3(N__94535),
            .lcout(),
            .ltout(\pid_front.g0_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIBIFG6_12_LC_16_28_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIBIFG6_12_LC_16_28_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIBIFG6_12_LC_16_28_4 .LUT_INIT=16'b1101001001001011;
    LogicCell40 \pid_front.error_p_reg_esr_RNIBIFG6_12_LC_16_28_4  (
            .in0(N__71863),
            .in1(N__67528),
            .in2(N__67519),
            .in3(N__71869),
            .lcout(\pid_front.error_p_reg_esr_RNIBIFG6Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNISKLO_0_20_LC_17_4_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNISKLO_0_20_LC_17_4_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNISKLO_0_20_LC_17_4_0 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNISKLO_0_20_LC_17_4_0  (
            .in0(N__91594),
            .in1(N__67491),
            .in2(_gnd_net_),
            .in3(N__91085),
            .lcout(\pid_side.error_d_reg_prev_esr_RNISKLO_0Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_20_LC_17_4_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_20_LC_17_4_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_20_LC_17_4_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_20_LC_17_4_1  (
            .in0(N__91087),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94107),
            .ce(N__88078),
            .sr(N__87950));
    defparam \pid_side.error_d_reg_prev_esr_RNISKLO_20_LC_17_4_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNISKLO_20_LC_17_4_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNISKLO_20_LC_17_4_2 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNISKLO_20_LC_17_4_2  (
            .in0(N__91595),
            .in1(N__67492),
            .in2(_gnd_net_),
            .in3(N__91086),
            .lcout(\pid_side.error_d_reg_prev_esr_RNISKLOZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNI5SNH3_7_LC_17_4_3 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNI5SNH3_7_LC_17_4_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNI5SNH3_7_LC_17_4_3 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_side.error_p_reg_esr_RNI5SNH3_7_LC_17_4_3  (
            .in0(N__72358),
            .in1(N__72223),
            .in2(_gnd_net_),
            .in3(N__72199),
            .lcout(\pid_side.error_p_reg_esr_RNI5SNH3Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIOUJE2_6_LC_17_5_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIOUJE2_6_LC_17_5_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIOUJE2_6_LC_17_5_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIOUJE2_6_LC_17_5_2  (
            .in0(N__72238),
            .in1(N__76129),
            .in2(_gnd_net_),
            .in3(N__76249),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIOUJE2Z0Z_6 ),
            .ltout(\pid_side.error_d_reg_prev_esr_RNIOUJE2Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI44E63_6_LC_17_5_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI44E63_6_LC_17_5_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI44E63_6_LC_17_5_3 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI44E63_6_LC_17_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__67864),
            .in3(N__67850),
            .lcout(),
            .ltout(\pid_side.un1_pid_prereg_66_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIRH187_5_LC_17_5_4 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIRH187_5_LC_17_5_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIRH187_5_LC_17_5_4 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pid_side.error_p_reg_esr_RNIRH187_5_LC_17_5_4  (
            .in0(N__76078),
            .in1(N__76119),
            .in2(N__67861),
            .in3(N__76060),
            .lcout(\pid_side.error_p_reg_esr_RNIRH187Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_5_LC_17_5_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_5_LC_17_5_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_5_LC_17_5_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_5_LC_17_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78622),
            .lcout(\pid_side.error_d_reg_prevZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94114),
            .ce(N__88088),
            .sr(N__87947));
    defparam \pid_side.error_p_reg_esr_RNIBABR4_5_LC_17_5_6 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIBABR4_5_LC_17_5_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIBABR4_5_LC_17_5_6 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_side.error_p_reg_esr_RNIBABR4_5_LC_17_5_6  (
            .in0(N__67851),
            .in1(N__67825),
            .in2(_gnd_net_),
            .in3(N__76120),
            .lcout(\pid_side.error_p_reg_esr_RNIBABR4Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI8UIO_0_15_LC_17_6_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI8UIO_0_15_LC_17_6_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI8UIO_0_15_LC_17_6_0 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI8UIO_0_15_LC_17_6_0  (
            .in0(N__90813),
            .in1(N__67791),
            .in2(_gnd_net_),
            .in3(N__91538),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI8UIO_0Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_15_LC_17_6_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_15_LC_17_6_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_15_LC_17_6_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_15_LC_17_6_1  (
            .in0(N__91540),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94121),
            .ce(N__88087),
            .sr(N__87945));
    defparam \pid_side.error_d_reg_prev_esr_RNI8UIO_15_LC_17_6_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI8UIO_15_LC_17_6_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI8UIO_15_LC_17_6_2 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI8UIO_15_LC_17_6_2  (
            .in0(N__90814),
            .in1(N__67792),
            .in2(_gnd_net_),
            .in3(N__91539),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI8UIOZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIE4JO_17_LC_17_6_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIE4JO_17_LC_17_6_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIE4JO_17_LC_17_6_3 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIE4JO_17_LC_17_6_3  (
            .in0(N__90790),
            .in1(N__67749),
            .in2(_gnd_net_),
            .in3(N__91169),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIE4JOZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_17_LC_17_6_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_17_LC_17_6_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_17_LC_17_6_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_17_LC_17_6_4  (
            .in0(N__91170),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94121),
            .ce(N__88087),
            .sr(N__87945));
    defparam \pid_side.error_d_reg_prev_esr_RNIGI4KK_12_LC_17_6_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIGI4KK_12_LC_17_6_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIGI4KK_12_LC_17_6_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIGI4KK_12_LC_17_6_5  (
            .in0(N__76485),
            .in1(N__68036),
            .in2(_gnd_net_),
            .in3(N__68588),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIGI4KKZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNICCO8B_12_LC_17_6_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNICCO8B_12_LC_17_6_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNICCO8B_12_LC_17_6_6 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNICCO8B_12_LC_17_6_6  (
            .in0(N__68589),
            .in1(_gnd_net_),
            .in2(N__68041),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prev_esr_RNICCO8BZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIBNLL9_18_LC_17_7_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIBNLL9_18_LC_17_7_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIBNLL9_18_LC_17_7_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIBNLL9_18_LC_17_7_0  (
            .in0(N__67929),
            .in1(N__68071),
            .in2(N__68110),
            .in3(N__67943),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIBNLL9Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI2BI34_21_LC_17_7_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI2BI34_21_LC_17_7_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI2BI34_21_LC_17_7_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI2BI34_21_LC_17_7_1  (
            .in0(_gnd_net_),
            .in1(N__67956),
            .in2(_gnd_net_),
            .in3(N__67917),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI2BI34Z0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIKSEL1_0_21_LC_17_7_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIKSEL1_0_21_LC_17_7_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIKSEL1_0_21_LC_17_7_2 .LUT_INIT=16'b0001100011100111;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIKSEL1_0_21_LC_17_7_2  (
            .in0(N__91647),
            .in1(N__91379),
            .in2(N__72951),
            .in3(N__67989),
            .lcout(\pid_side.un1_pid_prereg_0_13 ),
            .ltout(\pid_side.un1_pid_prereg_0_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIR9TU8_21_LC_17_7_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIR9TU8_21_LC_17_7_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIR9TU8_21_LC_17_7_3 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIR9TU8_21_LC_17_7_3  (
            .in0(N__67944),
            .in1(N__67930),
            .in2(N__67921),
            .in3(N__67916),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIR9TU8Z0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNO_0_30_LC_17_7_4 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNO_0_30_LC_17_7_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNO_0_30_LC_17_7_4 .LUT_INIT=16'b1000011101111000;
    LogicCell40 \pid_side.pid_prereg_esr_RNO_0_30_LC_17_7_4  (
            .in0(N__72585),
            .in1(N__72756),
            .in2(N__72589),
            .in3(N__72757),
            .lcout(\pid_side.un1_pid_prereg_0_axb_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIUBKL1_21_LC_17_7_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIUBKL1_21_LC_17_7_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIUBKL1_21_LC_17_7_5 .LUT_INIT=16'b1110111100001000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIUBKL1_21_LC_17_7_5  (
            .in0(N__91380),
            .in1(N__91648),
            .in2(N__72952),
            .in3(N__67891),
            .lcout(\pid_side.un1_pid_prereg_0_24 ),
            .ltout(\pid_side.un1_pid_prereg_0_24_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNINEHM6_21_LC_17_7_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNINEHM6_21_LC_17_7_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNINEHM6_21_LC_17_7_6 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNINEHM6_21_LC_17_7_6  (
            .in0(N__72748),
            .in1(N__68350),
            .in2(N__68329),
            .in3(N__68326),
            .lcout(\pid_side.error_d_reg_prev_esr_RNINEHM6Z0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIRLKM6_21_LC_17_7_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIRLKM6_21_LC_17_7_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIRLKM6_21_LC_17_7_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIRLKM6_21_LC_17_7_7  (
            .in0(N__72579),
            .in1(N__72750),
            .in2(N__72730),
            .in3(N__72749),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIRLKM6Z0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIO2HL1_0_21_LC_17_8_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIO2HL1_0_21_LC_17_8_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIO2HL1_0_21_LC_17_8_0 .LUT_INIT=16'b0001100011100111;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIO2HL1_0_21_LC_17_8_0  (
            .in0(N__91377),
            .in1(N__91641),
            .in2(N__72927),
            .in3(N__68175),
            .lcout(\pid_side.un1_pid_prereg_0_17 ),
            .ltout(\pid_side.un1_pid_prereg_0_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIOUVL6_21_LC_17_8_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIOUVL6_21_LC_17_8_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIOUVL6_21_LC_17_8_1 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIOUVL6_21_LC_17_8_1  (
            .in0(N__68293),
            .in1(N__68281),
            .in2(N__68266),
            .in3(N__68141),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIOUVL6Z0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIMVFL1_21_LC_17_8_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIMVFL1_21_LC_17_8_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIMVFL1_21_LC_17_8_2 .LUT_INIT=16'b1110111100001000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIMVFL1_21_LC_17_8_2  (
            .in0(N__91376),
            .in1(N__91640),
            .in2(N__72926),
            .in3(N__68252),
            .lcout(\pid_side.un1_pid_prereg_0_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNISR7K9_16_LC_17_8_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNISR7K9_16_LC_17_8_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNISR7K9_16_LC_17_8_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNISR7K9_16_LC_17_8_3  (
            .in0(N__68224),
            .in1(N__68118),
            .in2(N__68206),
            .in3(N__68085),
            .lcout(\pid_side.error_d_reg_prev_esr_RNISR7K9Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIO2HL1_21_LC_17_8_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIO2HL1_21_LC_17_8_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIO2HL1_21_LC_17_8_4 .LUT_INIT=16'b1110111100001000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIO2HL1_21_LC_17_8_4  (
            .in0(N__91375),
            .in1(N__91639),
            .in2(N__72925),
            .in3(N__68176),
            .lcout(\pid_side.un1_pid_prereg_0_18 ),
            .ltout(\pid_side.un1_pid_prereg_0_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI0B4M6_21_LC_17_8_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI0B4M6_21_LC_17_8_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI0B4M6_21_LC_17_8_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI0B4M6_21_LC_17_8_5  (
            .in0(N__68155),
            .in1(N__68142),
            .in2(N__68128),
            .in3(N__72630),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI0B4M6Z0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIOVFK9_17_LC_17_8_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIOVFK9_17_LC_17_8_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIOVFK9_17_LC_17_8_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIOVFK9_17_LC_17_8_6  (
            .in0(N__68119),
            .in1(N__68100),
            .in2(N__68089),
            .in3(N__68064),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIOVFK9Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNII83B3_21_LC_17_8_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNII83B3_21_LC_17_8_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNII83B3_21_LC_17_8_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNII83B3_21_LC_17_8_7  (
            .in0(_gnd_net_),
            .in1(N__68436),
            .in2(_gnd_net_),
            .in3(N__72629),
            .lcout(\pid_side.error_d_reg_prev_esr_RNII83B3Z0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNI4O091_0_10_LC_17_9_0 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNI4O091_0_10_LC_17_9_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNI4O091_0_10_LC_17_9_0 .LUT_INIT=16'b1000111011001111;
    LogicCell40 \pid_side.error_p_reg_esr_RNI4O091_0_10_LC_17_9_0  (
            .in0(N__79222),
            .in1(N__72989),
            .in2(N__73033),
            .in3(N__73097),
            .lcout(),
            .ltout(\pid_side.error_p_reg_esr_RNI4O091_0Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIV62K2_10_LC_17_9_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIV62K2_10_LC_17_9_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIV62K2_10_LC_17_9_1 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIV62K2_10_LC_17_9_1  (
            .in0(_gnd_net_),
            .in1(N__73073),
            .in2(N__68413),
            .in3(N__68407),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIV62K2Z0Z_10 ),
            .ltout(\pid_side.error_d_reg_prev_esr_RNIV62K2Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNID3GT3_0_10_LC_17_9_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNID3GT3_0_10_LC_17_9_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNID3GT3_0_10_LC_17_9_2 .LUT_INIT=16'b1011010001001011;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNID3GT3_0_10_LC_17_9_2  (
            .in0(N__73029),
            .in1(N__73077),
            .in2(N__68410),
            .in3(N__82341),
            .lcout(\pid_side.error_d_reg_prev_esr_RNID3GT3_0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNI4O091_10_LC_17_9_3 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNI4O091_10_LC_17_9_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNI4O091_10_LC_17_9_3 .LUT_INIT=16'b1111110011010100;
    LogicCell40 \pid_side.error_p_reg_esr_RNI4O091_10_LC_17_9_3  (
            .in0(N__73096),
            .in1(N__73025),
            .in2(N__72991),
            .in3(N__79221),
            .lcout(\pid_side.error_p_reg_esr_RNI4O091Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNI80KL2_12_LC_17_9_4 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNI80KL2_12_LC_17_9_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNI80KL2_12_LC_17_9_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_side.error_p_reg_esr_RNI80KL2_12_LC_17_9_4  (
            .in0(_gnd_net_),
            .in1(N__68622),
            .in2(_gnd_net_),
            .in3(N__68369),
            .lcout(),
            .ltout(\pid_side.un1_pid_prereg_153_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNII28CB_10_LC_17_9_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNII28CB_10_LC_17_9_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNII28CB_10_LC_17_9_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNII28CB_10_LC_17_9_5  (
            .in0(N__72525),
            .in1(N__72568),
            .in2(N__68401),
            .in3(N__68380),
            .lcout(\pid_side.error_d_reg_prev_esr_RNII28CBZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNID3GT3_10_LC_17_9_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNID3GT3_10_LC_17_9_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNID3GT3_10_LC_17_9_6 .LUT_INIT=16'b1110111110001100;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNID3GT3_10_LC_17_9_6  (
            .in0(N__73030),
            .in1(N__82342),
            .in2(N__73078),
            .in3(N__68386),
            .lcout(\pid_side.error_d_reg_prev_esr_RNID3GT3Z0Z_10 ),
            .ltout(\pid_side.error_d_reg_prev_esr_RNID3GT3Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIUOPVA_10_LC_17_9_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIUOPVA_10_LC_17_9_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIUOPVA_10_LC_17_9_7 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIUOPVA_10_LC_17_9_7  (
            .in0(N__68370),
            .in1(N__68649),
            .in2(N__68626),
            .in3(N__68623),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIUOPVAZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIQVAP2_12_LC_17_10_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIQVAP2_12_LC_17_10_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIQVAP2_12_LC_17_10_0 .LUT_INIT=16'b1101000011011101;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIQVAP2_12_LC_17_10_0  (
            .in0(N__79452),
            .in1(N__91247),
            .in2(N__68503),
            .in3(N__68569),
            .lcout(),
            .ltout(\pid_side.un1_pid_prereg_167_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI59QR8_12_LC_17_10_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI59QR8_12_LC_17_10_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI59QR8_12_LC_17_10_1 .LUT_INIT=16'b1110111111100000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI59QR8_12_LC_17_10_1  (
            .in0(N__68518),
            .in1(N__68484),
            .in2(N__68596),
            .in3(N__68458),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI59QR8Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIL0VP1_0_12_LC_17_10_2 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIL0VP1_0_12_LC_17_10_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIL0VP1_0_12_LC_17_10_2 .LUT_INIT=16'b0000110001001101;
    LogicCell40 \pid_side.error_p_reg_esr_RNIL0VP1_0_12_LC_17_10_2  (
            .in0(N__68562),
            .in1(N__69657),
            .in2(N__90978),
            .in3(N__82403),
            .lcout(\pid_side.un1_pid_prereg_167_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_fast_esr_RNIPEC11_12_LC_17_10_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_fast_esr_RNIPEC11_12_LC_17_10_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_fast_esr_RNIPEC11_12_LC_17_10_3 .LUT_INIT=16'b1101111001001000;
    LogicCell40 \pid_side.error_d_reg_fast_esr_RNIPEC11_12_LC_17_10_3  (
            .in0(N__79326),
            .in1(N__90968),
            .in2(N__76226),
            .in3(N__68561),
            .lcout(),
            .ltout(\pid_side.error_d_reg_fast_esr_RNIPEC11Z0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_fast_esr_RNIEIJH2_12_LC_17_10_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_fast_esr_RNIEIJH2_12_LC_17_10_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_fast_esr_RNIEIJH2_12_LC_17_10_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \pid_side.error_d_reg_fast_esr_RNIEIJH2_12_LC_17_10_4  (
            .in0(_gnd_net_),
            .in1(N__68524),
            .in2(N__68548),
            .in3(N__82402),
            .lcout(\pid_side.error_d_reg_fast_esr_RNIEIJH2Z0Z_12 ),
            .ltout(\pid_side.error_d_reg_fast_esr_RNIEIJH2Z0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIJHVG3_12_LC_17_10_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIJHVG3_12_LC_17_10_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIJHVG3_12_LC_17_10_5 .LUT_INIT=16'b1001011011000011;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIJHVG3_12_LC_17_10_5  (
            .in0(N__91248),
            .in1(N__68502),
            .in2(N__68545),
            .in3(N__79453),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIJHVG3Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_fast_esr_RNIPHKN_12_LC_17_10_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_fast_esr_RNIPHKN_12_LC_17_10_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_fast_esr_RNIPHKN_12_LC_17_10_6 .LUT_INIT=16'b1011101111101110;
    LogicCell40 \pid_side.error_d_reg_fast_esr_RNIPHKN_12_LC_17_10_6  (
            .in0(N__90967),
            .in1(N__76216),
            .in2(_gnd_net_),
            .in3(N__79325),
            .lcout(\pid_side.error_d_reg_fast_esr_RNIPHKNZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI4M9H4_14_LC_17_10_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI4M9H4_14_LC_17_10_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI4M9H4_14_LC_17_10_7 .LUT_INIT=16'b1110100010100000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI4M9H4_14_LC_17_10_7  (
            .in0(N__68517),
            .in1(N__68498),
            .in2(N__68485),
            .in3(N__68464),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI4M9H4Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_2_13_LC_17_11_0 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_2_13_LC_17_11_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_2_13_LC_17_11_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_2_13_LC_17_11_0  (
            .in0(N__84256),
            .in1(N__87138),
            .in2(N__84833),
            .in3(N__69583),
            .lcout(\pid_front.error_i_reg_9_rn_2_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_ki_esr_4_LC_17_11_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_esr_4_LC_17_11_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_esr_4_LC_17_11_1 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_esr_4_LC_17_11_1  (
            .in0(_gnd_net_),
            .in1(N__88860),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(xy_ki_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94170),
            .ce(N__83905),
            .sr(N__86429));
    defparam \Commands_frame_decoder.source_xy_ki_esr_7_LC_17_11_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_esr_7_LC_17_11_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_esr_7_LC_17_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_esr_7_LC_17_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__92124),
            .lcout(xy_ki_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94170),
            .ce(N__83905),
            .sr(N__86429));
    defparam \Commands_frame_decoder.source_xy_ki_esr_5_LC_17_11_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_esr_5_LC_17_11_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_esr_5_LC_17_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_esr_5_LC_17_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88701),
            .lcout(xy_ki_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94170),
            .ce(N__83905),
            .sr(N__86429));
    defparam \Commands_frame_decoder.source_xy_ki_esr_6_LC_17_11_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_esr_6_LC_17_11_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_esr_6_LC_17_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_esr_6_LC_17_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88510),
            .lcout(xy_ki_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94170),
            .ce(N__83905),
            .sr(N__86429));
    defparam \pid_side.m78_0_a2_4_LC_17_11_5 .C_ON=1'b0;
    defparam \pid_side.m78_0_a2_4_LC_17_11_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.m78_0_a2_4_LC_17_11_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_side.m78_0_a2_4_LC_17_11_5  (
            .in0(N__70001),
            .in1(N__68699),
            .in2(N__70057),
            .in3(N__84255),
            .lcout(pid_side_N_490),
            .ltout(pid_side_N_490_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_4_11_LC_17_11_6 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_4_11_LC_17_11_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_4_11_LC_17_11_6 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_4_11_LC_17_11_6  (
            .in0(N__87418),
            .in1(N__78503),
            .in2(N__68683),
            .in3(N__80213),
            .lcout(),
            .ltout(\pid_side.m78_0_a2_sx_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_3_11_LC_17_11_7 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_3_11_LC_17_11_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_3_11_LC_17_11_7 .LUT_INIT=16'b0000111000000100;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_3_11_LC_17_11_7  (
            .in0(N__89794),
            .in1(N__85938),
            .in2(N__68680),
            .in3(N__81648),
            .lcout(\pid_side.N_394 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_11_LC_17_12_0 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_11_LC_17_12_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_11_LC_17_12_0 .LUT_INIT=16'b1110101010101010;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_11_LC_17_12_0  (
            .in0(N__68764),
            .in1(N__74962),
            .in2(N__83375),
            .in3(N__68773),
            .lcout(),
            .ltout(\pid_side.m78_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_11_LC_17_12_1 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_11_LC_17_12_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_11_LC_17_12_1 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \pid_side.error_i_reg_esr_11_LC_17_12_1  (
            .in0(N__68671),
            .in1(N__68797),
            .in2(N__68791),
            .in3(N__77029),
            .lcout(\pid_side.error_i_regZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94185),
            .ce(N__86760),
            .sr(N__86419));
    defparam \pid_side.error_cry_2_0_c_RNIEAJ82_LC_17_12_2 .C_ON=1'b0;
    defparam \pid_side.error_cry_2_0_c_RNIEAJ82_LC_17_12_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_2_0_c_RNIEAJ82_LC_17_12_2 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \pid_side.error_cry_2_0_c_RNIEAJ82_LC_17_12_2  (
            .in0(N__82685),
            .in1(N__82850),
            .in2(N__89113),
            .in3(N__83636),
            .lcout(\pid_side.N_626 ),
            .ltout(\pid_side.N_626_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_3_c_RNI8N5S3_LC_17_12_3 .C_ON=1'b0;
    defparam \pid_side.error_cry_3_c_RNI8N5S3_LC_17_12_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_3_c_RNI8N5S3_LC_17_12_3 .LUT_INIT=16'b1111001000000000;
    LogicCell40 \pid_side.error_cry_3_c_RNI8N5S3_LC_17_12_3  (
            .in0(N__77224),
            .in1(N__87775),
            .in2(N__68767),
            .in3(N__83476),
            .lcout(\pid_side.N_576 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_2_11_LC_17_12_4 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_2_11_LC_17_12_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_2_11_LC_17_12_4 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_2_11_LC_17_12_4  (
            .in0(N__87776),
            .in1(N__84092),
            .in2(N__83374),
            .in3(N__76648),
            .lcout(\pid_side.N_398 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_3_c_RNI0N8Q2_LC_17_12_5 .C_ON=1'b0;
    defparam \pid_side.error_cry_3_c_RNI0N8Q2_LC_17_12_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_3_c_RNI0N8Q2_LC_17_12_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \pid_side.error_cry_3_c_RNI0N8Q2_LC_17_12_5  (
            .in0(N__77223),
            .in1(N__85128),
            .in2(_gnd_net_),
            .in3(N__84922),
            .lcout(\pid_side.N_161 ),
            .ltout(\pid_side.N_161_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_3_c_RNI96FF3_LC_17_12_6 .C_ON=1'b0;
    defparam \pid_side.error_cry_3_c_RNI96FF3_LC_17_12_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_3_c_RNI96FF3_LC_17_12_6 .LUT_INIT=16'b0011000000000000;
    LogicCell40 \pid_side.error_cry_3_c_RNI96FF3_LC_17_12_6  (
            .in0(_gnd_net_),
            .in1(N__84091),
            .in2(N__68758),
            .in3(N__76820),
            .lcout(\pid_side.m13_2_03_4_i_0_o2_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_10_c_RNII20I1_LC_17_13_0 .C_ON=1'b0;
    defparam \pid_side.error_cry_10_c_RNII20I1_LC_17_13_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_10_c_RNII20I1_LC_17_13_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \pid_side.error_cry_10_c_RNII20I1_LC_17_13_0  (
            .in0(_gnd_net_),
            .in1(N__84768),
            .in2(_gnd_net_),
            .in3(N__85919),
            .lcout(\pid_side.N_594 ),
            .ltout(\pid_side.N_594_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_2_13_LC_17_13_1 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_2_13_LC_17_13_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_2_13_LC_17_13_1 .LUT_INIT=16'b0001010100000000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_2_13_LC_17_13_1  (
            .in0(N__84491),
            .in1(N__87777),
            .in2(N__68734),
            .in3(N__87140),
            .lcout(),
            .ltout(\pid_side.error_i_reg_9_sn_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_13_LC_17_13_2 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_13_LC_17_13_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_13_LC_17_13_2 .LUT_INIT=16'b0001111100010000;
    LogicCell40 \pid_side.error_i_reg_esr_13_LC_17_13_2  (
            .in0(N__77104),
            .in1(N__77011),
            .in2(N__68731),
            .in3(N__68833),
            .lcout(\pid_side.error_i_regZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94197),
            .ce(N__86782),
            .sr(N__86408));
    defparam \pid_side.error_i_reg_esr_17_LC_17_13_3 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_17_LC_17_13_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_17_LC_17_13_3 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \pid_side.error_i_reg_esr_17_LC_17_13_3  (
            .in0(N__84492),
            .in1(N__68878),
            .in2(N__87128),
            .in3(N__73192),
            .lcout(\pid_side.error_i_regZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94197),
            .ce(N__86782),
            .sr(N__86408));
    defparam \pid_side.error_i_reg_esr_RNO_0_12_LC_17_13_4 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_12_LC_17_13_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_12_LC_17_13_4 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_12_LC_17_13_4  (
            .in0(N__80936),
            .in1(N__84770),
            .in2(N__87417),
            .in3(N__89828),
            .lcout(),
            .ltout(\pid_side.m0_2_03_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_12_LC_17_13_5 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_12_LC_17_13_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_12_LC_17_13_5 .LUT_INIT=16'b1100000001000100;
    LogicCell40 \pid_side.error_i_reg_esr_12_LC_17_13_5  (
            .in0(N__68860),
            .in1(N__87141),
            .in2(N__68854),
            .in3(N__84404),
            .lcout(\pid_side.error_i_regZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94197),
            .ce(N__86782),
            .sr(N__86408));
    defparam \pid_side.error_cry_0_c_RNI4F3S_LC_17_13_6 .C_ON=1'b0;
    defparam \pid_side.error_cry_0_c_RNI4F3S_LC_17_13_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_c_RNI4F3S_LC_17_13_6 .LUT_INIT=16'b0000101100001000;
    LogicCell40 \pid_side.error_cry_0_c_RNI4F3S_LC_17_13_6  (
            .in0(N__80935),
            .in1(N__83008),
            .in2(N__83132),
            .in3(N__81009),
            .lcout(\pid_side.m1_0_03 ),
            .ltout(\pid_side.m1_0_03_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_1_13_LC_17_13_7 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_1_13_LC_17_13_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_1_13_LC_17_13_7 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_1_13_LC_17_13_7  (
            .in0(N__84769),
            .in1(N__87139),
            .in2(N__68836),
            .in3(N__84403),
            .lcout(\pid_side.error_i_reg_9_rn_1_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_3_c_RNIQD011_LC_17_14_0 .C_ON=1'b0;
    defparam \pid_side.error_cry_3_c_RNIQD011_LC_17_14_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_3_c_RNIQD011_LC_17_14_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \pid_side.error_cry_3_c_RNIQD011_LC_17_14_0  (
            .in0(N__82265),
            .in1(N__77222),
            .in2(_gnd_net_),
            .in3(N__80866),
            .lcout(\pid_side.N_232 ),
            .ltout(\pid_side.N_232_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_3_c_RNI32EI1_LC_17_14_1 .C_ON=1'b0;
    defparam \pid_side.error_cry_3_c_RNI32EI1_LC_17_14_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_3_c_RNI32EI1_LC_17_14_1 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \pid_side.error_cry_3_c_RNI32EI1_LC_17_14_1  (
            .in0(_gnd_net_),
            .in1(N__89097),
            .in2(N__68824),
            .in3(N__83477),
            .lcout(\pid_side.N_549 ),
            .ltout(\pid_side.N_549_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_6_LC_17_14_2 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_6_LC_17_14_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_6_LC_17_14_2 .LUT_INIT=16'b1111110011110000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_6_LC_17_14_2  (
            .in0(_gnd_net_),
            .in1(N__69482),
            .in2(N__68821),
            .in3(N__69514),
            .lcout(),
            .ltout(\pid_side.error_i_reg_esr_RNO_0_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_6_LC_17_14_3 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_6_LC_17_14_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_6_LC_17_14_3 .LUT_INIT=16'b1010101010100000;
    LogicCell40 \pid_side.error_i_reg_esr_6_LC_17_14_3  (
            .in0(N__83350),
            .in1(_gnd_net_),
            .in2(N__68818),
            .in3(N__73687),
            .lcout(\pid_side.error_i_regZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94214),
            .ce(N__86774),
            .sr(N__86399));
    defparam \pid_side.error_cry_3_0_c_RNINVTD2_LC_17_14_4 .C_ON=1'b0;
    defparam \pid_side.error_cry_3_0_c_RNINVTD2_LC_17_14_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_3_0_c_RNINVTD2_LC_17_14_4 .LUT_INIT=16'b0100011100000000;
    LogicCell40 \pid_side.error_cry_3_0_c_RNINVTD2_LC_17_14_4  (
            .in0(N__83637),
            .in1(N__82742),
            .in2(N__85246),
            .in3(N__74942),
            .lcout(\pid_side.N_580 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_3_0_c_RNIO3R61_LC_17_14_5 .C_ON=1'b0;
    defparam \pid_side.error_cry_3_0_c_RNIO3R61_LC_17_14_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_3_0_c_RNIO3R61_LC_17_14_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \pid_side.error_cry_3_0_c_RNIO3R61_LC_17_14_5  (
            .in0(N__78498),
            .in1(N__80948),
            .in2(_gnd_net_),
            .in3(N__85233),
            .lcout(\pid_side.N_156 ),
            .ltout(\pid_side.N_156_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_2_0_c_RNIMM2O2_LC_17_14_6 .C_ON=1'b0;
    defparam \pid_side.error_cry_2_0_c_RNIMM2O2_LC_17_14_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_2_0_c_RNIMM2O2_LC_17_14_6 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \pid_side.error_cry_2_0_c_RNIMM2O2_LC_17_14_6  (
            .in0(N__83638),
            .in1(N__85084),
            .in2(N__69517),
            .in3(N__82743),
            .lcout(\pid_side.N_182 ),
            .ltout(\pid_side.N_182_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_1_22_LC_17_14_7 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_1_22_LC_17_14_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_1_22_LC_17_14_7 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_1_22_LC_17_14_7  (
            .in0(N__69481),
            .in1(N__69451),
            .in2(N__69445),
            .in3(N__73686),
            .lcout(\pid_side.m10_2_03_3_i_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_5_LC_17_15_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_5_LC_17_15_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_5_LC_17_15_0 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \Commands_frame_decoder.state_5_LC_17_15_0  (
            .in0(N__69342),
            .in1(N__69442),
            .in2(_gnd_net_),
            .in3(N__69416),
            .lcout(\Commands_frame_decoder.stateZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94230),
            .ce(),
            .sr(N__86389));
    defparam \dron_frame_decoder_1.state_7_LC_17_15_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_7_LC_17_15_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_7_LC_17_15_1 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \dron_frame_decoder_1.state_7_LC_17_15_1  (
            .in0(N__69222),
            .in1(N__69322),
            .in2(_gnd_net_),
            .in3(N__69298),
            .lcout(\dron_frame_decoder_1.stateZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94230),
            .ce(),
            .sr(N__86389));
    defparam \pid_alt.state_0_LC_17_15_2 .C_ON=1'b0;
    defparam \pid_alt.state_0_LC_17_15_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.state_0_LC_17_15_2 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \pid_alt.state_0_LC_17_15_2  (
            .in0(N__69045),
            .in1(N__69198),
            .in2(_gnd_net_),
            .in3(N__68912),
            .lcout(\pid_alt.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94230),
            .ce(),
            .sr(N__86389));
    defparam \pid_alt.state_1_LC_17_15_3 .C_ON=1'b0;
    defparam \pid_alt.state_1_LC_17_15_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.state_1_LC_17_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.state_1_LC_17_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69046),
            .lcout(\pid_alt.N_72_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94230),
            .ce(),
            .sr(N__86389));
    defparam \pid_front.error_p_reg_esr_RNICMVCG_14_LC_17_15_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNICMVCG_14_LC_17_15_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNICMVCG_14_LC_17_15_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_front.error_p_reg_esr_RNICMVCG_14_LC_17_15_4  (
            .in0(_gnd_net_),
            .in1(N__71091),
            .in2(_gnd_net_),
            .in3(N__71563),
            .lcout(\pid_front.error_p_reg_esr_RNICMVCGZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_fast_esr_RNIGBTF_12_LC_17_15_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_fast_esr_RNIGBTF_12_LC_17_15_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_fast_esr_RNIGBTF_12_LC_17_15_5 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \pid_side.error_d_reg_fast_esr_RNIGBTF_12_LC_17_15_5  (
            .in0(N__76227),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79327),
            .lcout(\pid_side.N_2601_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIMERG_1_12_LC_17_15_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIMERG_1_12_LC_17_15_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIMERG_1_12_LC_17_15_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIMERG_1_12_LC_17_15_6  (
            .in0(_gnd_net_),
            .in1(N__79468),
            .in2(_gnd_net_),
            .in3(N__91249),
            .lcout(\pid_side.g1_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNITU3P4_0_10_LC_17_15_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNITU3P4_0_10_LC_17_15_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNITU3P4_0_10_LC_17_15_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNITU3P4_0_10_LC_17_15_7  (
            .in0(_gnd_net_),
            .in1(N__72567),
            .in2(_gnd_net_),
            .in3(N__72526),
            .lcout(\pid_side.error_d_reg_prev_esr_RNITU3P4_0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_1_c_RNITUNK1_LC_17_16_0 .C_ON=1'b0;
    defparam \pid_front.error_cry_1_c_RNITUNK1_LC_17_16_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_1_c_RNITUNK1_LC_17_16_0 .LUT_INIT=16'b0010000000101010;
    LogicCell40 \pid_front.error_cry_1_c_RNITUNK1_LC_17_16_0  (
            .in0(N__83009),
            .in1(N__80004),
            .in2(N__90649),
            .in3(N__79903),
            .lcout(\pid_front.N_429 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_0_c_RNIT3D41_LC_17_16_1 .C_ON=1'b0;
    defparam \pid_front.error_cry_0_0_c_RNIT3D41_LC_17_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_0_c_RNIT3D41_LC_17_16_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \pid_front.error_cry_0_0_c_RNIT3D41_LC_17_16_1  (
            .in0(N__83011),
            .in1(N__90600),
            .in2(_gnd_net_),
            .in3(N__77968),
            .lcout(),
            .ltout(\pid_front.N_332_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_2_c_RNID2UK3_LC_17_16_2 .C_ON=1'b0;
    defparam \pid_front.error_cry_2_c_RNID2UK3_LC_17_16_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_2_c_RNID2UK3_LC_17_16_2 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \pid_front.error_cry_2_c_RNID2UK3_LC_17_16_2  (
            .in0(N__85748),
            .in1(N__69637),
            .in2(N__69631),
            .in3(N__74081),
            .lcout(\pid_front.N_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_0_17_LC_17_16_3 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_17_LC_17_16_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_17_LC_17_16_3 .LUT_INIT=16'b0000000100010001;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_17_LC_17_16_3  (
            .in0(N__74542),
            .in1(N__77047),
            .in2(N__87443),
            .in3(N__69628),
            .lcout(),
            .ltout(\pid_front.error_i_reg_esr_RNO_0Z0Z_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_17_LC_17_16_4 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_17_LC_17_16_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_17_LC_17_16_4 .LUT_INIT=16'b1010100000100000;
    LogicCell40 \pid_front.error_i_reg_esr_17_LC_17_16_4  (
            .in0(N__87104),
            .in1(N__84413),
            .in2(N__69622),
            .in3(N__69532),
            .lcout(\pid_front.error_i_regZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94246),
            .ce(N__78137),
            .sr(N__86381));
    defparam \pid_front.error_i_reg_esr_RNO_1_17_LC_17_16_5 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_1_17_LC_17_16_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_1_17_LC_17_16_5 .LUT_INIT=16'b0101000100000001;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_1_17_LC_17_16_5  (
            .in0(N__89338),
            .in1(N__69594),
            .in2(N__84187),
            .in3(N__69581),
            .lcout(\pid_front.error_i_reg_esr_RNO_1Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_2_0_c_RNI8A562_LC_17_17_0 .C_ON=1'b0;
    defparam \pid_front.error_cry_2_0_c_RNI8A562_LC_17_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_2_0_c_RNI8A562_LC_17_17_0 .LUT_INIT=16'b0010000001110000;
    LogicCell40 \pid_front.error_cry_2_0_c_RNI8A562_LC_17_17_0  (
            .in0(N__83010),
            .in1(N__77743),
            .in2(N__74967),
            .in3(N__74858),
            .lcout(\pid_front.N_580 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_2_12_LC_17_17_1 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_2_12_LC_17_17_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_2_12_LC_17_17_1 .LUT_INIT=16'b1000000010001010;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_2_12_LC_17_17_1  (
            .in0(N__89028),
            .in1(N__73483),
            .in2(N__89815),
            .in3(N__78205),
            .lcout(),
            .ltout(\pid_front.m16_2_03_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_1_12_LC_17_17_2 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_1_12_LC_17_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_1_12_LC_17_17_2 .LUT_INIT=16'b1111010111110100;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_1_12_LC_17_17_2  (
            .in0(N__87434),
            .in1(N__74372),
            .in2(N__69745),
            .in3(N__69675),
            .lcout(),
            .ltout(\pid_front.m16_2_03_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_12_LC_17_17_3 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_12_LC_17_17_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_12_LC_17_17_3 .LUT_INIT=16'b1000100000001100;
    LogicCell40 \pid_front.error_i_reg_esr_12_LC_17_17_3  (
            .in0(N__84595),
            .in1(N__86936),
            .in2(N__69742),
            .in3(N__84414),
            .lcout(\pid_front.error_i_regZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94264),
            .ce(N__78131),
            .sr(N__86375));
    defparam \pid_front.error_i_reg_esr_RNO_1_14_LC_17_17_4 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_1_14_LC_17_17_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_1_14_LC_17_17_4 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_1_14_LC_17_17_4  (
            .in0(N__87435),
            .in1(N__69676),
            .in2(N__69763),
            .in3(N__74373),
            .lcout(),
            .ltout(\pid_front.m18_2_03_4_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_14_LC_17_17_5 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_14_LC_17_17_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_14_LC_17_17_5 .LUT_INIT=16'b1000100000001000;
    LogicCell40 \pid_front.error_i_reg_esr_14_LC_17_17_5  (
            .in0(N__69769),
            .in1(N__86937),
            .in2(N__69724),
            .in3(N__84415),
            .lcout(\pid_front.error_i_regZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94264),
            .ce(N__78131),
            .sr(N__86375));
    defparam \pid_front.error_cry_2_0_c_RNITT5E5_LC_17_17_6 .C_ON=1'b0;
    defparam \pid_front.error_cry_2_0_c_RNITT5E5_LC_17_17_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_2_0_c_RNITT5E5_LC_17_17_6 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \pid_front.error_cry_2_0_c_RNITT5E5_LC_17_17_6  (
            .in0(N__89576),
            .in1(N__69709),
            .in2(_gnd_net_),
            .in3(N__69701),
            .lcout(\pid_front.N_263 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_c_RNIEOA53_LC_17_18_0 .C_ON=1'b0;
    defparam \pid_front.error_cry_0_c_RNIEOA53_LC_17_18_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_c_RNIEOA53_LC_17_18_0 .LUT_INIT=16'b1111111111001110;
    LogicCell40 \pid_front.error_cry_0_c_RNIEOA53_LC_17_18_0  (
            .in0(N__74146),
            .in1(N__73653),
            .in2(N__87774),
            .in3(N__79782),
            .lcout(\pid_front.N_54_i_1 ),
            .ltout(\pid_front.N_54_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_5_16_LC_17_18_1 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_5_16_LC_17_18_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_5_16_LC_17_18_1 .LUT_INIT=16'b0000000010111000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_5_16_LC_17_18_1  (
            .in0(N__82296),
            .in1(N__84181),
            .in2(N__69661),
            .in3(N__89307),
            .lcout(),
            .ltout(\pid_front.error_i_reg_esr_RNO_5Z0Z_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_1_16_LC_17_18_2 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_1_16_LC_17_18_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_1_16_LC_17_18_2 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_1_16_LC_17_18_2  (
            .in0(N__87030),
            .in1(_gnd_net_),
            .in2(N__69832),
            .in3(N__84487),
            .lcout(),
            .ltout(\pid_front.error_i_reg_9_rn_0_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_16_LC_17_18_3 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_16_LC_17_18_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_16_LC_17_18_3 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \pid_front.error_i_reg_esr_16_LC_17_18_3  (
            .in0(N__69982),
            .in1(N__74380),
            .in2(N__69829),
            .in3(N__69811),
            .lcout(\pid_front.error_i_regZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94282),
            .ce(N__78142),
            .sr(N__86370));
    defparam \pid_front.error_i_reg_esr_RNO_2_16_LC_17_18_4 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_2_16_LC_17_18_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_2_16_LC_17_18_4 .LUT_INIT=16'b0001000001010000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_2_16_LC_17_18_4  (
            .in0(N__84402),
            .in1(N__85750),
            .in2(N__87089),
            .in3(N__69793),
            .lcout(\pid_front.error_i_reg_9_sn_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_5_c_RNIOO142_LC_17_18_5 .C_ON=1'b0;
    defparam \pid_front.error_cry_5_c_RNIOO142_LC_17_18_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_5_c_RNIOO142_LC_17_18_5 .LUT_INIT=16'b0000010011110100;
    LogicCell40 \pid_front.error_cry_5_c_RNIOO142_LC_17_18_5  (
            .in0(N__78412),
            .in1(N__89306),
            .in2(N__89592),
            .in3(N__69805),
            .lcout(\pid_front.N_259 ),
            .ltout(\pid_front.N_259_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_0_14_LC_17_18_6 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_14_LC_17_18_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_14_LC_17_18_6 .LUT_INIT=16'b0001010110111111;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_14_LC_17_18_6  (
            .in0(N__84401),
            .in1(N__81259),
            .in2(N__69787),
            .in3(N__69784),
            .lcout(\pid_front.error_i_reg_9_1_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_3_14_LC_17_19_0 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_3_14_LC_17_19_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_3_14_LC_17_19_0 .LUT_INIT=16'b1000100010101000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_3_14_LC_17_19_0  (
            .in0(N__76896),
            .in1(N__69974),
            .in2(N__83522),
            .in3(N__73893),
            .lcout(\pid_front.N_454 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_4_c_RNIMV991_LC_17_19_1 .C_ON=1'b0;
    defparam \pid_front.error_cry_4_c_RNIMV991_LC_17_19_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_4_c_RNIMV991_LC_17_19_1 .LUT_INIT=16'b0000001010100010;
    LogicCell40 \pid_front.error_cry_4_c_RNIMV991_LC_17_19_1  (
            .in0(N__90223),
            .in1(N__73769),
            .in2(N__90435),
            .in3(N__77974),
            .lcout(\pid_front.N_515 ),
            .ltout(\pid_front.N_515_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_7_15_LC_17_19_2 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_7_15_LC_17_19_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_7_15_LC_17_19_2 .LUT_INIT=16'b1100000011001000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_7_15_LC_17_19_2  (
            .in0(N__83515),
            .in1(N__85749),
            .in2(N__69751),
            .in3(N__73896),
            .lcout(),
            .ltout(\pid_front.N_450_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_3_15_LC_17_19_3 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_3_15_LC_17_19_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_3_15_LC_17_19_3 .LUT_INIT=16'b1111000011110100;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_3_15_LC_17_19_3  (
            .in0(N__89293),
            .in1(N__81325),
            .in2(N__69748),
            .in3(N__80629),
            .lcout(\pid_front.m19_2_03_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_6_16_LC_17_19_4 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_6_16_LC_17_19_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_6_16_LC_17_19_4 .LUT_INIT=16'b0000110000001110;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_6_16_LC_17_19_4  (
            .in0(N__83514),
            .in1(N__69975),
            .in2(N__87805),
            .in3(N__73894),
            .lcout(),
            .ltout(\pid_front.N_446_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_3_16_LC_17_19_5 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_3_16_LC_17_19_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_3_16_LC_17_19_5 .LUT_INIT=16'b1111000011110001;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_3_16_LC_17_19_5  (
            .in0(N__87428),
            .in1(N__89292),
            .in2(N__69985),
            .in3(N__80630),
            .lcout(\pid_front.m20_2_03_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_5_13_LC_17_19_6 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_5_13_LC_17_19_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_5_13_LC_17_19_6 .LUT_INIT=16'b1000100010101000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_5_13_LC_17_19_6  (
            .in0(N__81324),
            .in1(N__69976),
            .in2(N__83523),
            .in3(N__73895),
            .lcout(),
            .ltout(\pid_front.N_438_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_3_13_LC_17_19_7 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_3_13_LC_17_19_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_3_13_LC_17_19_7 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_3_13_LC_17_19_7  (
            .in0(N__86934),
            .in1(N__84486),
            .in2(N__69964),
            .in3(N__69838),
            .lcout(\pid_front.error_i_reg_9_sn_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNI6EER_0_14_LC_17_20_0 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI6EER_0_14_LC_17_20_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI6EER_0_14_LC_17_20_0 .LUT_INIT=16'b0101111111111111;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNI6EER_0_14_LC_17_20_0  (
            .in0(N__69849),
            .in1(_gnd_net_),
            .in2(N__69931),
            .in3(N__69894),
            .lcout(\pid_front.error_i_acumm_13_i_o2_0_7_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_14_LC_17_20_1 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_14_LC_17_20_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_14_LC_17_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_14_LC_17_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69950),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94313),
            .ce(N__75327),
            .sr(N__86363));
    defparam \pid_front.error_i_acumm_prereg_esr_22_LC_17_20_2 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_22_LC_17_20_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_22_LC_17_20_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_22_LC_17_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69916),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94313),
            .ce(N__75327),
            .sr(N__86363));
    defparam \pid_front.error_i_acumm_prereg_esr_27_LC_17_20_3 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_27_LC_17_20_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_27_LC_17_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_27_LC_17_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69882),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94313),
            .ce(N__75327),
            .sr(N__86363));
    defparam \pid_front.error_i_reg_esr_RNO_6_13_LC_17_20_4 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_6_13_LC_17_20_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_6_13_LC_17_20_4 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_6_13_LC_17_20_4  (
            .in0(N__87773),
            .in1(N__84816),
            .in2(_gnd_net_),
            .in3(N__80681),
            .lcout(\pid_front.N_439 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_4_15_LC_17_20_5 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_4_15_LC_17_20_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_4_15_LC_17_20_5 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_4_15_LC_17_20_5  (
            .in0(N__84815),
            .in1(N__80788),
            .in2(_gnd_net_),
            .in3(N__80773),
            .lcout(\pid_side.N_109 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI0GC61_0_19_LC_17_20_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI0GC61_0_19_LC_17_20_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI0GC61_0_19_LC_17_20_6 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_p_reg_esr_RNI0GC61_0_19_LC_17_20_6  (
            .in0(N__70224),
            .in1(N__70236),
            .in2(_gnd_net_),
            .in3(N__91811),
            .lcout(\pid_front.error_p_reg_esr_RNI0GC61_0Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI0GC61_19_LC_17_20_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI0GC61_19_LC_17_20_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI0GC61_19_LC_17_20_7 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \pid_front.error_p_reg_esr_RNI0GC61_19_LC_17_20_7  (
            .in0(N__91812),
            .in1(_gnd_net_),
            .in2(N__70240),
            .in3(N__70225),
            .lcout(\pid_front.error_p_reg_esr_RNI0GC61Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNIQVBR_10_LC_17_21_0 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIQVBR_10_LC_17_21_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIQVBR_10_LC_17_21_0 .LUT_INIT=16'b0000000001011111;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNIQVBR_10_LC_17_21_0  (
            .in0(N__75101),
            .in1(_gnd_net_),
            .in2(N__75026),
            .in3(N__75670),
            .lcout(),
            .ltout(\pid_front.N_531_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNIR6LR5_28_LC_17_21_1 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIR6LR5_28_LC_17_21_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIR6LR5_28_LC_17_21_1 .LUT_INIT=16'b1110111011101100;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNIR6LR5_28_LC_17_21_1  (
            .in0(N__75964),
            .in1(N__75868),
            .in2(N__70186),
            .in3(N__75056),
            .lcout(\pid_front.N_255 ),
            .ltout(\pid_front.N_255_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_9_LC_17_21_2 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_9_LC_17_21_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_9_LC_17_21_2 .LUT_INIT=16'b0000101000001011;
    LogicCell40 \pid_front.error_i_acumm_9_LC_17_21_2  (
            .in0(N__70174),
            .in1(N__70145),
            .in2(N__70132),
            .in3(N__75965),
            .lcout(\pid_front.error_i_acummZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94329),
            .ce(N__75765),
            .sr(_gnd_net_));
    defparam \pid_front.state_RNI0V2N_1_LC_17_21_3 .C_ON=1'b0;
    defparam \pid_front.state_RNI0V2N_1_LC_17_21_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.state_RNI0V2N_1_LC_17_21_3 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \pid_front.state_RNI0V2N_1_LC_17_21_3  (
            .in0(N__75963),
            .in1(N__70495),
            .in2(_gnd_net_),
            .in3(N__71063),
            .lcout(\pid_front.N_276 ),
            .ltout(\pid_front.N_276_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNIU9HN5_3_LC_17_21_4 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIU9HN5_3_LC_17_21_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIU9HN5_3_LC_17_21_4 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNIU9HN5_3_LC_17_21_4  (
            .in0(N__75057),
            .in1(N__74623),
            .in2(N__70099),
            .in3(N__70411),
            .lcout(\pid_front.N_632 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.state_RNI2NLV1_0_LC_17_21_5 .C_ON=1'b0;
    defparam \pid_front.state_RNI2NLV1_0_LC_17_21_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.state_RNI2NLV1_0_LC_17_21_5 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \pid_front.state_RNI2NLV1_0_LC_17_21_5  (
            .in0(N__70078),
            .in1(N__70061),
            .in2(N__70612),
            .in3(N__70027),
            .lcout(),
            .ltout(\pid_front.N_382_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.state_RNIOKAI2_0_LC_17_21_6 .C_ON=1'b0;
    defparam \pid_front.state_RNIOKAI2_0_LC_17_21_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.state_RNIOKAI2_0_LC_17_21_6 .LUT_INIT=16'b1111101111111010;
    LogicCell40 \pid_front.state_RNIOKAI2_0_LC_17_21_6  (
            .in0(N__71064),
            .in1(N__70610),
            .in2(N__70525),
            .in3(N__70497),
            .lcout(\pid_front.N_64 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNIRU7I_10_LC_17_21_7 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIRU7I_10_LC_17_21_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIRU7I_10_LC_17_21_7 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNIRU7I_10_LC_17_21_7  (
            .in0(_gnd_net_),
            .in1(N__75013),
            .in2(_gnd_net_),
            .in3(N__75100),
            .lcout(\pid_front.N_217 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNILQ6F_9_LC_17_22_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNILQ6F_9_LC_17_22_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNILQ6F_9_LC_17_22_0 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \pid_front.error_p_reg_esr_RNILQ6F_9_LC_17_22_0  (
            .in0(N__78808),
            .in1(N__71344),
            .in2(N__71320),
            .in3(N__71337),
            .lcout(\pid_front.error_p_reg_esr_RNILQ6FZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIQK6U_10_LC_17_22_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIQK6U_10_LC_17_22_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIQK6U_10_LC_17_22_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIQK6U_10_LC_17_22_1  (
            .in0(_gnd_net_),
            .in1(N__70268),
            .in2(_gnd_net_),
            .in3(N__81896),
            .lcout(),
            .ltout(\pid_front.N_2382_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIFM3D1_10_LC_17_22_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIFM3D1_10_LC_17_22_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIFM3D1_10_LC_17_22_2 .LUT_INIT=16'b0101101010010110;
    LogicCell40 \pid_front.error_p_reg_esr_RNIFM3D1_10_LC_17_22_2  (
            .in0(N__70399),
            .in1(N__71362),
            .in2(N__70375),
            .in3(N__78738),
            .lcout(\pid_front.error_p_reg_esr_RNIFM3D1Z0Z_10 ),
            .ltout(\pid_front.error_p_reg_esr_RNIFM3D1Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIS5CU3_9_LC_17_22_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIS5CU3_9_LC_17_22_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIS5CU3_9_LC_17_22_3 .LUT_INIT=16'b1001011010010110;
    LogicCell40 \pid_front.error_p_reg_esr_RNIS5CU3_9_LC_17_22_3  (
            .in0(N__75170),
            .in1(N__70332),
            .in2(N__70372),
            .in3(N__70365),
            .lcout(\pid_front.error_p_reg_esr_RNIS5CU3Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNINU9V7_9_LC_17_22_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNINU9V7_9_LC_17_22_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNINU9V7_9_LC_17_22_4 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_front.error_p_reg_esr_RNINU9V7_9_LC_17_22_4  (
            .in0(N__70333),
            .in1(N__75171),
            .in2(N__70324),
            .in3(N__70303),
            .lcout(\pid_front.error_p_reg_esr_RNINU9V7Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_10_LC_17_22_5 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_10_LC_17_22_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_10_LC_17_22_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_10_LC_17_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81897),
            .lcout(\pid_front.error_d_reg_prevZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94344),
            .ce(N__71785),
            .sr(N__71683));
    defparam \pid_front.error_d_reg_prev_esr_RNIA2O6_9_LC_17_22_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIA2O6_9_LC_17_22_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIA2O6_9_LC_17_22_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIA2O6_9_LC_17_22_6  (
            .in0(_gnd_net_),
            .in1(N__71361),
            .in2(_gnd_net_),
            .in3(N__78737),
            .lcout(\pid_front.N_2376_i ),
            .ltout(\pid_front.N_2376_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNILQ6F_0_9_LC_17_22_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNILQ6F_0_9_LC_17_22_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNILQ6F_0_9_LC_17_22_7 .LUT_INIT=16'b0011110010010110;
    LogicCell40 \pid_front.error_p_reg_esr_RNILQ6F_0_9_LC_17_22_7  (
            .in0(N__71336),
            .in1(N__71316),
            .in2(N__71293),
            .in3(N__78807),
            .lcout(\pid_front.error_p_reg_esr_RNILQ6F_0Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNIBKH41_0_15_LC_17_23_0 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIBKH41_0_15_LC_17_23_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIBKH41_0_15_LC_17_23_0 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNIBKH41_0_15_LC_17_23_0  (
            .in0(N__71193),
            .in1(N__71232),
            .in2(N__71160),
            .in3(N__71265),
            .lcout(\pid_front.error_i_acumm_13_i_o2_0_9_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_15_LC_17_23_1 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_15_LC_17_23_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_15_LC_17_23_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_15_LC_17_23_1  (
            .in0(N__71115),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94359),
            .ce(N__75325),
            .sr(N__86356));
    defparam \pid_front.error_i_acumm_prereg_esr_RNIBKH41_15_LC_17_23_2 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIBKH41_15_LC_17_23_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIBKH41_15_LC_17_23_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNIBKH41_15_LC_17_23_2  (
            .in0(N__71194),
            .in1(N__71233),
            .in2(N__71161),
            .in3(N__71266),
            .lcout(\pid_front.error_i_acumm_13_i_o2_0_9_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_16_LC_17_23_3 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_16_LC_17_23_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_16_LC_17_23_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_16_LC_17_23_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71257),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94359),
            .ce(N__75325),
            .sr(N__86356));
    defparam \pid_front.error_i_acumm_prereg_esr_17_LC_17_23_4 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_17_LC_17_23_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_17_LC_17_23_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_17_LC_17_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71223),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94359),
            .ce(N__75325),
            .sr(N__86356));
    defparam \pid_front.error_i_acumm_prereg_esr_24_LC_17_23_5 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_24_LC_17_23_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_24_LC_17_23_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_24_LC_17_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71185),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94359),
            .ce(N__75325),
            .sr(N__86356));
    defparam \pid_front.error_p_reg_esr_RNIBJ5B3_0_14_LC_17_23_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIBJ5B3_0_14_LC_17_23_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIBJ5B3_0_14_LC_17_23_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_p_reg_esr_RNIBJ5B3_0_14_LC_17_23_6  (
            .in0(N__71142),
            .in1(N__71127),
            .in2(_gnd_net_),
            .in3(N__71114),
            .lcout(\pid_front.error_p_reg_esr_RNIBJ5B3_0Z0Z_14 ),
            .ltout(\pid_front.error_p_reg_esr_RNIBJ5B3_0Z0Z_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI4820U_12_LC_17_23_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI4820U_12_LC_17_23_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI4820U_12_LC_17_23_7 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_front.error_p_reg_esr_RNI4820U_12_LC_17_23_7  (
            .in0(N__71596),
            .in1(_gnd_net_),
            .in2(N__71566),
            .in3(N__71552),
            .lcout(\pid_front.error_p_reg_esr_RNI4820UZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNI18694_0_13_LC_17_24_1 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI18694_0_13_LC_17_24_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI18694_0_13_LC_17_24_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNI18694_0_13_LC_17_24_1  (
            .in0(N__71518),
            .in1(N__71440),
            .in2(N__71512),
            .in3(N__71497),
            .lcout(\pid_front.N_227 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNI18694_13_LC_17_24_3 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI18694_13_LC_17_24_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI18694_13_LC_17_24_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNI18694_13_LC_17_24_3  (
            .in0(N__71485),
            .in1(N__71455),
            .in2(N__71479),
            .in3(N__71464),
            .lcout(\pid_front.N_203 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNI4FJ41_0_19_LC_17_25_0 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI4FJ41_0_19_LC_17_25_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI4FJ41_0_19_LC_17_25_0 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNI4FJ41_0_19_LC_17_25_0  (
            .in0(N__71370),
            .in1(N__71406),
            .in2(N__72105),
            .in3(N__71448),
            .lcout(\pid_front.error_i_acumm_13_i_o2_0_8_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_19_LC_17_25_1 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_19_LC_17_25_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_19_LC_17_25_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_19_LC_17_25_1  (
            .in0(N__72057),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94376),
            .ce(N__75323),
            .sr(N__86352));
    defparam \pid_front.error_i_acumm_prereg_esr_RNI4FJ41_19_LC_17_25_2 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI4FJ41_19_LC_17_25_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI4FJ41_19_LC_17_25_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNI4FJ41_19_LC_17_25_2  (
            .in0(N__71371),
            .in1(N__71407),
            .in2(N__72106),
            .in3(N__71449),
            .lcout(\pid_front.error_i_acumm_13_i_o2_0_8_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_20_LC_17_25_3 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_20_LC_17_25_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_20_LC_17_25_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_20_LC_17_25_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71434),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94376),
            .ce(N__75323),
            .sr(N__86352));
    defparam \pid_front.error_i_acumm_prereg_esr_21_LC_17_25_4 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_21_LC_17_25_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_21_LC_17_25_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_21_LC_17_25_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71398),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94376),
            .ce(N__75323),
            .sr(N__86352));
    defparam \pid_front.error_i_acumm_prereg_esr_23_LC_17_25_5 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_23_LC_17_25_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_23_LC_17_25_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_23_LC_17_25_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72136),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94376),
            .ce(N__75323),
            .sr(N__86352));
    defparam \pid_front.error_p_reg_esr_RNIBOAB3_0_18_LC_17_25_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIBOAB3_0_18_LC_17_25_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIBOAB3_0_18_LC_17_25_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_front.error_p_reg_esr_RNIBOAB3_0_18_LC_17_25_6  (
            .in0(N__76140),
            .in1(_gnd_net_),
            .in2(N__72084),
            .in3(N__72056),
            .lcout(\pid_front.un1_pid_prereg_0_7 ),
            .ltout(\pid_front.un1_pid_prereg_0_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIE7KM6_17_LC_17_25_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIE7KM6_17_LC_17_25_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIE7KM6_17_LC_17_25_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIE7KM6_17_LC_17_25_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__72016),
            .in3(N__72012),
            .lcout(\pid_front.error_p_reg_esr_RNIE7KM6Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_fast_esr_12_LC_17_26_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_fast_esr_12_LC_17_26_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_fast_esr_12_LC_17_26_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_fast_esr_12_LC_17_26_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81859),
            .lcout(\pid_front.error_d_reg_fastZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94384),
            .ce(N__93406),
            .sr(N__93007));
    defparam \pid_front.error_p_reg_esr_RNI8NB61_2_11_LC_17_27_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI8NB61_2_11_LC_17_27_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI8NB61_2_11_LC_17_27_3 .LUT_INIT=16'b0111011100010001;
    LogicCell40 \pid_front.error_p_reg_esr_RNI8NB61_2_11_LC_17_27_3  (
            .in0(N__94588),
            .in1(N__71939),
            .in2(_gnd_net_),
            .in3(N__71844),
            .lcout(),
            .ltout(\pid_front.g0_1_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIJHNC2_12_LC_17_27_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIJHNC2_12_LC_17_27_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIJHNC2_12_LC_17_27_4 .LUT_INIT=16'b1001000011111001;
    LogicCell40 \pid_front.error_p_reg_esr_RNIJHNC2_12_LC_17_27_4  (
            .in0(N__81827),
            .in1(N__78694),
            .in2(N__71917),
            .in3(N__71903),
            .lcout(\pid_front.g0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIUO6U_0_12_LC_17_27_5 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIUO6U_0_12_LC_17_27_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIUO6U_0_12_LC_17_27_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIUO6U_0_12_LC_17_27_5  (
            .in0(_gnd_net_),
            .in1(N__78690),
            .in2(_gnd_net_),
            .in3(N__81826),
            .lcout(\pid_front.N_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_11_LC_17_27_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_11_LC_17_27_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_11_LC_17_27_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_11_LC_17_27_7  (
            .in0(N__94589),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prevZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94389),
            .ce(N__71816),
            .sr(N__71716));
    defparam \pid_side.error_p_reg_esr_RNIFJGD3_6_LC_18_5_0 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIFJGD3_6_LC_18_5_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIFJGD3_6_LC_18_5_0 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_side.error_p_reg_esr_RNIFJGD3_6_LC_18_5_0  (
            .in0(N__72292),
            .in1(N__72286),
            .in2(_gnd_net_),
            .in3(N__72274),
            .lcout(\pid_side.error_p_reg_esr_RNIFJGD3Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNISPEI_6_LC_18_5_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNISPEI_6_LC_18_5_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNISPEI_6_LC_18_5_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNISPEI_6_LC_18_5_1  (
            .in0(_gnd_net_),
            .in1(N__72239),
            .in2(_gnd_net_),
            .in3(N__78553),
            .lcout(),
            .ltout(\pid_side.N_2565_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIIFTC1_6_LC_18_5_2 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIIFTC1_6_LC_18_5_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIIFTC1_6_LC_18_5_2 .LUT_INIT=16'b1010111100101011;
    LogicCell40 \pid_side.error_p_reg_esr_RNIIFTC1_6_LC_18_5_2  (
            .in0(N__90015),
            .in1(N__76272),
            .in2(N__72295),
            .in3(N__78621),
            .lcout(\pid_side.error_p_reg_esr_RNIIFTC1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNINKTC1_0_7_LC_18_5_3 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNINKTC1_0_7_LC_18_5_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNINKTC1_0_7_LC_18_5_3 .LUT_INIT=16'b0101101010010110;
    LogicCell40 \pid_side.error_p_reg_esr_RNINKTC1_0_7_LC_18_5_3  (
            .in0(N__72489),
            .in1(N__72240),
            .in2(N__89971),
            .in3(N__78554),
            .lcout(\pid_side.error_p_reg_esr_RNINKTC1_0Z0Z_7 ),
            .ltout(\pid_side.error_p_reg_esr_RNINKTC1_0Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIFJGD3_0_6_LC_18_5_4 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIFJGD3_0_6_LC_18_5_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIFJGD3_0_6_LC_18_5_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_p_reg_esr_RNIFJGD3_0_6_LC_18_5_4  (
            .in0(_gnd_net_),
            .in1(N__72285),
            .in2(N__72277),
            .in3(N__72273),
            .lcout(\pid_side.error_p_reg_esr_RNIFJGD3_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_6_LC_18_5_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_6_LC_18_5_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_6_LC_18_5_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_6_LC_18_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78556),
            .lcout(\pid_side.error_d_reg_prevZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94122),
            .ce(N__88053),
            .sr(N__87951));
    defparam \pid_side.error_p_reg_esr_RNINKTC1_7_LC_18_5_6 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNINKTC1_7_LC_18_5_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNINKTC1_7_LC_18_5_6 .LUT_INIT=16'b1000110011101111;
    LogicCell40 \pid_side.error_p_reg_esr_RNINKTC1_7_LC_18_5_6  (
            .in0(N__78555),
            .in1(N__89970),
            .in2(N__72244),
            .in3(N__72490),
            .lcout(\pid_side.error_p_reg_esr_RNINKTC1Z0Z_7 ),
            .ltout(\pid_side.error_p_reg_esr_RNINKTC1Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIKF8V6_7_LC_18_5_7 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIKF8V6_7_LC_18_5_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIKF8V6_7_LC_18_5_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_p_reg_esr_RNIKF8V6_7_LC_18_5_7  (
            .in0(N__72216),
            .in1(N__72351),
            .in2(N__72202),
            .in3(N__72191),
            .lcout(\pid_side.error_p_reg_esr_RNIKF8V6Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_8_LC_18_6_0 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_8_LC_18_6_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_8_LC_18_6_0 .LUT_INIT=16'b1010101000001000;
    LogicCell40 \pid_side.error_i_reg_esr_8_LC_18_6_0  (
            .in0(N__83367),
            .in1(N__73456),
            .in2(N__87430),
            .in3(N__73318),
            .lcout(\pid_side.error_i_regZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94130),
            .ce(N__86777),
            .sr(N__86444));
    defparam \pid_front.error_i_reg_9_sn_rn_1_15_LC_18_6_1 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_9_sn_rn_1_15_LC_18_6_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_9_sn_rn_1_15_LC_18_6_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \pid_front.error_i_reg_9_sn_rn_1_15_LC_18_6_1  (
            .in0(_gnd_net_),
            .in1(N__89377),
            .in2(_gnd_net_),
            .in3(N__87399),
            .lcout(pid_side_error_i_reg_9_sn_rn_1_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNISPTC1_8_LC_18_6_2 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNISPTC1_8_LC_18_6_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNISPTC1_8_LC_18_6_2 .LUT_INIT=16'b1000110011101111;
    LogicCell40 \pid_side.error_p_reg_esr_RNISPTC1_8_LC_18_6_2  (
            .in0(N__79054),
            .in1(N__87823),
            .in2(N__72478),
            .in3(N__72367),
            .lcout(\pid_side.error_p_reg_esr_RNISPTC1Z0Z_8 ),
            .ltout(\pid_side.error_p_reg_esr_RNISPTC1Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIECBV6_8_LC_18_6_3 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIECBV6_8_LC_18_6_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIECBV6_8_LC_18_6_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_side.error_p_reg_esr_RNIECBV6_8_LC_18_6_3  (
            .in0(N__72375),
            .in1(N__72442),
            .in2(N__72424),
            .in3(N__72408),
            .lcout(\pid_side.error_p_reg_esr_RNIECBV6Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNI9GJD3_8_LC_18_6_4 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNI9GJD3_8_LC_18_6_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNI9GJD3_8_LC_18_6_4 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_side.error_p_reg_esr_RNI9GJD3_8_LC_18_6_4  (
            .in0(N__72409),
            .in1(_gnd_net_),
            .in2(N__72385),
            .in3(N__72376),
            .lcout(\pid_side.error_p_reg_esr_RNI9GJD3Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNI1VTC1_0_9_LC_18_6_5 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNI1VTC1_0_9_LC_18_6_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNI1VTC1_0_9_LC_18_6_5 .LUT_INIT=16'b0110001110011100;
    LogicCell40 \pid_side.error_p_reg_esr_RNI1VTC1_0_9_LC_18_6_5  (
            .in0(N__81684),
            .in1(N__89940),
            .in2(N__72835),
            .in3(N__72772),
            .lcout(\pid_side.error_p_reg_esr_RNI1VTC1_0Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI0UEI_8_LC_18_6_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI0UEI_8_LC_18_6_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI0UEI_8_LC_18_6_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI0UEI_8_LC_18_6_6  (
            .in0(_gnd_net_),
            .in1(N__72831),
            .in2(_gnd_net_),
            .in3(N__81683),
            .lcout(\pid_side.N_2577_i ),
            .ltout(\pid_side.N_2577_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNISPTC1_0_8_LC_18_6_7 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNISPTC1_0_8_LC_18_6_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNISPTC1_0_8_LC_18_6_7 .LUT_INIT=16'b0101101010010110;
    LogicCell40 \pid_side.error_p_reg_esr_RNISPTC1_0_8_LC_18_6_7  (
            .in0(N__87822),
            .in1(N__72474),
            .in2(N__72361),
            .in3(N__79053),
            .lcout(\pid_side.error_p_reg_esr_RNISPTC1_0Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNI98EQ_1_LC_18_7_1 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNI98EQ_1_LC_18_7_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNI98EQ_1_LC_18_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_p_reg_esr_RNI98EQ_1_LC_18_7_1  (
            .in0(N__90715),
            .in1(N__82534),
            .in2(_gnd_net_),
            .in3(N__82497),
            .lcout(),
            .ltout(\pid_side.un1_pid_prereg_9_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIM6H42_0_LC_18_7_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIM6H42_0_LC_18_7_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIM6H42_0_LC_18_7_2 .LUT_INIT=16'b0010110100101101;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIM6H42_0_LC_18_7_2  (
            .in0(N__76735),
            .in1(N__79399),
            .in2(N__72340),
            .in3(N__72337),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIM6H42Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIVDLL1_0_21_LC_18_7_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIVDLL1_0_21_LC_18_7_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIVDLL1_0_21_LC_18_7_3 .LUT_INIT=16'b0001111010000111;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIVDLL1_0_21_LC_18_7_3  (
            .in0(N__91383),
            .in1(N__91651),
            .in2(N__72616),
            .in3(N__72924),
            .lcout(\pid_side.un1_pid_prereg_0_25 ),
            .ltout(\pid_side.un1_pid_prereg_0_25_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNITP9B3_21_LC_18_7_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNITP9B3_21_LC_18_7_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNITP9B3_21_LC_18_7_4 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNITP9B3_21_LC_18_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__72733),
            .in3(N__72726),
            .lcout(\pid_side.error_d_reg_prev_esr_RNITP9B3Z0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIHEJ01_0_LC_18_7_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIHEJ01_0_LC_18_7_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIHEJ01_0_LC_18_7_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIHEJ01_0_LC_18_7_5  (
            .in0(N__72703),
            .in1(N__76734),
            .in2(_gnd_net_),
            .in3(N__79398),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIHEJ01Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIQ5IL1_0_21_LC_18_7_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIQ5IL1_0_21_LC_18_7_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIQ5IL1_0_21_LC_18_7_6 .LUT_INIT=16'b0001100011100111;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIQ5IL1_0_21_LC_18_7_6  (
            .in0(N__91649),
            .in1(N__91381),
            .in2(N__72947),
            .in3(N__72664),
            .lcout(\pid_side.un1_pid_prereg_0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIVDLL1_21_LC_18_7_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIVDLL1_21_LC_18_7_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIVDLL1_21_LC_18_7_7 .LUT_INIT=16'b1110000011111000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIVDLL1_21_LC_18_7_7  (
            .in0(N__91382),
            .in1(N__91650),
            .in2(N__72615),
            .in3(N__72923),
            .lcout(\pid_side.un1_pid_prereg_0_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNITU3P4_10_LC_18_8_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNITU3P4_10_LC_18_8_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNITU3P4_10_LC_18_8_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNITU3P4_10_LC_18_8_0  (
            .in0(_gnd_net_),
            .in1(N__72565),
            .in2(_gnd_net_),
            .in3(N__72524),
            .lcout(\pid_side.error_d_reg_prev_esr_RNITU3P4Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIUREI_7_LC_18_8_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIUREI_7_LC_18_8_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIUREI_7_LC_18_8_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIUREI_7_LC_18_8_1  (
            .in0(_gnd_net_),
            .in1(N__72468),
            .in2(_gnd_net_),
            .in3(N__79046),
            .lcout(\pid_side.N_2571_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_7_LC_18_8_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_7_LC_18_8_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_7_LC_18_8_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_7_LC_18_8_2  (
            .in0(N__79047),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94147),
            .ce(N__87991),
            .sr(N__87961));
    defparam \pid_side.state_RNI7OA81_0_LC_18_8_3 .C_ON=1'b0;
    defparam \pid_side.state_RNI7OA81_0_LC_18_8_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.state_RNI7OA81_0_LC_18_8_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pid_side.state_RNI7OA81_0_LC_18_8_3  (
            .in0(_gnd_net_),
            .in1(N__72457),
            .in2(_gnd_net_),
            .in3(N__87960),
            .lcout(\pid_side.N_834_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_8_LC_18_8_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_8_LC_18_8_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_8_LC_18_8_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_8_LC_18_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81682),
            .lcout(\pid_side.error_d_reg_prevZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94147),
            .ce(N__87991),
            .sr(N__87961));
    defparam \pid_side.error_d_reg_prev_esr_14_LC_18_8_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_14_LC_18_8_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_14_LC_18_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_14_LC_18_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__91441),
            .lcout(\pid_side.error_d_reg_prevZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94147),
            .ce(N__87991),
            .sr(N__87961));
    defparam \pid_side.error_d_reg_prev_fast_esr_12_LC_18_8_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_fast_esr_12_LC_18_8_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_fast_esr_12_LC_18_8_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_prev_fast_esr_12_LC_18_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__91243),
            .lcout(\pid_side.error_d_reg_prev_fastZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94147),
            .ce(N__87991),
            .sr(N__87961));
    defparam \pid_side.error_d_reg_prev_esr_21_LC_18_8_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_21_LC_18_8_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_21_LC_18_8_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_21_LC_18_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__91378),
            .lcout(\pid_side.error_d_reg_prevZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94147),
            .ce(N__87991),
            .sr(N__87961));
    defparam \pid_side.error_p_reg_esr_RNI1VTC1_9_LC_18_9_0 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNI1VTC1_9_LC_18_9_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNI1VTC1_9_LC_18_9_0 .LUT_INIT=16'b1011000011111011;
    LogicCell40 \pid_side.error_p_reg_esr_RNI1VTC1_9_LC_18_9_0  (
            .in0(N__81688),
            .in1(N__72830),
            .in2(N__89941),
            .in3(N__72771),
            .lcout(\pid_side.error_p_reg_esr_RNI1VTC1Z0Z_9 ),
            .ltout(\pid_side.error_p_reg_esr_RNI1VTC1Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIBMBO6_10_LC_18_9_1 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIBMBO6_10_LC_18_9_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIBMBO6_10_LC_18_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_p_reg_esr_RNIBMBO6_10_LC_18_9_1  (
            .in0(N__72810),
            .in1(N__73122),
            .in2(N__72790),
            .in3(N__73175),
            .lcout(\pid_side.error_p_reg_esr_RNIBMBO6Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIIARG_10_LC_18_9_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIIARG_10_LC_18_9_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIIARG_10_LC_18_9_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIIARG_10_LC_18_9_2  (
            .in0(_gnd_net_),
            .in1(N__73064),
            .in2(_gnd_net_),
            .in3(N__73031),
            .lcout(),
            .ltout(\pid_side.N_2589_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIRE1B1_10_LC_18_9_3 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIRE1B1_10_LC_18_9_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIRE1B1_10_LC_18_9_3 .LUT_INIT=16'b0100101110110100;
    LogicCell40 \pid_side.error_p_reg_esr_RNIRE1B1_10_LC_18_9_3  (
            .in0(N__79224),
            .in1(N__73099),
            .in2(N__72775),
            .in3(N__72990),
            .lcout(\pid_side.error_p_reg_esr_RNIRE1B1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI20FI_9_LC_18_9_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI20FI_9_LC_18_9_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI20FI_9_LC_18_9_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI20FI_9_LC_18_9_4  (
            .in0(_gnd_net_),
            .in1(N__73098),
            .in2(_gnd_net_),
            .in3(N__79223),
            .lcout(\pid_side.N_2583_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIV4S38_10_LC_18_9_5 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIV4S38_10_LC_18_9_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIV4S38_10_LC_18_9_5 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_side.error_p_reg_esr_RNIV4S38_10_LC_18_9_5  (
            .in0(N__73186),
            .in1(N__73176),
            .in2(N__73156),
            .in3(N__73123),
            .lcout(\pid_side.error_p_reg_esr_RNIV4S38Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_9_LC_18_9_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_9_LC_18_9_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_9_LC_18_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_9_LC_18_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79225),
            .lcout(\pid_side.error_d_reg_prevZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94159),
            .ce(N__88020),
            .sr(N__87942));
    defparam \pid_side.error_d_reg_prev_esr_10_LC_18_9_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_10_LC_18_9_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_10_LC_18_9_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_10_LC_18_9_7  (
            .in0(N__73032),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94159),
            .ce(N__88020),
            .sr(N__87942));
    defparam \pid_side.error_d_reg_esr_10_LC_18_10_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_10_LC_18_10_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_10_LC_18_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_10_LC_18_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73051),
            .lcout(\pid_side.error_d_regZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94171),
            .ce(N__92619),
            .sr(N__92980));
    defparam \pid_side.error_p_reg_esr_10_LC_18_10_2 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_10_LC_18_10_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_10_LC_18_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_10_LC_18_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73006),
            .lcout(\pid_side.error_p_regZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94171),
            .ce(N__92619),
            .sr(N__92980));
    defparam \pid_front.m27_2_03_0_a2_0_0_LC_18_11_0 .C_ON=1'b0;
    defparam \pid_front.m27_2_03_0_a2_0_0_LC_18_11_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.m27_2_03_0_a2_0_0_LC_18_11_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \pid_front.m27_2_03_0_a2_0_0_LC_18_11_0  (
            .in0(N__89346),
            .in1(N__89793),
            .in2(_gnd_net_),
            .in3(N__89525),
            .lcout(pid_side_m27_2_03_0_a2_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_6_15_LC_18_11_1 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_6_15_LC_18_11_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_6_15_LC_18_11_1 .LUT_INIT=16'b0010001100100010;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_6_15_LC_18_11_1  (
            .in0(N__89526),
            .in1(N__87780),
            .in2(N__74872),
            .in3(N__89347),
            .lcout(),
            .ltout(\pid_front.m19_2_03_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_2_15_LC_18_11_2 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_2_15_LC_18_11_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_2_15_LC_18_11_2 .LUT_INIT=16'b1101110011111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_2_15_LC_18_11_2  (
            .in0(N__84093),
            .in1(N__74371),
            .in2(N__72973),
            .in3(N__72970),
            .lcout(\pid_front.m19_2_03_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_1_23_LC_18_11_4 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_1_23_LC_18_11_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_1_23_LC_18_11_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_1_23_LC_18_11_4  (
            .in0(N__88984),
            .in1(N__81654),
            .in2(_gnd_net_),
            .in3(N__84934),
            .lcout(),
            .ltout(\pid_side.N_253_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_23_LC_18_11_5 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_23_LC_18_11_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_23_LC_18_11_5 .LUT_INIT=16'b1111111100001100;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_23_LC_18_11_5  (
            .in0(_gnd_net_),
            .in1(N__73275),
            .in2(N__73258),
            .in3(N__76912),
            .lcout(),
            .ltout(\pid_side.m27_2_03_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_23_LC_18_11_6 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_23_LC_18_11_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_23_LC_18_11_6 .LUT_INIT=16'b1000101000000010;
    LogicCell40 \pid_side.error_i_reg_esr_23_LC_18_11_6  (
            .in0(N__87143),
            .in1(N__84323),
            .in2(N__73255),
            .in3(N__73230),
            .lcout(\pid_side.error_i_regZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94186),
            .ce(N__86751),
            .sr(N__86420));
    defparam \pid_side.error_cry_3_c_RNIV5H5C_LC_18_11_7 .C_ON=1'b0;
    defparam \pid_side.error_cry_3_c_RNIV5H5C_LC_18_11_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_3_c_RNIV5H5C_LC_18_11_7 .LUT_INIT=16'b1011111110111011;
    LogicCell40 \pid_side.error_cry_3_c_RNIV5H5C_LC_18_11_7  (
            .in0(N__73240),
            .in1(N__73924),
            .in2(N__84193),
            .in3(N__77028),
            .lcout(\pid_side.m11_2_03_3_i_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_3_14_LC_18_12_0 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_3_14_LC_18_12_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_3_14_LC_18_12_0 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_3_14_LC_18_12_0  (
            .in0(N__85929),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84761),
            .lcout(\pid_side.error_i_reg_esr_RNO_3Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.m66_i_o2_LC_18_12_1 .C_ON=1'b0;
    defparam \pid_side.m66_i_o2_LC_18_12_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.m66_i_o2_LC_18_12_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pid_side.m66_i_o2_LC_18_12_1  (
            .in0(_gnd_net_),
            .in1(N__78502),
            .in2(_gnd_net_),
            .in3(N__80204),
            .lcout(pid_side_N_216),
            .ltout(pid_side_N_216_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_3_17_LC_18_12_2 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_3_17_LC_18_12_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_3_17_LC_18_12_2 .LUT_INIT=16'b1100110100000101;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_3_17_LC_18_12_2  (
            .in0(N__85930),
            .in1(N__76855),
            .in2(N__73207),
            .in3(N__85600),
            .lcout(\pid_side.m21_2_03_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_6_17_LC_18_12_4 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_6_17_LC_18_12_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_6_17_LC_18_12_4 .LUT_INIT=16'b0000001100010111;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_6_17_LC_18_12_4  (
            .in0(N__85928),
            .in1(N__87422),
            .in2(N__89849),
            .in3(N__85133),
            .lcout(),
            .ltout(\pid_side.error_i_reg_esr_RNO_6Z0Z_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_4_17_LC_18_12_5 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_4_17_LC_18_12_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_4_17_LC_18_12_5 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_4_17_LC_18_12_5  (
            .in0(_gnd_net_),
            .in1(N__80340),
            .in2(N__73204),
            .in3(N__73411),
            .lcout(),
            .ltout(\pid_side.m21_2_03_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_17_LC_18_12_6 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_17_LC_18_12_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_17_LC_18_12_6 .LUT_INIT=16'b0000000100000011;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_17_LC_18_12_6  (
            .in0(N__87429),
            .in1(N__73201),
            .in2(N__73195),
            .in3(N__76990),
            .lcout(\pid_side.error_i_reg_esr_RNO_0_0_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_5_17_LC_18_12_7 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_5_17_LC_18_12_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_5_17_LC_18_12_7 .LUT_INIT=16'b0000000000010101;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_5_17_LC_18_12_7  (
            .in0(N__85132),
            .in1(N__89838),
            .in2(N__87436),
            .in3(N__85927),
            .lcout(\pid_side.error_i_reg_esr_RNO_5Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_1_sqmuxa_1_i_o2_LC_18_13_0 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_1_sqmuxa_1_i_o2_LC_18_13_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_1_sqmuxa_1_i_o2_LC_18_13_0 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \pid_front.error_i_acumm_1_sqmuxa_1_i_o2_LC_18_13_0  (
            .in0(N__73405),
            .in1(N__82240),
            .in2(N__83176),
            .in3(N__80187),
            .lcout(pid_side_N_235),
            .ltout(pid_side_N_235_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_3_24_LC_18_13_1 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_3_24_LC_18_13_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_3_24_LC_18_13_1 .LUT_INIT=16'b0000001110101011;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_3_24_LC_18_13_1  (
            .in0(N__76956),
            .in1(N__80410),
            .in2(N__73345),
            .in3(N__81630),
            .lcout(),
            .ltout(\pid_side.m28_2_03_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_2_24_LC_18_13_2 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_2_24_LC_18_13_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_2_24_LC_18_13_2 .LUT_INIT=16'b1111000011111011;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_2_24_LC_18_13_2  (
            .in0(N__81425),
            .in1(N__87388),
            .in2(N__73342),
            .in3(N__85923),
            .lcout(),
            .ltout(\pid_side.m28_2_03_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_24_LC_18_13_3 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_24_LC_18_13_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_24_LC_18_13_3 .LUT_INIT=16'b1000110000000100;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_24_LC_18_13_3  (
            .in0(N__84469),
            .in1(N__87094),
            .in2(N__73339),
            .in3(N__73311),
            .lcout(),
            .ltout(\pid_side.error_i_reg_9_rn_0_24_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_24_LC_18_13_4 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_24_LC_18_13_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_24_LC_18_13_4 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \pid_side.error_i_reg_esr_24_LC_18_13_4  (
            .in0(N__73449),
            .in1(_gnd_net_),
            .in2(N__73336),
            .in3(N__73297),
            .lcout(\pid_side.error_i_regZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94215),
            .ce(N__86759),
            .sr(N__86400));
    defparam \pid_side.error_cry_5_c_RNIR4S86_LC_18_13_6 .C_ON=1'b0;
    defparam \pid_side.error_cry_5_c_RNIR4S86_LC_18_13_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_5_c_RNIR4S86_LC_18_13_6 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \pid_side.error_cry_5_c_RNIR4S86_LC_18_13_6  (
            .in0(N__89837),
            .in1(N__73717),
            .in2(N__87416),
            .in3(N__73702),
            .lcout(\pid_side.m56_0_o2_0 ),
            .ltout(\pid_side.m56_0_o2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_1_24_LC_18_13_7 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_1_24_LC_18_13_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_1_24_LC_18_13_7 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_1_24_LC_18_13_7  (
            .in0(N__84468),
            .in1(N__87374),
            .in2(N__73300),
            .in3(N__87093),
            .lcout(\pid_side.error_i_reg_9_sn_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_2_c_RNI1TK51_LC_18_14_0 .C_ON=1'b0;
    defparam \pid_front.error_cry_2_c_RNI1TK51_LC_18_14_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_2_c_RNI1TK51_LC_18_14_0 .LUT_INIT=16'b0010010101110101;
    LogicCell40 \pid_front.error_cry_2_c_RNI1TK51_LC_18_14_0  (
            .in0(N__82252),
            .in1(N__80011),
            .in2(N__79626),
            .in3(N__74082),
            .lcout(\pid_front.m78_0_m2_1_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_ki_fast_3_rep1_esr_LC_18_14_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_fast_3_rep1_esr_LC_18_14_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_fast_3_rep1_esr_LC_18_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_fast_3_rep1_esr_LC_18_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__92327),
            .lcout(xy_ki_fast_3_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94231),
            .ce(N__83901),
            .sr(N__86390));
    defparam \pid_side.error_cry_2_c_RNI7GEC1_LC_18_14_2 .C_ON=1'b0;
    defparam \pid_side.error_cry_2_c_RNI7GEC1_LC_18_14_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_2_c_RNI7GEC1_LC_18_14_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \pid_side.error_cry_2_c_RNI7GEC1_LC_18_14_2  (
            .in0(N__90235),
            .in1(N__87560),
            .in2(_gnd_net_),
            .in3(N__80867),
            .lcout(\pid_side.N_155 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_2_0_c_RNI7C2S_LC_18_14_3 .C_ON=1'b0;
    defparam \pid_side.error_cry_2_0_c_RNI7C2S_LC_18_14_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_2_0_c_RNI7C2S_LC_18_14_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \pid_side.error_cry_2_0_c_RNI7C2S_LC_18_14_3  (
            .in0(_gnd_net_),
            .in1(N__79612),
            .in2(_gnd_net_),
            .in3(N__83639),
            .lcout(),
            .ltout(\pid_side.error_cry_2_0_c_RNI7C2SZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_2_0_c_RNI7A6P2_LC_18_14_4 .C_ON=1'b0;
    defparam \pid_side.error_cry_2_0_c_RNI7A6P2_LC_18_14_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_2_0_c_RNI7A6P2_LC_18_14_4 .LUT_INIT=16'b0001100101011101;
    LogicCell40 \pid_side.error_cry_2_0_c_RNI7A6P2_LC_18_14_4  (
            .in0(N__82744),
            .in1(N__89562),
            .in2(N__73468),
            .in3(N__83659),
            .lcout(),
            .ltout(\pid_side.error_cry_2_0_c_RNI7A6PZ0Z2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_2_c_RNIKE157_LC_18_14_5 .C_ON=1'b0;
    defparam \pid_side.error_cry_2_c_RNIKE157_LC_18_14_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_2_c_RNIKE157_LC_18_14_5 .LUT_INIT=16'b0101111000001110;
    LogicCell40 \pid_side.error_cry_2_c_RNIKE157_LC_18_14_5  (
            .in0(N__84056),
            .in1(N__73465),
            .in2(N__73459),
            .in3(N__76657),
            .lcout(\pid_side.N_204 ),
            .ltout(\pid_side.N_204_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_0_c_RNIOEIJA_LC_18_14_6 .C_ON=1'b0;
    defparam \pid_side.error_cry_0_c_RNIOEIJA_LC_18_14_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_c_RNIOEIJA_LC_18_14_6 .LUT_INIT=16'b1010000011100100;
    LogicCell40 \pid_side.error_cry_0_c_RNIOEIJA_LC_18_14_6  (
            .in0(N__87403),
            .in1(N__89851),
            .in2(N__73438),
            .in3(N__73435),
            .lcout(\pid_side.m51_0_o2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_1_c_RNI4CLP1_LC_18_15_0 .C_ON=1'b0;
    defparam \pid_side.error_cry_1_c_RNI4CLP1_LC_18_15_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_1_c_RNI4CLP1_LC_18_15_0 .LUT_INIT=16'b0000011110100111;
    LogicCell40 \pid_side.error_cry_1_c_RNI4CLP1_LC_18_15_0  (
            .in0(N__85137),
            .in1(N__82828),
            .in2(N__84186),
            .in3(N__81098),
            .lcout(),
            .ltout(\pid_side.g0_16_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_5_c_RNI1JA04_LC_18_15_1 .C_ON=1'b0;
    defparam \pid_side.error_cry_5_c_RNI1JA04_LC_18_15_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_5_c_RNI1JA04_LC_18_15_1 .LUT_INIT=16'b0100111101001010;
    LogicCell40 \pid_side.error_cry_5_c_RNI1JA04_LC_18_15_1  (
            .in0(N__85127),
            .in1(N__81640),
            .in2(N__73417),
            .in3(N__81525),
            .lcout(\pid_side.N_228 ),
            .ltout(\pid_side.N_228_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_26_LC_18_15_2 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_26_LC_18_15_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_26_LC_18_15_2 .LUT_INIT=16'b0011111101010101;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_26_LC_18_15_2  (
            .in0(N__85909),
            .in1(N__81327),
            .in2(N__73414),
            .in3(N__84560),
            .lcout(),
            .ltout(\pid_side.error_i_reg_9_1_26_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_26_LC_18_15_3 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_26_LC_18_15_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_26_LC_18_15_3 .LUT_INIT=16'b1000110000001100;
    LogicCell40 \pid_side.error_i_reg_esr_26_LC_18_15_3  (
            .in0(N__84562),
            .in1(N__87103),
            .in2(N__73570),
            .in3(N__73542),
            .lcout(\pid_side.error_i_regZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94247),
            .ce(N__86755),
            .sr(N__86382));
    defparam \pid_side.error_cry_1_c_RNI21KO1_LC_18_15_4 .C_ON=1'b0;
    defparam \pid_side.error_cry_1_c_RNI21KO1_LC_18_15_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_1_c_RNI21KO1_LC_18_15_4 .LUT_INIT=16'b0000100001011101;
    LogicCell40 \pid_side.error_cry_1_c_RNI21KO1_LC_18_15_4  (
            .in0(N__90396),
            .in1(N__82827),
            .in2(N__85159),
            .in3(N__81097),
            .lcout(),
            .ltout(\pid_side.m10_2_03_3_i_0_o2_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_5_c_RNIG3A13_LC_18_15_5 .C_ON=1'b0;
    defparam \pid_side.error_cry_5_c_RNIG3A13_LC_18_15_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_5_c_RNIG3A13_LC_18_15_5 .LUT_INIT=16'b1101001111000010;
    LogicCell40 \pid_side.error_cry_5_c_RNIG3A13_LC_18_15_5  (
            .in0(N__78501),
            .in1(N__90397),
            .in2(N__73549),
            .in3(N__81524),
            .lcout(\pid_side.N_207 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_10_LC_18_15_6 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_10_LC_18_15_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_10_LC_18_15_6 .LUT_INIT=16'b1010100010100000;
    LogicCell40 \pid_side.error_i_reg_esr_10_LC_18_15_6  (
            .in0(N__83376),
            .in1(N__81328),
            .in2(N__73546),
            .in3(N__73534),
            .lcout(\pid_side.error_i_regZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94247),
            .ce(N__86755),
            .sr(N__86382));
    defparam \pid_side.error_i_reg_esr_22_LC_18_15_7 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_22_LC_18_15_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_22_LC_18_15_7 .LUT_INIT=16'b1100010010000000;
    LogicCell40 \pid_side.error_i_reg_esr_22_LC_18_15_7  (
            .in0(N__84561),
            .in1(N__87102),
            .in2(N__73510),
            .in3(N__77644),
            .lcout(\pid_side.error_i_regZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94247),
            .ce(N__86755),
            .sr(N__86382));
    defparam \pid_front.error_i_reg_esr_RNO_3_12_LC_18_16_0 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_3_12_LC_18_16_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_3_12_LC_18_16_0 .LUT_INIT=16'b1111001100000101;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_3_12_LC_18_16_0  (
            .in0(N__73796),
            .in1(N__73907),
            .in2(N__90255),
            .in3(N__73477),
            .lcout(\pid_front.N_186_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_5_12_LC_18_16_1 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_5_12_LC_18_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_5_12_LC_18_16_1 .LUT_INIT=16'b0010010101110101;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_5_12_LC_18_16_1  (
            .in0(N__80193),
            .in1(N__74171),
            .in2(N__90253),
            .in3(N__77966),
            .lcout(\pid_front.error_i_reg_esr_RNO_5_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_0_c_RNI1VVU_LC_18_16_2 .C_ON=1'b0;
    defparam \pid_side.error_cry_0_c_RNI1VVU_LC_18_16_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_c_RNI1VVU_LC_18_16_2 .LUT_INIT=16'b0101001100000011;
    LogicCell40 \pid_side.error_cry_0_c_RNI1VVU_LC_18_16_2  (
            .in0(N__90395),
            .in1(N__80192),
            .in2(N__85160),
            .in3(N__81013),
            .lcout(),
            .ltout(\pid_side.m10_2_03_3_i_0_o2_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_4_c_RNI2AAT2_LC_18_16_3 .C_ON=1'b0;
    defparam \pid_side.error_cry_4_c_RNI2AAT2_LC_18_16_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_4_c_RNI2AAT2_LC_18_16_3 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \pid_side.error_cry_4_c_RNI2AAT2_LC_18_16_3  (
            .in0(N__85161),
            .in1(N__80472),
            .in2(N__73471),
            .in3(N__80303),
            .lcout(\pid_side.N_185 ),
            .ltout(\pid_side.N_185_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_4_c_RNI5SCD3_LC_18_16_4 .C_ON=1'b0;
    defparam \pid_side.error_cry_4_c_RNI5SCD3_LC_18_16_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_4_c_RNI5SCD3_LC_18_16_4 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \pid_side.error_cry_4_c_RNI5SCD3_LC_18_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__73927),
            .in3(N__85746),
            .lcout(\pid_side.m11_2_03_3_i_0_o2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_5_19_LC_18_16_5 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_5_19_LC_18_16_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_5_19_LC_18_16_5 .LUT_INIT=16'b0000010011000100;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_5_19_LC_18_16_5  (
            .in0(N__73906),
            .in1(N__85747),
            .in2(N__80214),
            .in3(N__73795),
            .lcout(\pid_front.error_i_reg_esr_RNO_5Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_0_c_RNINCAV_LC_18_16_6 .C_ON=1'b0;
    defparam \pid_front.error_cry_0_0_c_RNINCAV_LC_18_16_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_0_c_RNINCAV_LC_18_16_6 .LUT_INIT=16'b0000111101010101;
    LogicCell40 \pid_front.error_cry_0_0_c_RNINCAV_LC_18_16_6  (
            .in0(N__77967),
            .in1(_gnd_net_),
            .in2(N__74183),
            .in3(N__80194),
            .lcout(\pid_front.N_183 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_5_c_RNIQLS66_LC_18_16_7 .C_ON=1'b0;
    defparam \pid_side.error_cry_5_c_RNIQLS66_LC_18_16_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_5_c_RNIQLS66_LC_18_16_7 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \pid_side.error_cry_5_c_RNIQLS66_LC_18_16_7  (
            .in0(N__89037),
            .in1(N__73713),
            .in2(N__89822),
            .in3(N__73698),
            .lcout(\pid_side.m10_2_03_3_i_0_o2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_4_11_LC_18_17_0 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_4_11_LC_18_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_4_11_LC_18_17_0 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_4_11_LC_18_17_0  (
            .in0(N__78499),
            .in1(N__83318),
            .in2(N__89072),
            .in3(N__80217),
            .lcout(\pid_front.m78_0_a2_sx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_1_c_RNIJE4M2_LC_18_17_1 .C_ON=1'b0;
    defparam \pid_front.error_cry_1_c_RNIJE4M2_LC_18_17_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_1_c_RNIJE4M2_LC_18_17_1 .LUT_INIT=16'b0101010101110111;
    LogicCell40 \pid_front.error_cry_1_c_RNIJE4M2_LC_18_17_1  (
            .in0(N__83491),
            .in1(N__73657),
            .in2(_gnd_net_),
            .in3(N__79783),
            .lcout(),
            .ltout(\pid_front.error_cry_1_c_RNIJE4MZ0Z2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_2_0_c_RNIT6OP8_LC_18_17_2 .C_ON=1'b0;
    defparam \pid_front.error_cry_2_0_c_RNIT6OP8_LC_18_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_2_0_c_RNIT6OP8_LC_18_17_2 .LUT_INIT=16'b1011111100111111;
    LogicCell40 \pid_front.error_cry_2_0_c_RNIT6OP8_LC_18_17_2  (
            .in0(N__73579),
            .in1(N__74194),
            .in2(N__73636),
            .in3(N__73632),
            .lcout(\pid_front.m8_2_03_3_i_0 ),
            .ltout(\pid_front.m8_2_03_3_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_4_LC_18_17_3 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_4_LC_18_17_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_4_LC_18_17_3 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \pid_front.error_i_reg_4_LC_18_17_3  (
            .in0(N__83319),
            .in1(N__82131),
            .in2(N__73600),
            .in3(N__73593),
            .lcout(\pid_front.error_i_regZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94283),
            .ce(),
            .sr(N__86371));
    defparam \pid_front.m58_0_o2_N_2L1_LC_18_17_4 .C_ON=1'b0;
    defparam \pid_front.m58_0_o2_N_2L1_LC_18_17_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.m58_0_o2_N_2L1_LC_18_17_4 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \pid_front.m58_0_o2_N_2L1_LC_18_17_4  (
            .in0(N__89027),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__89563),
            .lcout(\pid_front.m58_0_o2_N_2LZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_1_0_c_RNI590G1_LC_18_17_5 .C_ON=1'b0;
    defparam \pid_front.error_cry_1_0_c_RNI590G1_LC_18_17_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_1_0_c_RNI590G1_LC_18_17_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \pid_front.error_cry_1_0_c_RNI590G1_LC_18_17_5  (
            .in0(N__80218),
            .in1(N__78500),
            .in2(N__85770),
            .in3(N__77857),
            .lcout(),
            .ltout(\pid_front.error_cry_1_0_c_RNI590GZ0Z1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_1_0_c_RNINT963_LC_18_17_6 .C_ON=1'b0;
    defparam \pid_front.error_cry_1_0_c_RNINT963_LC_18_17_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_1_0_c_RNINT963_LC_18_17_6 .LUT_INIT=16'b0000111100001110;
    LogicCell40 \pid_front.error_cry_1_0_c_RNINT963_LC_18_17_6  (
            .in0(N__89233),
            .in1(N__87751),
            .in2(N__74224),
            .in3(N__74207),
            .lcout(\pid_front.error_cry_1_0_c_RNINTZ0Z963 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_c_RNIT3C71_LC_18_18_0 .C_ON=1'b0;
    defparam \pid_front.error_cry_0_c_RNIT3C71_LC_18_18_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_c_RNIT3C71_LC_18_18_0 .LUT_INIT=16'b0001000000011010;
    LogicCell40 \pid_front.error_cry_0_c_RNIT3C71_LC_18_18_0  (
            .in0(N__82253),
            .in1(N__74134),
            .in2(N__83182),
            .in3(N__79998),
            .lcout(),
            .ltout(\pid_front.N_40_0_i_i_o2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_2_c_RNIKGVO2_LC_18_18_1 .C_ON=1'b0;
    defparam \pid_front.error_cry_2_c_RNIKGVO2_LC_18_18_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_2_c_RNIKGVO2_LC_18_18_1 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \pid_front.error_cry_2_c_RNIKGVO2_LC_18_18_1  (
            .in0(N__81244),
            .in1(N__82147),
            .in2(N__74089),
            .in3(N__74077),
            .lcout(\pid_front.error_cry_2_c_RNIKGVOZ0Z2 ),
            .ltout(\pid_front.error_cry_2_c_RNIKGVOZ0Z2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_0_15_LC_18_18_2 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_15_LC_18_18_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_15_LC_18_18_2 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_15_LC_18_18_2  (
            .in0(N__84548),
            .in1(N__84787),
            .in2(N__73993),
            .in3(N__87025),
            .lcout(\pid_front.error_i_reg_9_rn_1_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_4_15_LC_18_18_3 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_4_15_LC_18_18_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_4_15_LC_18_18_3 .LUT_INIT=16'b0010001000000010;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_4_15_LC_18_18_3  (
            .in0(N__87026),
            .in1(N__84549),
            .in2(N__76702),
            .in3(N__73990),
            .lcout(),
            .ltout(\pid_front.error_i_reg_9_sn_rn_0_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_1_15_LC_18_18_4 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_1_15_LC_18_18_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_1_15_LC_18_18_4 .LUT_INIT=16'b0101000011111010;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_1_15_LC_18_18_4  (
            .in0(N__79486),
            .in1(_gnd_net_),
            .in2(N__73972),
            .in3(N__74690),
            .lcout(),
            .ltout(\pid_front.error_i_reg_9_sn_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_15_LC_18_18_5 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_15_LC_18_18_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_15_LC_18_18_5 .LUT_INIT=16'b0000110001011100;
    LogicCell40 \pid_front.error_i_reg_esr_15_LC_18_18_5  (
            .in0(N__73969),
            .in1(N__73960),
            .in2(N__73951),
            .in3(N__73948),
            .lcout(\pid_front.error_i_regZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94298),
            .ce(N__78130),
            .sr(N__86367));
    defparam \pid_front.error_i_reg_esr_RNO_4_19_LC_18_19_0 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_4_19_LC_18_19_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_4_19_LC_18_19_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_4_19_LC_18_19_0  (
            .in0(_gnd_net_),
            .in1(N__87760),
            .in2(_gnd_net_),
            .in3(N__74390),
            .lcout(\pid_front.error_i_reg_esr_RNO_4Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_3_0_c_RNIKJAS1_LC_18_19_1 .C_ON=1'b0;
    defparam \pid_front.error_cry_3_0_c_RNIKJAS1_LC_18_19_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_3_0_c_RNIKJAS1_LC_18_19_1 .LUT_INIT=16'b0000010011000100;
    LogicCell40 \pid_front.error_cry_3_0_c_RNIKJAS1_LC_18_19_1  (
            .in0(N__74266),
            .in1(N__90234),
            .in2(N__90441),
            .in3(N__74814),
            .lcout(\pid_front.N_226 ),
            .ltout(\pid_front.N_226_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_3_17_LC_18_19_2 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_3_17_LC_18_19_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_3_17_LC_18_19_2 .LUT_INIT=16'b1111000100010001;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_3_17_LC_18_19_2  (
            .in0(N__80620),
            .in1(N__84786),
            .in2(N__74545),
            .in3(N__76867),
            .lcout(\pid_front.m21_2_03_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_3_18_LC_18_19_3 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_3_18_LC_18_19_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_3_18_LC_18_19_3 .LUT_INIT=16'b1000100011111000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_3_18_LC_18_19_3  (
            .in0(N__74391),
            .in1(N__85777),
            .in2(N__85573),
            .in3(N__74404),
            .lcout(\pid_front.m22_2_03_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_2_0_c_RNI5ON81_LC_18_19_4 .C_ON=1'b0;
    defparam \pid_front.error_cry_2_0_c_RNI5ON81_LC_18_19_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_2_0_c_RNI5ON81_LC_18_19_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \pid_front.error_cry_2_0_c_RNI5ON81_LC_18_19_4  (
            .in0(N__90431),
            .in1(N__77739),
            .in2(_gnd_net_),
            .in3(N__74496),
            .lcout(\pid_front.N_254 ),
            .ltout(\pid_front.N_254_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_4_16_LC_18_19_5 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_4_16_LC_18_19_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_4_16_LC_18_19_5 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_4_16_LC_18_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__74398),
            .in3(N__81130),
            .lcout(),
            .ltout(\pid_front.error_i_reg_9_N_2L1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_0_16_LC_18_19_6 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_16_LC_18_19_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_16_LC_18_19_6 .LUT_INIT=16'b0000000100000011;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_16_LC_18_19_6  (
            .in0(N__81326),
            .in1(N__74356),
            .in2(N__74395),
            .in3(N__74392),
            .lcout(\pid_front.error_i_reg_esr_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_10_c_RNIUJG21_LC_18_19_7 .C_ON=1'b0;
    defparam \pid_front.error_cry_10_c_RNIUJG21_LC_18_19_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_10_c_RNIUJG21_LC_18_19_7 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \pid_front.error_cry_10_c_RNIUJG21_LC_18_19_7  (
            .in0(N__84785),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80619),
            .lcout(\pid_front.N_594 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_7_c_RNIULJO1_LC_18_20_0 .C_ON=1'b0;
    defparam \pid_front.error_cry_7_c_RNIULJO1_LC_18_20_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_7_c_RNIULJO1_LC_18_20_0 .LUT_INIT=16'b0011001000000010;
    LogicCell40 \pid_front.error_cry_7_c_RNIULJO1_LC_18_20_0  (
            .in0(N__74311),
            .in1(N__90436),
            .in2(N__85180),
            .in3(N__79904),
            .lcout(\pid_front.N_611 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_4_13_LC_18_20_1 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_4_13_LC_18_20_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_4_13_LC_18_20_1 .LUT_INIT=16'b0100000001110000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_4_13_LC_18_20_1  (
            .in0(N__79905),
            .in1(N__90222),
            .in2(N__90442),
            .in3(N__74312),
            .lcout(),
            .ltout(\pid_front.N_569_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_0_13_LC_18_20_2 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_13_LC_18_20_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_13_LC_18_20_2 .LUT_INIT=16'b1010000010101000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_13_LC_18_20_2  (
            .in0(N__76900),
            .in1(N__74968),
            .in2(N__74875),
            .in3(N__74856),
            .lcout(),
            .ltout(\pid_front.N_436_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_13_LC_18_20_3 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_13_LC_18_20_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_13_LC_18_20_3 .LUT_INIT=16'b0100010001001110;
    LogicCell40 \pid_front.error_i_reg_esr_13_LC_18_20_3  (
            .in0(N__74761),
            .in1(N__74755),
            .in2(N__74740),
            .in3(N__74644),
            .lcout(\pid_front.error_i_regZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94330),
            .ce(N__78110),
            .sr(N__86360));
    defparam \pid_front.error_i_reg_esr_RNO_1_13_LC_18_20_4 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_1_13_LC_18_20_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_1_13_LC_18_20_4 .LUT_INIT=16'b0010101000100000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_1_13_LC_18_20_4  (
            .in0(N__89043),
            .in1(N__74722),
            .in2(N__89586),
            .in3(N__74691),
            .lcout(\pid_front.N_437 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.m10_2_03_3_i_0_a2_0_0_LC_18_20_5 .C_ON=1'b0;
    defparam \pid_front.m10_2_03_3_i_0_a2_0_0_LC_18_20_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.m10_2_03_3_i_0_a2_0_0_LC_18_20_5 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \pid_front.m10_2_03_3_i_0_a2_0_0_LC_18_20_5  (
            .in0(N__90437),
            .in1(N__90675),
            .in2(_gnd_net_),
            .in3(N__90221),
            .lcout(\pid_front.m10_2_03_3_i_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNI2405_3_LC_18_21_0 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI2405_3_LC_18_21_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI2405_3_LC_18_21_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNI2405_3_LC_18_21_0  (
            .in0(N__75243),
            .in1(N__75188),
            .in2(N__74568),
            .in3(N__75471),
            .lcout(\pid_front.error_i_acumm_13_0_a2_2_2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNIU2OK_5_LC_18_21_1 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIU2OK_5_LC_18_21_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIU2OK_5_LC_18_21_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNIU2OK_5_LC_18_21_1  (
            .in0(N__75242),
            .in1(N__75020),
            .in2(N__75192),
            .in3(N__75108),
            .lcout(\pid_front.N_603 ),
            .ltout(\pid_front.N_603_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNI3CD01_3_LC_18_21_2 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI3CD01_3_LC_18_21_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI3CD01_3_LC_18_21_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNI3CD01_3_LC_18_21_2  (
            .in0(N__75966),
            .in1(N__74564),
            .in2(N__74608),
            .in3(N__75470),
            .lcout(\pid_front.error_i_acumm_13_0_a2_3_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_3_LC_18_21_3 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_3_LC_18_21_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_3_LC_18_21_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_3_LC_18_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74593),
            .lcout(\pid_front.error_i_acumm16lto3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94345),
            .ce(N__75328),
            .sr(N__86358));
    defparam \pid_front.error_i_acumm_prereg_esr_5_LC_18_21_4 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_5_LC_18_21_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_5_LC_18_21_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_5_LC_18_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75283),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94345),
            .ce(N__75328),
            .sr(N__86358));
    defparam \pid_front.error_i_acumm_prereg_esr_6_LC_18_21_5 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_6_LC_18_21_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_6_LC_18_21_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_6_LC_18_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75224),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94345),
            .ce(N__75328),
            .sr(N__86358));
    defparam \pid_front.error_i_acumm_prereg_esr_10_LC_18_21_6 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_10_LC_18_21_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_10_LC_18_21_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_10_LC_18_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75172),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94345),
            .ce(N__75328),
            .sr(N__86358));
    defparam \pid_front.error_i_acumm_prereg_esr_11_LC_18_21_7 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_11_LC_18_21_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_11_LC_18_21_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_11_LC_18_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75144),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94345),
            .ce(N__75328),
            .sr(N__86358));
    defparam \pid_front.error_i_acumm_RNO_0_10_LC_18_22_0 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_RNO_0_10_LC_18_22_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_RNO_0_10_LC_18_22_0 .LUT_INIT=16'b0000111100001011;
    LogicCell40 \pid_front.error_i_acumm_RNO_0_10_LC_18_22_0  (
            .in0(N__75653),
            .in1(N__75109),
            .in2(N__75956),
            .in3(N__75999),
            .lcout(),
            .ltout(\pid_front.N_355_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_10_LC_18_22_1 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_10_LC_18_22_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_10_LC_18_22_1 .LUT_INIT=16'b0000001100000010;
    LogicCell40 \pid_front.error_i_acumm_10_LC_18_22_1  (
            .in0(N__75110),
            .in1(N__75865),
            .in2(N__75073),
            .in3(N__75791),
            .lcout(\pid_front.error_i_acummZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94360),
            .ce(N__75766),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNI09AI4_12_LC_18_22_2 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI09AI4_12_LC_18_22_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI09AI4_12_LC_18_22_2 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNI09AI4_12_LC_18_22_2  (
            .in0(_gnd_net_),
            .in1(N__75651),
            .in2(_gnd_net_),
            .in3(N__75058),
            .lcout(\pid_front.N_285 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_RNO_0_11_LC_18_22_4 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_RNO_0_11_LC_18_22_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_RNO_0_11_LC_18_22_4 .LUT_INIT=16'b0000111100001011;
    LogicCell40 \pid_front.error_i_acumm_RNO_0_11_LC_18_22_4  (
            .in0(N__75654),
            .in1(N__75024),
            .in2(N__75957),
            .in3(N__76000),
            .lcout(),
            .ltout(\pid_front.N_353_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_11_LC_18_22_5 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_11_LC_18_22_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_11_LC_18_22_5 .LUT_INIT=16'b0000001100000010;
    LogicCell40 \pid_front.error_i_acumm_11_LC_18_22_5  (
            .in0(N__75025),
            .in1(N__75866),
            .in2(N__74983),
            .in3(N__75792),
            .lcout(\pid_front.error_i_acummZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94360),
            .ce(N__75766),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_RNO_0_12_LC_18_22_6 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_RNO_0_12_LC_18_22_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_RNO_0_12_LC_18_22_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pid_front.error_i_acumm_RNO_0_12_LC_18_22_6  (
            .in0(_gnd_net_),
            .in1(N__75652),
            .in2(_gnd_net_),
            .in3(N__75998),
            .lcout(),
            .ltout(\pid_front.N_242_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_12_LC_18_22_7 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_12_LC_18_22_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_12_LC_18_22_7 .LUT_INIT=16'b0001000000110000;
    LogicCell40 \pid_front.error_i_acumm_12_LC_18_22_7  (
            .in0(N__75933),
            .in1(N__75867),
            .in2(N__75796),
            .in3(N__75793),
            .lcout(\pid_front.error_i_acummZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94360),
            .ce(N__75766),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_12_LC_18_23_0 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_12_LC_18_23_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_12_LC_18_23_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_12_LC_18_23_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75700),
            .lcout(\pid_front.un10lto12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94368),
            .ce(N__75326),
            .sr(N__86354));
    defparam \pid_front.error_i_acumm_prereg_esr_1_LC_18_23_1 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_1_LC_18_23_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_1_LC_18_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_1_LC_18_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75615),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94368),
            .ce(N__75326),
            .sr(N__86354));
    defparam \pid_front.error_i_acumm_prereg_esr_2_LC_18_23_2 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_2_LC_18_23_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_2_LC_18_23_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_2_LC_18_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75557),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94368),
            .ce(N__75326),
            .sr(N__86354));
    defparam \pid_front.error_i_acumm_prereg_esr_4_LC_18_23_3 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_4_LC_18_23_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_4_LC_18_23_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_4_LC_18_23_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75511),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94368),
            .ce(N__75326),
            .sr(N__86354));
    defparam \pid_front.error_i_acumm_prereg_esr_7_LC_18_23_4 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_7_LC_18_23_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_7_LC_18_23_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_7_LC_18_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75449),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94368),
            .ce(N__75326),
            .sr(N__86354));
    defparam \pid_front.error_i_acumm_prereg_esr_8_LC_18_23_5 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_8_LC_18_23_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_8_LC_18_23_5 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_8_LC_18_23_5  (
            .in0(_gnd_net_),
            .in1(N__75382),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94368),
            .ce(N__75326),
            .sr(N__86354));
    defparam \pid_front.error_p_reg_esr_RNITCC61_18_LC_18_24_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNITCC61_18_LC_18_24_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNITCC61_18_LC_18_24_2 .LUT_INIT=16'b1000100011101110;
    LogicCell40 \pid_front.error_p_reg_esr_RNITCC61_18_LC_18_24_2  (
            .in0(N__81958),
            .in1(N__76192),
            .in2(_gnd_net_),
            .in3(N__76165),
            .lcout(\pid_front.error_p_reg_esr_RNITCC61Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNI6FM11_6_LC_20_5_6 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNI6FM11_6_LC_20_5_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNI6FM11_6_LC_20_5_6 .LUT_INIT=16'b1100001101101001;
    LogicCell40 \pid_side.error_p_reg_esr_RNI6FM11_6_LC_20_5_6  (
            .in0(N__76273),
            .in1(N__78542),
            .in2(N__90014),
            .in3(N__78613),
            .lcout(\pid_side.error_p_reg_esr_RNI6FM11Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_1_LC_20_6_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_1_LC_20_6_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_1_LC_20_6_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_1_LC_20_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82498),
            .lcout(\pid_side.error_d_reg_prevZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94148),
            .ce(N__88106),
            .sr(N__87953));
    defparam \pid_side.error_p_reg_esr_RNI76TK1_5_LC_20_7_7 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNI76TK1_5_LC_20_7_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNI76TK1_5_LC_20_7_7 .LUT_INIT=16'b1011001011101000;
    LogicCell40 \pid_side.error_p_reg_esr_RNI76TK1_5_LC_20_7_7  (
            .in0(N__76105),
            .in1(N__76285),
            .in2(N__89908),
            .in3(N__78607),
            .lcout(\pid_side.error_p_reg_esr_RNI76TK1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIIHEQ_4_LC_20_8_0 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIIHEQ_4_LC_20_8_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIIHEQ_4_LC_20_8_0 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_side.error_p_reg_esr_RNIIHEQ_4_LC_20_8_0  (
            .in0(N__82545),
            .in1(N__76371),
            .in2(_gnd_net_),
            .in3(N__87881),
            .lcout(\pid_side.error_p_reg_esr_RNIIHEQZ0Z_4 ),
            .ltout(\pid_side.error_p_reg_esr_RNIIHEQZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNI76TK1_0_5_LC_20_8_1 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNI76TK1_0_5_LC_20_8_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNI76TK1_0_5_LC_20_8_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \pid_side.error_p_reg_esr_RNI76TK1_0_5_LC_20_8_1  (
            .in0(N__89901),
            .in1(N__76284),
            .in2(N__76099),
            .in3(N__78606),
            .lcout(\pid_side.error_p_reg_esr_RNI76TK1_0Z0Z_5 ),
            .ltout(\pid_side.error_p_reg_esr_RNI76TK1_0Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIG7MC2_5_LC_20_8_2 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIG7MC2_5_LC_20_8_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIG7MC2_5_LC_20_8_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_side.error_p_reg_esr_RNIG7MC2_5_LC_20_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__76096),
            .in3(N__76052),
            .lcout(\pid_side.error_p_reg_esr_RNIG7MC2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_4_LC_20_8_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_4_LC_20_8_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_4_LC_20_8_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_4_LC_20_8_3  (
            .in0(N__87883),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94172),
            .ce(N__88054),
            .sr(N__87948));
    defparam \pid_side.error_p_reg_esr_RNIG7MC2_0_5_LC_20_8_4 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIG7MC2_0_5_LC_20_8_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIG7MC2_0_5_LC_20_8_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_side.error_p_reg_esr_RNIG7MC2_0_5_LC_20_8_4  (
            .in0(_gnd_net_),
            .in1(N__76071),
            .in2(_gnd_net_),
            .in3(N__76051),
            .lcout(\pid_side.error_p_reg_esr_RNIG7MC2_0Z0Z_5 ),
            .ltout(\pid_side.error_p_reg_esr_RNIG7MC2_0Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIN4BP4_3_LC_20_8_5 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIN4BP4_3_LC_20_8_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIN4BP4_3_LC_20_8_5 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_side.error_p_reg_esr_RNIN4BP4_3_LC_20_8_5  (
            .in0(N__79249),
            .in1(N__76363),
            .in2(N__76390),
            .in3(N__76353),
            .lcout(\pid_side.error_p_reg_esr_RNIN4BP4Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIIHEQ_0_4_LC_20_8_6 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIIHEQ_0_4_LC_20_8_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIIHEQ_0_4_LC_20_8_6 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_p_reg_esr_RNIIHEQ_0_4_LC_20_8_6  (
            .in0(N__82546),
            .in1(N__76372),
            .in2(_gnd_net_),
            .in3(N__87882),
            .lcout(\pid_side.error_p_reg_esr_RNIIHEQ_0Z0Z_4 ),
            .ltout(\pid_side.error_p_reg_esr_RNIIHEQ_0Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNISL2L4_3_LC_20_8_7 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNISL2L4_3_LC_20_8_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNISL2L4_3_LC_20_8_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_side.error_p_reg_esr_RNISL2L4_3_LC_20_8_7  (
            .in0(N__79248),
            .in1(N__78927),
            .in2(N__76357),
            .in3(N__76352),
            .lcout(\pid_side.error_p_reg_esr_RNISL2L4Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIKAJO_19_LC_20_9_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIKAJO_19_LC_20_9_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIKAJO_19_LC_20_9_1 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIKAJO_19_LC_20_9_1  (
            .in0(N__91129),
            .in1(_gnd_net_),
            .in2(N__82423),
            .in3(N__91051),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIKAJOZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIKAJO_0_19_LC_20_9_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIKAJO_0_19_LC_20_9_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIKAJO_0_19_LC_20_9_2 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIKAJO_0_19_LC_20_9_2  (
            .in0(N__91050),
            .in1(N__82419),
            .in2(_gnd_net_),
            .in3(N__91128),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIKAJO_0Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNI6FM11_0_6_LC_20_9_3 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNI6FM11_0_6_LC_20_9_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNI6FM11_0_6_LC_20_9_3 .LUT_INIT=16'b0101101010010110;
    LogicCell40 \pid_side.error_p_reg_esr_RNI6FM11_0_6_LC_20_9_3  (
            .in0(N__78543),
            .in1(N__76283),
            .in2(N__90016),
            .in3(N__78614),
            .lcout(\pid_side.error_p_reg_esr_RNI6FM11_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_esr_RNI2OIO_3_13_LC_20_10_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_RNI2OIO_3_13_LC_20_10_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_esr_RNI2OIO_3_13_LC_20_10_0 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_d_reg_esr_RNI2OIO_3_13_LC_20_10_0  (
            .in0(N__90899),
            .in1(N__79106),
            .in2(_gnd_net_),
            .in3(N__91482),
            .lcout(\pid_side.error_d_reg_esr_RNI2OIO_3Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_fast_esr_RNIC6BT_12_LC_20_10_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_fast_esr_RNIC6BT_12_LC_20_10_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_fast_esr_RNIC6BT_12_LC_20_10_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \pid_side.error_d_reg_fast_esr_RNIC6BT_12_LC_20_10_1  (
            .in0(N__91483),
            .in1(N__90900),
            .in2(N__79120),
            .in3(N__79316),
            .lcout(),
            .ltout(\pid_side.error_d_reg_fast_esr_RNIC6BTZ0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_fast_esr_RNIKR212_12_LC_20_10_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_fast_esr_RNIKR212_12_LC_20_10_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_fast_esr_RNIKR212_12_LC_20_10_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \pid_side.error_d_reg_prev_fast_esr_RNIKR212_12_LC_20_10_2  (
            .in0(_gnd_net_),
            .in1(N__76237),
            .in2(N__76231),
            .in3(N__76228),
            .lcout(),
            .ltout(\pid_side.g0_3_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIF28I3_12_LC_20_10_3 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIF28I3_12_LC_20_10_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIF28I3_12_LC_20_10_3 .LUT_INIT=16'b1110000110000111;
    LogicCell40 \pid_side.error_p_reg_esr_RNIF28I3_12_LC_20_10_3  (
            .in0(N__76570),
            .in1(N__90974),
            .in2(N__76555),
            .in3(N__82381),
            .lcout(),
            .ltout(\pid_side.g1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNI46CB9_12_LC_20_10_4 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNI46CB9_12_LC_20_10_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNI46CB9_12_LC_20_10_4 .LUT_INIT=16'b1101010001000100;
    LogicCell40 \pid_side.error_p_reg_esr_RNI46CB9_12_LC_20_10_4  (
            .in0(N__79129),
            .in1(N__76552),
            .in2(N__76522),
            .in3(N__76519),
            .lcout(\pid_side.error_p_reg_esr_RNI46CB9Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_13_LC_20_10_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_13_LC_20_10_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_13_LC_20_10_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_13_LC_20_10_5  (
            .in0(N__91484),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94199),
            .ce(N__88119),
            .sr(N__87944));
    defparam \pid_side.error_d_reg_esr_RNI2OIO_0_13_LC_20_10_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_RNI2OIO_0_13_LC_20_10_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_esr_RNI2OIO_0_13_LC_20_10_6 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_side.error_d_reg_esr_RNI2OIO_0_13_LC_20_10_6  (
            .in0(N__90898),
            .in1(N__79105),
            .in2(_gnd_net_),
            .in3(N__91481),
            .lcout(),
            .ltout(\pid_side.N_2608_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI7J5H1_14_LC_20_10_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI7J5H1_14_LC_20_10_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI7J5H1_14_LC_20_10_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI7J5H1_14_LC_20_10_7  (
            .in0(N__90851),
            .in1(N__79173),
            .in2(N__76465),
            .in3(N__91436),
            .lcout(\pid_side.g0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI905J4_1_LC_20_11_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI905J4_1_LC_20_11_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI905J4_1_LC_20_11_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI905J4_1_LC_20_11_0  (
            .in0(N__76710),
            .in1(N__82456),
            .in2(N__76453),
            .in3(N__76396),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI905J4Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIIQL11_1_LC_20_11_1 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIIQL11_1_LC_20_11_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIIQL11_1_LC_20_11_1 .LUT_INIT=16'b1111110011010100;
    LogicCell40 \pid_side.error_p_reg_esr_RNIIQL11_1_LC_20_11_1  (
            .in0(N__76725),
            .in1(N__82479),
            .in2(N__90714),
            .in3(N__79385),
            .lcout(),
            .ltout(\pid_side.error_p_reg_esr_RNIIQL11Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIBGIE2_1_LC_20_11_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIBGIE2_1_LC_20_11_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIBGIE2_1_LC_20_11_2 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIBGIE2_1_LC_20_11_2  (
            .in0(_gnd_net_),
            .in1(N__82532),
            .in2(N__76399),
            .in3(N__76741),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIBGIE2Z0Z_1 ),
            .ltout(\pid_side.error_d_reg_prev_esr_RNIBGIE2Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI9BFR3_1_LC_20_11_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI9BFR3_1_LC_20_11_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI9BFR3_1_LC_20_11_3 .LUT_INIT=16'b1111110011010100;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI9BFR3_1_LC_20_11_3  (
            .in0(N__82533),
            .in1(N__76711),
            .in2(N__76744),
            .in3(N__82480),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI9BFR3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIIQL11_0_1_LC_20_11_5 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIIQL11_0_1_LC_20_11_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIIQL11_0_1_LC_20_11_5 .LUT_INIT=16'b1111001101110001;
    LogicCell40 \pid_side.error_p_reg_esr_RNIIQL11_0_1_LC_20_11_5  (
            .in0(N__76724),
            .in1(N__82478),
            .in2(N__90713),
            .in3(N__79384),
            .lcout(\pid_side.error_p_reg_esr_RNIIQL11_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_0_LC_20_11_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_0_LC_20_11_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_0_LC_20_11_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_0_LC_20_11_6  (
            .in0(N__79386),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94217),
            .ce(N__88089),
            .sr(N__87943));
    defparam \pid_side.error_p_reg_esr_RNICBEQ_0_2_LC_20_11_7 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNICBEQ_0_2_LC_20_11_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNICBEQ_0_2_LC_20_11_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_p_reg_esr_RNICBEQ_0_2_LC_20_11_7  (
            .in0(N__79344),
            .in1(N__78904),
            .in2(_gnd_net_),
            .in3(N__79275),
            .lcout(\pid_side.error_p_reg_esr_RNICBEQ_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_5_15_LC_20_12_0 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_5_15_LC_20_12_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_5_15_LC_20_12_0 .LUT_INIT=16'b0100010000000100;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_5_15_LC_20_12_0  (
            .in0(N__84546),
            .in1(N__87114),
            .in2(N__76698),
            .in3(N__76999),
            .lcout(),
            .ltout(\pid_side.error_i_reg_9_sn_rn_0_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_1_15_LC_20_12_1 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_1_15_LC_20_12_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_1_15_LC_20_12_1 .LUT_INIT=16'b0101010111110000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_1_15_LC_20_12_1  (
            .in0(N__80080),
            .in1(_gnd_net_),
            .in2(N__76669),
            .in3(N__76666),
            .lcout(\pid_side.error_i_reg_9_sn_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_3_0_c_RNI58HU3_LC_20_12_2 .C_ON=1'b0;
    defparam \pid_side.error_cry_3_0_c_RNI58HU3_LC_20_12_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_3_0_c_RNI58HU3_LC_20_12_2 .LUT_INIT=16'b0011001100001010;
    LogicCell40 \pid_side.error_cry_3_0_c_RNI58HU3_LC_20_12_2  (
            .in0(N__89246),
            .in1(N__76656),
            .in2(N__85252),
            .in3(N__84082),
            .lcout(\pid_side.N_258 ),
            .ltout(\pid_side.N_258_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_2_15_LC_20_12_3 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_2_15_LC_20_12_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_2_15_LC_20_12_3 .LUT_INIT=16'b0011000001110101;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_2_15_LC_20_12_3  (
            .in0(N__84827),
            .in1(N__87750),
            .in2(N__76618),
            .in3(N__85926),
            .lcout(),
            .ltout(\pid_side.m19_2_03_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_15_LC_20_12_4 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_15_LC_20_12_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_15_LC_20_12_4 .LUT_INIT=16'b0000001110101010;
    LogicCell40 \pid_side.error_i_reg_esr_15_LC_20_12_4  (
            .in0(N__76615),
            .in1(N__77344),
            .in2(N__76597),
            .in3(N__76594),
            .lcout(\pid_side.error_i_regZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94233),
            .ce(N__86775),
            .sr(N__86409));
    defparam \pid_side.error_cry_5_c_RNIJK882_LC_20_12_5 .C_ON=1'b0;
    defparam \pid_side.error_cry_5_c_RNIJK882_LC_20_12_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_5_c_RNIJK882_LC_20_12_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \pid_side.error_cry_5_c_RNIJK882_LC_20_12_5  (
            .in0(N__82757),
            .in1(N__81520),
            .in2(_gnd_net_),
            .in3(N__87558),
            .lcout(\pid_side.N_245 ),
            .ltout(\pid_side.N_245_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_2_17_LC_20_12_6 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_2_17_LC_20_12_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_2_17_LC_20_12_6 .LUT_INIT=16'b1100111000000010;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_2_17_LC_20_12_6  (
            .in0(N__89245),
            .in1(N__84081),
            .in2(N__76993),
            .in3(N__80079),
            .lcout(\pid_side.N_262 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.m27_2_03_0_o3_LC_20_13_0 .C_ON=1'b0;
    defparam \pid_front.m27_2_03_0_o3_LC_20_13_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.m27_2_03_0_o3_LC_20_13_0 .LUT_INIT=16'b0011011111111111;
    LogicCell40 \pid_front.m27_2_03_0_o3_LC_20_13_0  (
            .in0(N__90648),
            .in1(N__90378),
            .in2(N__82763),
            .in3(N__85115),
            .lcout(pid_side_N_306),
            .ltout(pid_side_N_306_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_2_23_LC_20_13_1 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_2_23_LC_20_13_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_2_23_LC_20_13_1 .LUT_INIT=16'b0010001011110010;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_2_23_LC_20_13_1  (
            .in0(N__76963),
            .in1(N__80409),
            .in2(N__76915),
            .in3(N__85924),
            .lcout(\pid_side.m27_2_03_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_4_c_RNI5TC22_LC_20_13_2 .C_ON=1'b0;
    defparam \pid_side.error_cry_4_c_RNI5TC22_LC_20_13_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_4_c_RNI5TC22_LC_20_13_2 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \pid_side.error_cry_4_c_RNI5TC22_LC_20_13_2  (
            .in0(N__80283),
            .in1(N__85114),
            .in2(N__80479),
            .in3(N__90376),
            .lcout(\pid_side.N_629 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_5_14_LC_20_13_3 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_5_14_LC_20_13_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_5_14_LC_20_13_3 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_5_14_LC_20_13_3  (
            .in0(N__90377),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80407),
            .lcout(),
            .ltout(\pid_side.error_i_reg_esr_RNO_5Z0Z_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_4_14_LC_20_13_4 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_4_14_LC_20_13_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_4_14_LC_20_13_4 .LUT_INIT=16'b0100000011001000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_4_14_LC_20_13_4  (
            .in0(N__85117),
            .in1(N__76869),
            .in2(N__76765),
            .in3(N__76753),
            .lcout(\pid_side.error_i_reg_esr_RNO_4Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_4_c_RNIEMUO1_LC_20_13_5 .C_ON=1'b0;
    defparam \pid_side.error_cry_4_c_RNIEMUO1_LC_20_13_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_4_c_RNIEMUO1_LC_20_13_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \pid_side.error_cry_4_c_RNIEMUO1_LC_20_13_5  (
            .in0(N__80188),
            .in1(N__80465),
            .in2(_gnd_net_),
            .in3(N__80282),
            .lcout(\pid_side.N_160 ),
            .ltout(\pid_side.N_160_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_8_c_RNIM6373_LC_20_13_6 .C_ON=1'b0;
    defparam \pid_side.error_cry_8_c_RNIM6373_LC_20_13_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_8_c_RNIM6373_LC_20_13_6 .LUT_INIT=16'b0001110100001100;
    LogicCell40 \pid_side.error_cry_8_c_RNIM6373_LC_20_13_6  (
            .in0(N__80408),
            .in1(N__85116),
            .in2(N__76747),
            .in3(N__90379),
            .lcout(\pid_side.N_224 ),
            .ltout(\pid_side.N_224_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_3_13_LC_20_13_7 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_3_13_LC_20_13_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_3_13_LC_20_13_7 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_3_13_LC_20_13_7  (
            .in0(N__89788),
            .in1(N__87279),
            .in2(N__77113),
            .in3(N__77110),
            .lcout(\pid_side.m17_2_03_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.m5_0_03_4_i_i_a2_2_LC_20_14_0 .C_ON=1'b0;
    defparam \pid_side.m5_0_03_4_i_i_a2_2_LC_20_14_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.m5_0_03_4_i_i_a2_2_LC_20_14_0 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \pid_side.m5_0_03_4_i_i_a2_2_LC_20_14_0  (
            .in0(N__82943),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83150),
            .lcout(pid_side_N_491),
            .ltout(pid_side_N_491_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_5_17_LC_20_14_1 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_5_17_LC_20_14_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_5_17_LC_20_14_1 .LUT_INIT=16'b0100111000001010;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_5_17_LC_20_14_1  (
            .in0(N__90131),
            .in1(N__83146),
            .in2(N__77095),
            .in3(N__82945),
            .lcout(),
            .ltout(\pid_front.m21_2_03_0_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_4_17_LC_20_14_2 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_4_17_LC_20_14_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_4_17_LC_20_14_2 .LUT_INIT=16'b0000000100001101;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_4_17_LC_20_14_2  (
            .in0(N__80698),
            .in1(N__89320),
            .in2(N__77092),
            .in3(N__77088),
            .lcout(\pid_front.m21_2_03_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_1_c_RNILA2U_LC_20_14_3 .C_ON=1'b0;
    defparam \pid_side.error_cry_1_c_RNILA2U_LC_20_14_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_1_c_RNILA2U_LC_20_14_3 .LUT_INIT=16'b0001001110011011;
    LogicCell40 \pid_side.error_cry_1_c_RNILA2U_LC_20_14_3  (
            .in0(N__90130),
            .in1(N__82944),
            .in2(N__80853),
            .in3(N__81067),
            .lcout(),
            .ltout(\pid_side.m78_0_m2_1_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_5_c_RNIBQN53_LC_20_14_4 .C_ON=1'b0;
    defparam \pid_side.error_cry_5_c_RNIBQN53_LC_20_14_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_5_c_RNIBQN53_LC_20_14_4 .LUT_INIT=16'b0101111000001110;
    LogicCell40 \pid_side.error_cry_5_c_RNIBQN53_LC_20_14_4  (
            .in0(N__85054),
            .in1(N__81499),
            .in2(N__77035),
            .in3(N__87533),
            .lcout(\pid_side.N_184 ),
            .ltout(\pid_side.N_184_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_5_c_RNICLQM4_LC_20_14_5 .C_ON=1'b0;
    defparam \pid_side.error_cry_5_c_RNICLQM4_LC_20_14_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_5_c_RNICLQM4_LC_20_14_5 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \pid_side.error_cry_5_c_RNICLQM4_LC_20_14_5  (
            .in0(N__89730),
            .in1(N__87270),
            .in2(N__77032),
            .in3(N__83675),
            .lcout(\pid_side.N_229 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_ki_0_rep1_esr_LC_20_14_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_0_rep1_esr_LC_20_14_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_0_rep1_esr_LC_20_14_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_0_rep1_esr_LC_20_14_6  (
            .in0(N__88321),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(xy_ki_0_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94266),
            .ce(N__83898),
            .sr(N__86391));
    defparam \pid_side.error_i_reg_esr_RNO_0_13_LC_20_14_7 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_13_LC_20_14_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_13_LC_20_14_7 .LUT_INIT=16'b0000100010101000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_13_LC_20_14_7  (
            .in0(N__87278),
            .in1(N__80073),
            .in2(N__84116),
            .in3(N__80051),
            .lcout(\pid_side.N_437 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_0_c_inv_LC_20_15_0 .C_ON=1'b1;
    defparam \pid_side.error_cry_0_c_inv_LC_20_15_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_c_inv_LC_20_15_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_side.error_cry_0_c_inv_LC_20_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__77317),
            .in3(N__77332),
            .lcout(\pid_side.error_axb_0 ),
            .ltout(),
            .carryin(bfn_20_15_0_),
            .carryout(\pid_side.error_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_0_c_RNI43F5_LC_20_15_1 .C_ON=1'b1;
    defparam \pid_side.error_cry_0_c_RNI43F5_LC_20_15_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_c_RNI43F5_LC_20_15_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_side.error_cry_0_c_RNI43F5_LC_20_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__77308),
            .in3(N__77290),
            .lcout(\pid_side.error_1 ),
            .ltout(),
            .carryin(\pid_side.error_cry_0 ),
            .carryout(\pid_side.error_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_1_c_RNI66G5_LC_20_15_2 .C_ON=1'b1;
    defparam \pid_side.error_cry_1_c_RNI66G5_LC_20_15_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_1_c_RNI66G5_LC_20_15_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_side.error_cry_1_c_RNI66G5_LC_20_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__77287),
            .in3(N__77269),
            .lcout(\pid_side.error_2 ),
            .ltout(),
            .carryin(\pid_side.error_cry_1 ),
            .carryout(\pid_side.error_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_2_c_RNI89H5_LC_20_15_3 .C_ON=1'b1;
    defparam \pid_side.error_cry_2_c_RNI89H5_LC_20_15_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_2_c_RNI89H5_LC_20_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_cry_2_c_RNI89H5_LC_20_15_3  (
            .in0(_gnd_net_),
            .in1(N__77266),
            .in2(_gnd_net_),
            .in3(N__77251),
            .lcout(\pid_side.error_3 ),
            .ltout(),
            .carryin(\pid_side.error_cry_2 ),
            .carryout(\pid_side.error_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_3_c_RNI1SDJ_LC_20_15_4 .C_ON=1'b1;
    defparam \pid_side.error_cry_3_c_RNI1SDJ_LC_20_15_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_3_c_RNI1SDJ_LC_20_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_3_c_RNI1SDJ_LC_20_15_4  (
            .in0(_gnd_net_),
            .in1(N__77248),
            .in2(N__83752),
            .in3(N__77164),
            .lcout(\pid_side.error_4 ),
            .ltout(),
            .carryin(\pid_side.error_cry_3 ),
            .carryout(\pid_side.error_cry_0_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_0_0_c_RNIF3ET_LC_20_15_5 .C_ON=1'b1;
    defparam \pid_side.error_cry_0_0_c_RNIF3ET_LC_20_15_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_0_c_RNIF3ET_LC_20_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_0_0_c_RNIF3ET_LC_20_15_5  (
            .in0(_gnd_net_),
            .in1(N__77161),
            .in2(N__85366),
            .in3(N__77146),
            .lcout(\pid_side.error_5 ),
            .ltout(),
            .carryin(\pid_side.error_cry_0_0 ),
            .carryout(\pid_side.error_cry_1_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_1_0_c_RNII9K11_LC_20_15_6 .C_ON=1'b1;
    defparam \pid_side.error_cry_1_0_c_RNII9K11_LC_20_15_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_1_0_c_RNII9K11_LC_20_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_1_0_c_RNII9K11_LC_20_15_6  (
            .in0(_gnd_net_),
            .in1(N__77143),
            .in2(N__85354),
            .in3(N__77128),
            .lcout(\pid_side.error_6 ),
            .ltout(),
            .carryin(\pid_side.error_cry_1_0 ),
            .carryout(\pid_side.error_cry_2_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_2_0_c_RNILFQL_LC_20_15_7 .C_ON=1'b1;
    defparam \pid_side.error_cry_2_0_c_RNILFQL_LC_20_15_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_2_0_c_RNILFQL_LC_20_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_2_0_c_RNILFQL_LC_20_15_7  (
            .in0(_gnd_net_),
            .in1(N__77125),
            .in2(N__85339),
            .in3(N__77116),
            .lcout(\pid_side.error_7 ),
            .ltout(),
            .carryin(\pid_side.error_cry_2_0 ),
            .carryout(\pid_side.error_cry_3_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_3_0_c_RNIOL0Q_LC_20_16_0 .C_ON=1'b1;
    defparam \pid_side.error_cry_3_0_c_RNIOL0Q_LC_20_16_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_3_0_c_RNIOL0Q_LC_20_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_3_0_c_RNIOL0Q_LC_20_16_0  (
            .in0(_gnd_net_),
            .in1(N__77563),
            .in2(N__85327),
            .in3(N__77548),
            .lcout(\pid_side.error_8 ),
            .ltout(),
            .carryin(bfn_20_16_0_),
            .carryout(\pid_side.error_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_4_c_RNIC8FJ_LC_20_16_1 .C_ON=1'b1;
    defparam \pid_side.error_cry_4_c_RNIC8FJ_LC_20_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_4_c_RNIC8FJ_LC_20_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_4_c_RNIC8FJ_LC_20_16_1  (
            .in0(_gnd_net_),
            .in1(N__77545),
            .in2(N__85312),
            .in3(N__77530),
            .lcout(\pid_side.error_9 ),
            .ltout(),
            .carryin(\pid_side.error_cry_4 ),
            .carryout(\pid_side.error_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_5_c_RNIM4IS_LC_20_16_2 .C_ON=1'b1;
    defparam \pid_side.error_cry_5_c_RNIM4IS_LC_20_16_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_5_c_RNIM4IS_LC_20_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_5_c_RNIM4IS_LC_20_16_2  (
            .in0(_gnd_net_),
            .in1(N__77527),
            .in2(N__85294),
            .in3(N__77518),
            .lcout(\pid_side.error_10 ),
            .ltout(),
            .carryin(\pid_side.error_cry_5 ),
            .carryout(\pid_side.error_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_6_c_RNIQBMT_LC_20_16_3 .C_ON=1'b1;
    defparam \pid_side.error_cry_6_c_RNIQBMT_LC_20_16_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_6_c_RNIQBMT_LC_20_16_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_cry_6_c_RNIQBMT_LC_20_16_3  (
            .in0(_gnd_net_),
            .in1(N__77515),
            .in2(_gnd_net_),
            .in3(N__77500),
            .lcout(\pid_side.error_11 ),
            .ltout(),
            .carryin(\pid_side.error_cry_6 ),
            .carryout(\pid_side.error_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_7_c_RNIPRDP1_LC_20_16_4 .C_ON=1'b1;
    defparam \pid_side.error_cry_7_c_RNIPRDP1_LC_20_16_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_7_c_RNIPRDP1_LC_20_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_7_c_RNIPRDP1_LC_20_16_4  (
            .in0(_gnd_net_),
            .in1(N__77497),
            .in2(N__77482),
            .in3(N__77449),
            .lcout(\pid_side.error_12 ),
            .ltout(),
            .carryin(\pid_side.error_cry_7 ),
            .carryout(\pid_side.error_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_8_c_RNIUUKS_LC_20_16_5 .C_ON=1'b1;
    defparam \pid_side.error_cry_8_c_RNIUUKS_LC_20_16_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_8_c_RNIUUKS_LC_20_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_8_c_RNIUUKS_LC_20_16_5  (
            .in0(_gnd_net_),
            .in1(N__77446),
            .in2(N__77437),
            .in3(N__77413),
            .lcout(\pid_side.error_13 ),
            .ltout(),
            .carryin(\pid_side.error_cry_8 ),
            .carryout(\pid_side.error_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_9_c_RNI13MS_LC_20_16_6 .C_ON=1'b1;
    defparam \pid_side.error_cry_9_c_RNI13MS_LC_20_16_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_9_c_RNI13MS_LC_20_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_9_c_RNI13MS_LC_20_16_6  (
            .in0(_gnd_net_),
            .in1(N__77410),
            .in2(N__77386),
            .in3(N__77401),
            .lcout(\pid_side.error_14 ),
            .ltout(),
            .carryin(\pid_side.error_cry_9 ),
            .carryout(\pid_side.error_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_10_c_RNIBCT11_LC_20_16_7 .C_ON=1'b0;
    defparam \pid_side.error_cry_10_c_RNIBCT11_LC_20_16_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_10_c_RNIBCT11_LC_20_16_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_cry_10_c_RNIBCT11_LC_20_16_7  (
            .in0(N__77398),
            .in1(N__77385),
            .in2(_gnd_net_),
            .in3(N__77371),
            .lcout(\pid_side.error_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_3_15_LC_20_17_0 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_3_15_LC_20_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_3_15_LC_20_17_0 .LUT_INIT=16'b0000111000000010;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_3_15_LC_20_17_0  (
            .in0(N__87586),
            .in1(N__87409),
            .in2(N__89747),
            .in3(N__77367),
            .lcout(\pid_side.m19_2_03_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_ki_esr_0_LC_20_17_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_esr_0_LC_20_17_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_esr_0_LC_20_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_esr_0_LC_20_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88322),
            .lcout(xy_ki_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94315),
            .ce(N__83890),
            .sr(N__86372));
    defparam \pid_side.error_i_reg_esr_RNO_3_22_LC_20_17_2 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_3_22_LC_20_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_3_22_LC_20_17_2 .LUT_INIT=16'b0000111000000100;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_3_22_LC_20_17_2  (
            .in0(N__89081),
            .in1(N__81577),
            .in2(N__89746),
            .in3(N__84896),
            .lcout(\pid_side.error_i_reg_esr_RNO_3Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_4_22_LC_20_17_3 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_4_22_LC_20_17_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_4_22_LC_20_17_3 .LUT_INIT=16'b1110111011111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_4_22_LC_20_17_3  (
            .in0(N__84897),
            .in1(N__89692),
            .in2(N__81602),
            .in3(N__89082),
            .lcout(),
            .ltout(\pid_side.error_i_reg_esr_RNO_4Z0Z_22_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_2_22_LC_20_17_4 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_2_22_LC_20_17_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_2_22_LC_20_17_4 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_2_22_LC_20_17_4  (
            .in0(_gnd_net_),
            .in1(N__77632),
            .in2(N__77656),
            .in3(N__77653),
            .lcout(),
            .ltout(\pid_side.N_297_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_22_LC_20_17_5 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_22_LC_20_17_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_22_LC_20_17_5 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_22_LC_20_17_5  (
            .in0(_gnd_net_),
            .in1(N__81444),
            .in2(N__77647),
            .in3(N__85849),
            .lcout(\pid_side.N_301 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_6_c_RNISNFT1_LC_20_17_6 .C_ON=1'b0;
    defparam \pid_side.error_cry_6_c_RNISNFT1_LC_20_17_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_6_c_RNISNFT1_LC_20_17_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \pid_side.error_cry_6_c_RNISNFT1_LC_20_17_6  (
            .in0(N__89080),
            .in1(N__80376),
            .in2(_gnd_net_),
            .in3(N__87529),
            .lcout(\pid_side.N_252 ),
            .ltout(\pid_side.N_252_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_3_21_LC_20_17_7 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_3_21_LC_20_17_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_3_21_LC_20_17_7 .LUT_INIT=16'b0001000100001111;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_3_21_LC_20_17_7  (
            .in0(N__84898),
            .in1(N__87410),
            .in2(N__77626),
            .in3(N__89696),
            .lcout(\pid_side.un4_error_i_reg_31_am_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_0_c_RNIB56C1_LC_20_18_0 .C_ON=1'b0;
    defparam \pid_side.error_cry_0_c_RNIB56C1_LC_20_18_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_c_RNIB56C1_LC_20_18_0 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \pid_side.error_cry_0_c_RNIB56C1_LC_20_18_0  (
            .in0(N__78496),
            .in1(N__80216),
            .in2(_gnd_net_),
            .in3(N__77623),
            .lcout(),
            .ltout(\pid_side.N_537_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_3_c_RNIDJI03_LC_20_18_1 .C_ON=1'b0;
    defparam \pid_side.error_cry_3_c_RNIDJI03_LC_20_18_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_3_c_RNIDJI03_LC_20_18_1 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \pid_side.error_cry_3_c_RNIDJI03_LC_20_18_1  (
            .in0(N__89748),
            .in1(N__83481),
            .in2(N__77587),
            .in3(N__77584),
            .lcout(\pid_side.m9_2_03_3_i_0_o2_0 ),
            .ltout(\pid_side.m9_2_03_3_i_0_o2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_1_21_LC_20_18_2 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_1_21_LC_20_18_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_1_21_LC_20_18_2 .LUT_INIT=16'b1111111111110100;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_1_21_LC_20_18_2  (
            .in0(N__84835),
            .in1(N__79737),
            .in2(N__78517),
            .in3(N__78193),
            .lcout(\pid_side.error_i_reg_esr_RNO_1Z0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_6_12_LC_20_18_3 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_6_12_LC_20_18_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_6_12_LC_20_18_3 .LUT_INIT=16'b0010010101110101;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_6_12_LC_20_18_3  (
            .in0(N__80215),
            .in1(N__80012),
            .in2(N__79659),
            .in3(N__77810),
            .lcout(),
            .ltout(\pid_front.error_i_reg_esr_RNO_6_0_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_4_12_LC_20_18_4 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_4_12_LC_20_18_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_4_12_LC_20_18_4 .LUT_INIT=16'b0101111000001110;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_4_12_LC_20_18_4  (
            .in0(N__78497),
            .in1(N__78417),
            .in2(N__78328),
            .in3(N__78323),
            .lcout(\pid_front.N_228_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_4_21_LC_20_18_5 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_4_21_LC_20_18_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_4_21_LC_20_18_5 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_4_21_LC_20_18_5  (
            .in0(N__81201),
            .in1(N__79576),
            .in2(_gnd_net_),
            .in3(N__79711),
            .lcout(\pid_side.un4_error_i_reg_31_bm_sx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_1_19_LC_20_19_0 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_1_19_LC_20_19_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_1_19_LC_20_19_0 .LUT_INIT=16'b0000101000011010;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_1_19_LC_20_19_0  (
            .in0(N__84540),
            .in1(N__78826),
            .in2(N__87144),
            .in3(N__78187),
            .lcout(),
            .ltout(\pid_front.error_i_reg_esr_RNO_1_0_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_19_LC_20_19_1 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_19_LC_20_19_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_19_LC_20_19_1 .LUT_INIT=16'b0100101000000000;
    LogicCell40 \pid_front.error_i_reg_esr_19_LC_20_19_1  (
            .in0(N__84541),
            .in1(N__78178),
            .in2(N__78166),
            .in3(N__78832),
            .lcout(\pid_front.error_i_regZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94347),
            .ce(N__78147),
            .sr(N__86364));
    defparam \pid_front.error_cry_0_0_c_RNI7FNK1_LC_20_19_2 .C_ON=1'b0;
    defparam \pid_front.error_cry_0_0_c_RNI7FNK1_LC_20_19_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_0_c_RNI7FNK1_LC_20_19_2 .LUT_INIT=16'b0001000010110000;
    LogicCell40 \pid_front.error_cry_0_0_c_RNI7FNK1_LC_20_19_2  (
            .in0(N__82996),
            .in1(N__77981),
            .in2(N__90685),
            .in3(N__79913),
            .lcout(\pid_front.N_27_0_i_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_2_0_c_RNIUGKS1_LC_20_19_3 .C_ON=1'b0;
    defparam \pid_front.error_cry_2_0_c_RNIUGKS1_LC_20_19_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_2_0_c_RNIUGKS1_LC_20_19_3 .LUT_INIT=16'b0000001000000111;
    LogicCell40 \pid_front.error_cry_2_0_c_RNIUGKS1_LC_20_19_3  (
            .in0(N__82997),
            .in1(N__77871),
            .in2(N__90677),
            .in3(N__77748),
            .lcout(),
            .ltout(\pid_front.N_426_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_0_c_RNIU6KI6_LC_20_19_4 .C_ON=1'b0;
    defparam \pid_front.error_cry_0_0_c_RNIU6KI6_LC_20_19_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_0_c_RNIU6KI6_LC_20_19_4 .LUT_INIT=16'b0000000110101011;
    LogicCell40 \pid_front.error_cry_0_0_c_RNIU6KI6_LC_20_19_4  (
            .in0(N__89535),
            .in1(N__78868),
            .in2(N__78862),
            .in3(N__78859),
            .lcout(\pid_front.m7_2_01 ),
            .ltout(\pid_front.m7_2_01_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_2_19_LC_20_19_5 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_2_19_LC_20_19_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_2_19_LC_20_19_5 .LUT_INIT=16'b0101000101110011;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_2_19_LC_20_19_5  (
            .in0(N__89286),
            .in1(N__84539),
            .in2(N__78847),
            .in3(N__78844),
            .lcout(\pid_front.error_i_reg_esr_RNO_2_0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_3_19_LC_20_20_4 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_3_19_LC_20_20_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_3_19_LC_20_20_4 .LUT_INIT=16'b0001010100010001;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_3_19_LC_20_20_4  (
            .in0(N__80691),
            .in1(N__89287),
            .in2(N__89605),
            .in3(N__81243),
            .lcout(\pid_front.error_i_reg_esr_RNO_3Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_esr_8_LC_20_23_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_8_LC_20_23_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_8_LC_20_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_8_LC_20_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78820),
            .lcout(\pid_front.error_d_regZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94386),
            .ce(N__93395),
            .sr(N__93008));
    defparam \pid_front.error_d_reg_esr_3_LC_20_23_5 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_3_LC_20_23_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_3_LC_20_23_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_3_LC_20_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78778),
            .lcout(\pid_front.error_d_regZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94386),
            .ce(N__93395),
            .sr(N__93008));
    defparam \pid_front.error_d_reg_esr_9_LC_20_24_3 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_9_LC_20_24_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_9_LC_20_24_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_9_LC_20_24_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78748),
            .lcout(\pid_front.error_d_regZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94391),
            .ce(N__93366),
            .sr(N__93009));
    defparam \pid_front.error_d_reg_prev_esr_RNIUO6U_12_LC_20_28_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIUO6U_12_LC_20_28_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIUO6U_12_LC_20_28_6 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIUO6U_12_LC_20_28_6  (
            .in0(_gnd_net_),
            .in1(N__78702),
            .in2(_gnd_net_),
            .in3(N__81819),
            .lcout(\pid_front.N_5_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_esr_5_LC_21_7_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_5_LC_21_7_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_5_LC_21_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_5_LC_21_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78634),
            .lcout(\pid_side.error_d_regZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94173),
            .ce(N__92657),
            .sr(N__92981));
    defparam \pid_side.error_d_reg_esr_6_LC_21_7_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_6_LC_21_7_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_6_LC_21_7_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_6_LC_21_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78574),
            .lcout(\pid_side.error_d_regZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94173),
            .ce(N__92657),
            .sr(N__92981));
    defparam \pid_side.error_d_reg_esr_7_LC_21_7_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_7_LC_21_7_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_7_LC_21_7_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_7_LC_21_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79072),
            .lcout(\pid_side.error_d_regZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94173),
            .ce(N__92657),
            .sr(N__92981));
    defparam \pid_side.error_p_reg_esr_3_LC_21_7_7 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_3_LC_21_7_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_3_LC_21_7_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_3_LC_21_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79027),
            .lcout(\pid_side.error_p_regZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94173),
            .ce(N__92657),
            .sr(N__92981));
    defparam \pid_side.error_p_reg_esr_RNIU3T36_2_LC_21_8_0 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIU3T36_2_LC_21_8_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIU3T36_2_LC_21_8_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_p_reg_esr_RNIU3T36_2_LC_21_8_0  (
            .in0(N__78970),
            .in1(N__78960),
            .in2(N__79014),
            .in3(N__78912),
            .lcout(\pid_side.error_p_reg_esr_RNIU3T36Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNICBEQ_2_LC_21_8_1 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNICBEQ_2_LC_21_8_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNICBEQ_2_LC_21_8_1 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_side.error_p_reg_esr_RNICBEQ_2_LC_21_8_1  (
            .in0(N__79345),
            .in1(N__78903),
            .in2(_gnd_net_),
            .in3(N__79284),
            .lcout(\pid_side.error_p_reg_esr_RNICBEQZ0Z_2 ),
            .ltout(\pid_side.error_p_reg_esr_RNICBEQZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNILOD82_2_LC_21_8_2 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNILOD82_2_LC_21_8_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNILOD82_2_LC_21_8_2 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \pid_side.error_p_reg_esr_RNILOD82_2_LC_21_8_2  (
            .in0(_gnd_net_),
            .in1(N__78913),
            .in2(N__78964),
            .in3(N__78961),
            .lcout(\pid_side.error_p_reg_esr_RNILOD82Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIFEEQ_0_3_LC_21_8_3 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIFEEQ_0_3_LC_21_8_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIFEEQ_0_3_LC_21_8_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_p_reg_esr_RNIFEEQ_0_3_LC_21_8_3  (
            .in0(N__78876),
            .in1(N__78885),
            .in2(_gnd_net_),
            .in3(N__79184),
            .lcout(\pid_side.error_p_reg_esr_RNIFEEQ_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_2_LC_21_8_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_2_LC_21_8_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_2_LC_21_8_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_2_LC_21_8_4  (
            .in0(N__79285),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94187),
            .ce(N__88080),
            .sr(N__87952));
    defparam \pid_side.error_d_reg_prev_esr_3_LC_21_8_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_3_LC_21_8_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_3_LC_21_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_3_LC_21_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79186),
            .lcout(\pid_side.error_d_reg_prevZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94187),
            .ce(N__88080),
            .sr(N__87952));
    defparam \pid_side.error_p_reg_esr_RNIFEEQ_3_LC_21_8_6 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIFEEQ_3_LC_21_8_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIFEEQ_3_LC_21_8_6 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \pid_side.error_p_reg_esr_RNIFEEQ_3_LC_21_8_6  (
            .in0(N__79185),
            .in1(_gnd_net_),
            .in2(N__78889),
            .in3(N__78877),
            .lcout(\pid_side.error_p_reg_esr_RNIFEEQZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_esr_9_LC_21_9_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_9_LC_21_9_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_9_LC_21_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_9_LC_21_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79240),
            .lcout(\pid_side.error_d_regZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94200),
            .ce(N__92656),
            .sr(N__92984));
    defparam \pid_side.error_d_reg_esr_3_LC_21_9_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_3_LC_21_9_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_3_LC_21_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_3_LC_21_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79198),
            .lcout(\pid_side.error_d_regZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94200),
            .ce(N__92656),
            .sr(N__92984));
    defparam \pid_side.error_d_reg_prev_esr_11_LC_21_10_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_11_LC_21_10_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_11_LC_21_10_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_11_LC_21_10_0  (
            .in0(N__83725),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94218),
            .ce(N__88120),
            .sr(N__87946));
    defparam \pid_side.error_d_reg_prev_esr_RNIMERG_0_12_LC_21_10_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIMERG_0_12_LC_21_10_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIMERG_0_12_LC_21_10_1 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIMERG_0_12_LC_21_10_1  (
            .in0(_gnd_net_),
            .in1(N__79466),
            .in2(_gnd_net_),
            .in3(N__91238),
            .lcout(\pid_side.N_5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_fast_esr_RNIFGGE_13_LC_21_10_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_fast_esr_RNIFGGE_13_LC_21_10_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_fast_esr_RNIFGGE_13_LC_21_10_2 .LUT_INIT=16'b1000100011101110;
    LogicCell40 \pid_side.error_d_reg_fast_esr_RNIFGGE_13_LC_21_10_2  (
            .in0(N__82317),
            .in1(N__90907),
            .in2(_gnd_net_),
            .in3(N__79118),
            .lcout(),
            .ltout(\pid_side.N_2608_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIKB371_14_LC_21_10_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIKB371_14_LC_21_10_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIKB371_14_LC_21_10_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIKB371_14_LC_21_10_3  (
            .in0(N__91437),
            .in1(N__79174),
            .in2(N__79141),
            .in3(N__90856),
            .lcout(),
            .ltout(\pid_side.g0_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI7PM14_12_LC_21_10_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI7PM14_12_LC_21_10_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI7PM14_12_LC_21_10_4 .LUT_INIT=16'b1011010000101101;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI7PM14_12_LC_21_10_4  (
            .in0(N__79417),
            .in1(N__79138),
            .in2(N__79132),
            .in3(N__79081),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI7PM14Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_esr_RNI2OIO_2_13_LC_21_10_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_RNI2OIO_2_13_LC_21_10_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_esr_RNI2OIO_2_13_LC_21_10_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_side.error_d_reg_esr_RNI2OIO_2_13_LC_21_10_5  (
            .in0(N__79119),
            .in1(_gnd_net_),
            .in2(N__90917),
            .in3(N__91488),
            .lcout(\pid_side.N_4_1_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNISHIO_2_11_LC_21_10_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNISHIO_2_11_LC_21_10_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNISHIO_2_11_LC_21_10_6 .LUT_INIT=16'b0111011100010001;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNISHIO_2_11_LC_21_10_6  (
            .in0(N__83724),
            .in1(N__91025),
            .in2(_gnd_net_),
            .in3(N__82371),
            .lcout(),
            .ltout(\pid_side.g0_1_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIR65H1_12_LC_21_10_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIR65H1_12_LC_21_10_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIR65H1_12_LC_21_10_7 .LUT_INIT=16'b1001000011111001;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIR65H1_12_LC_21_10_7  (
            .in0(N__79467),
            .in1(N__91239),
            .in2(N__79420),
            .in3(N__90972),
            .lcout(\pid_side.g0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_esr_0_LC_21_11_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_0_LC_21_11_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_0_LC_21_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_0_LC_21_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79411),
            .lcout(\pid_side.error_d_regZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94234),
            .ce(N__92655),
            .sr(N__92989));
    defparam \pid_side.error_d_reg_esr_1_LC_21_11_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_1_LC_21_11_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_1_LC_21_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_1_LC_21_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79369),
            .lcout(\pid_side.error_d_regZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94234),
            .ce(N__92655),
            .sr(N__92989));
    defparam \pid_side.error_p_reg_esr_2_LC_21_11_2 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_2_LC_21_11_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_2_LC_21_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_2_LC_21_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79357),
            .lcout(\pid_side.error_p_regZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94234),
            .ce(N__92655),
            .sr(N__92989));
    defparam \pid_side.error_d_reg_fast_esr_12_LC_21_11_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_fast_esr_12_LC_21_11_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_fast_esr_12_LC_21_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_fast_esr_12_LC_21_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__91270),
            .lcout(\pid_side.error_d_reg_fastZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94234),
            .ce(N__92655),
            .sr(N__92989));
    defparam \pid_side.error_d_reg_esr_2_LC_21_11_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_2_LC_21_11_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_2_LC_21_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_2_LC_21_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79297),
            .lcout(\pid_side.error_d_regZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94234),
            .ce(N__92655),
            .sr(N__92989));
    defparam \pid_side.error_cry_0_0_c_RNIFUCR2_LC_21_12_0 .C_ON=1'b0;
    defparam \pid_side.error_cry_0_0_c_RNIFUCR2_LC_21_12_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_0_c_RNIFUCR2_LC_21_12_0 .LUT_INIT=16'b0011000000111010;
    LogicCell40 \pid_side.error_cry_0_0_c_RNIFUCR2_LC_21_12_0  (
            .in0(N__82759),
            .in1(N__79264),
            .in2(N__90681),
            .in3(N__80287),
            .lcout(),
            .ltout(\pid_side.N_45_i_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_1_0_c_RNILHSE4_LC_21_12_1 .C_ON=1'b0;
    defparam \pid_side.error_cry_1_0_c_RNILHSE4_LC_21_12_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_1_0_c_RNILHSE4_LC_21_12_1 .LUT_INIT=16'b1111000011111100;
    LogicCell40 \pid_side.error_cry_1_0_c_RNILHSE4_LC_21_12_1  (
            .in0(_gnd_net_),
            .in1(N__81260),
            .in2(N__79252),
            .in3(N__82851),
            .lcout(\pid_side.N_8 ),
            .ltout(\pid_side.N_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_18_LC_21_12_2 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_18_LC_21_12_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_18_LC_21_12_2 .LUT_INIT=16'b0000000101000101;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_18_LC_21_12_2  (
            .in0(N__89252),
            .in1(N__84083),
            .in2(N__79558),
            .in3(N__79527),
            .lcout(),
            .ltout(\pid_side.error_i_reg_esr_RNO_0Z0Z_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_18_LC_21_12_3 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_18_LC_21_12_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_18_LC_21_12_3 .LUT_INIT=16'b0000000010110001;
    LogicCell40 \pid_side.error_i_reg_esr_18_LC_21_12_3  (
            .in0(N__84547),
            .in1(N__79534),
            .in2(N__79555),
            .in3(N__84199),
            .lcout(\pid_side.error_i_regZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94249),
            .ce(N__86776),
            .sr(N__86421));
    defparam \pid_side.error_i_reg_esr_RNO_2_18_LC_21_12_4 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_2_18_LC_21_12_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_2_18_LC_21_12_4 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_2_18_LC_21_12_4  (
            .in0(N__89820),
            .in1(N__80341),
            .in2(N__87358),
            .in3(N__87469),
            .lcout(\pid_side.m22_2_03_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_2_LC_21_12_5 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_2_LC_21_12_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_2_LC_21_12_5 .LUT_INIT=16'b0100000001001100;
    LogicCell40 \pid_side.error_i_reg_esr_2_LC_21_12_5  (
            .in0(N__79528),
            .in1(N__82087),
            .in2(N__84132),
            .in3(N__79510),
            .lcout(\pid_side.error_i_regZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94249),
            .ce(N__86776),
            .sr(N__86421));
    defparam \pid_front.error_i_reg_esr_RNO_5_15_LC_21_13_0 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_5_15_LC_21_13_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_5_15_LC_21_13_0 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_5_15_LC_21_13_0  (
            .in0(N__89438),
            .in1(N__87113),
            .in2(N__87330),
            .in3(N__84432),
            .lcout(\pid_front.error_i_reg_9_sn_sn_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_ki_esr_1_LC_21_13_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_esr_1_LC_21_13_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_esr_1_LC_21_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_esr_1_LC_21_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85534),
            .lcout(xy_ki_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94267),
            .ce(N__83877),
            .sr(N__86410));
    defparam \pid_side.error_i_reg_esr_RNO_5_20_LC_21_13_2 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_5_20_LC_21_13_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_5_20_LC_21_13_2 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_5_20_LC_21_13_2  (
            .in0(N__87258),
            .in1(N__89436),
            .in2(_gnd_net_),
            .in3(N__85910),
            .lcout(\pid_side.error_i_reg_esr_RNO_5Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_4_20_LC_21_13_3 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_4_20_LC_21_13_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_4_20_LC_21_13_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_4_20_LC_21_13_3  (
            .in0(N__82752),
            .in1(N__84915),
            .in2(_gnd_net_),
            .in3(N__87559),
            .lcout(),
            .ltout(\pid_side.N_314_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_2_20_LC_21_13_4 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_2_20_LC_21_13_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_2_20_LC_21_13_4 .LUT_INIT=16'b0000101000111011;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_2_20_LC_21_13_4  (
            .in0(N__90078),
            .in1(N__89163),
            .in2(N__79471),
            .in3(N__85912),
            .lcout(),
            .ltout(\pid_side.m24_2_03_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_1_20_LC_21_13_5 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_1_20_LC_21_13_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_1_20_LC_21_13_5 .LUT_INIT=16'b1111111111110100;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_1_20_LC_21_13_5  (
            .in0(N__87749),
            .in1(N__80339),
            .in2(N__79759),
            .in3(N__79747),
            .lcout(\pid_side.m24_2_03_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_6_20_LC_21_13_6 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_6_20_LC_21_13_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_6_20_LC_21_13_6 .LUT_INIT=16'b0101000001010011;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_6_20_LC_21_13_6  (
            .in0(N__89789),
            .in1(N__89437),
            .in2(N__87329),
            .in3(N__85911),
            .lcout(),
            .ltout(\pid_side.error_i_reg_esr_RNO_6Z0Z_20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_3_20_LC_21_13_7 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_3_20_LC_21_13_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_3_20_LC_21_13_7 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_3_20_LC_21_13_7  (
            .in0(N__87468),
            .in1(_gnd_net_),
            .in2(N__79756),
            .in3(N__79753),
            .lcout(\pid_side.m24_2_03_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_2_0_c_RNIO1GV1_LC_21_14_1 .C_ON=1'b0;
    defparam \pid_side.error_cry_2_0_c_RNIO1GV1_LC_21_14_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_2_0_c_RNIO1GV1_LC_21_14_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \pid_side.error_cry_2_0_c_RNIO1GV1_LC_21_14_1  (
            .in0(N__82212),
            .in1(N__82803),
            .in2(_gnd_net_),
            .in3(N__83588),
            .lcout(\pid_side.N_162 ),
            .ltout(\pid_side.N_162_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_3_0_c_RNIM4FM3_LC_21_14_2 .C_ON=1'b0;
    defparam \pid_side.error_cry_3_0_c_RNIM4FM3_LC_21_14_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_3_0_c_RNIM4FM3_LC_21_14_2 .LUT_INIT=16'b1110010010100000;
    LogicCell40 \pid_side.error_cry_3_0_c_RNIM4FM3_LC_21_14_2  (
            .in0(N__90662),
            .in1(N__82689),
            .in2(N__79741),
            .in3(N__85225),
            .lcout(\pid_side.N_206 ),
            .ltout(\pid_side.N_206_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_5_LC_21_14_3 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_5_LC_21_14_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_5_LC_21_14_3 .LUT_INIT=16'b1101110001010000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_5_LC_21_14_3  (
            .in0(N__84834),
            .in1(N__81187),
            .in2(N__79714),
            .in3(N__79710),
            .lcout(),
            .ltout(\pid_side.m9_2_03_3_i_0_o2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_5_LC_21_14_4 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_5_LC_21_14_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_5_LC_21_14_4 .LUT_INIT=16'b1010101010101000;
    LogicCell40 \pid_side.error_i_reg_esr_5_LC_21_14_4  (
            .in0(N__83354),
            .in1(N__79696),
            .in2(N__79684),
            .in3(N__79575),
            .lcout(\pid_side.error_i_regZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94285),
            .ce(N__86784),
            .sr(N__86401));
    defparam \pid_side.m17_2_03_4_a2_7_LC_21_14_5 .C_ON=1'b0;
    defparam \pid_side.m17_2_03_4_a2_7_LC_21_14_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.m17_2_03_4_a2_7_LC_21_14_5 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \pid_side.m17_2_03_4_a2_7_LC_21_14_5  (
            .in0(N__80205),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79625),
            .lcout(pid_side_N_496),
            .ltout(pid_side_N_496_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_2_c_RNILO2S_LC_21_14_6 .C_ON=1'b0;
    defparam \pid_side.error_cry_2_c_RNILO2S_LC_21_14_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_2_c_RNILO2S_LC_21_14_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \pid_side.error_cry_2_c_RNILO2S_LC_21_14_6  (
            .in0(N__89816),
            .in1(N__88971),
            .in2(N__79579),
            .in3(N__80832),
            .lcout(\pid_side.N_536 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_3_12_LC_21_15_0 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_3_12_LC_21_15_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_3_12_LC_21_15_0 .LUT_INIT=16'b1111001100000101;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_3_12_LC_21_15_0  (
            .in0(N__80455),
            .in1(N__80370),
            .in2(N__85077),
            .in3(N__80497),
            .lcout(\pid_side.N_186_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_5_12_LC_21_15_1 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_5_12_LC_21_15_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_5_12_LC_21_15_1 .LUT_INIT=16'b0001010110110101;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_5_12_LC_21_15_1  (
            .in0(N__80207),
            .in1(N__80253),
            .in2(N__85065),
            .in3(N__80978),
            .lcout(\pid_side.error_i_reg_esr_RNO_5Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_4_c_RNILSP52_LC_21_15_2 .C_ON=1'b0;
    defparam \pid_side.error_cry_4_c_RNILSP52_LC_21_15_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_4_c_RNILSP52_LC_21_15_2 .LUT_INIT=16'b0100000001001100;
    LogicCell40 \pid_side.error_cry_4_c_RNILSP52_LC_21_15_2  (
            .in0(N__80454),
            .in1(N__85005),
            .in2(N__89521),
            .in3(N__80369),
            .lcout(\pid_side.N_606 ),
            .ltout(\pid_side.N_606_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_4_c_RNI0E0R2_LC_21_15_3 .C_ON=1'b0;
    defparam \pid_side.error_cry_4_c_RNI0E0R2_LC_21_15_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_4_c_RNI0E0R2_LC_21_15_3 .LUT_INIT=16'b0000010101010101;
    LogicCell40 \pid_side.error_cry_4_c_RNI0E0R2_LC_21_15_3  (
            .in0(N__84419),
            .in1(_gnd_net_),
            .in2(N__80317),
            .in3(N__85776),
            .lcout(\pid_side.un4_error_i_reg_29_ns_sn ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_0_c_RNI6HUA1_LC_21_15_4 .C_ON=1'b0;
    defparam \pid_side.error_cry_0_c_RNI6HUA1_LC_21_15_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_c_RNI6HUA1_LC_21_15_4 .LUT_INIT=16'b0101010100001111;
    LogicCell40 \pid_side.error_cry_0_c_RNI6HUA1_LC_21_15_4  (
            .in0(N__80979),
            .in1(_gnd_net_),
            .in2(N__80281),
            .in3(N__80206),
            .lcout(\pid_side.N_183 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_1_0_c_RNIPBNB2_LC_21_15_5 .C_ON=1'b0;
    defparam \pid_side.error_cry_1_0_c_RNIPBNB2_LC_21_15_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_1_0_c_RNIPBNB2_LC_21_15_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \pid_side.error_cry_1_0_c_RNIPBNB2_LC_21_15_5  (
            .in0(N__81575),
            .in1(N__85025),
            .in2(_gnd_net_),
            .in3(N__82820),
            .lcout(\pid_side.N_188 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_9_c_RNI28JN3_LC_21_15_6 .C_ON=1'b0;
    defparam \pid_side.error_cry_9_c_RNI28JN3_LC_21_15_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_9_c_RNI28JN3_LC_21_15_6 .LUT_INIT=16'b0011000000111010;
    LogicCell40 \pid_side.error_cry_9_c_RNI28JN3_LC_21_15_6  (
            .in0(N__82758),
            .in1(N__80733),
            .in2(N__85076),
            .in3(N__81574),
            .lcout(\pid_side.N_231 ),
            .ltout(\pid_side.N_231_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_1_27_LC_21_15_7 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_1_27_LC_21_15_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_1_27_LC_21_15_7 .LUT_INIT=16'b0001000001010100;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_1_27_LC_21_15_7  (
            .in0(N__87348),
            .in1(N__84087),
            .in2(N__80059),
            .in3(N__80052),
            .lcout(\pid_side.N_339 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_1_c_RNIR72C1_0_LC_21_16_0 .C_ON=1'b0;
    defparam \pid_front.error_cry_1_c_RNIR72C1_0_LC_21_16_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_1_c_RNIR72C1_0_LC_21_16_0 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \pid_front.error_cry_1_c_RNIR72C1_0_LC_21_16_0  (
            .in0(N__82211),
            .in1(N__80003),
            .in2(N__83184),
            .in3(N__79912),
            .lcout(\pid_front.N_525 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_ki_fast_esr_0_LC_21_16_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_fast_esr_0_LC_21_16_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_fast_esr_0_LC_21_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_fast_esr_0_LC_21_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88323),
            .lcout(xy_ki_fast_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94316),
            .ce(N__83878),
            .sr(N__86383));
    defparam \pid_side.error_cry_0_c_RNIDR1R_LC_21_16_2 .C_ON=1'b0;
    defparam \pid_side.error_cry_0_c_RNIDR1R_LC_21_16_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_c_RNIDR1R_LC_21_16_2 .LUT_INIT=16'b0000010000100110;
    LogicCell40 \pid_side.error_cry_0_c_RNIDR1R_LC_21_16_2  (
            .in0(N__83169),
            .in1(N__82186),
            .in2(N__81081),
            .in3(N__80977),
            .lcout(\pid_side.N_40_0_i_i_o2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_2_c_RNINTCQ_LC_21_16_3 .C_ON=1'b0;
    defparam \pid_side.error_cry_2_c_RNINTCQ_LC_21_16_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_2_c_RNINTCQ_LC_21_16_3 .LUT_INIT=16'b0000100000011001;
    LogicCell40 \pid_side.error_cry_2_c_RNINTCQ_LC_21_16_3  (
            .in0(N__82187),
            .in1(N__83170),
            .in2(N__80947),
            .in3(N__80816),
            .lcout(\pid_side.N_40_0_i_i_o2_1 ),
            .ltout(\pid_side.N_40_0_i_i_o2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_0_c_RNIBKF82_LC_21_16_4 .C_ON=1'b0;
    defparam \pid_side.error_cry_0_c_RNIBKF82_LC_21_16_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_c_RNIBKF82_LC_21_16_4 .LUT_INIT=16'b0001000100011101;
    LogicCell40 \pid_side.error_cry_0_c_RNIBKF82_LC_21_16_4  (
            .in0(N__90670),
            .in1(N__90434),
            .in2(N__80776),
            .in3(N__80769),
            .lcout(),
            .ltout(\pid_side.m7_2_01_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_3_c_RNIVVTQ6_LC_21_16_5 .C_ON=1'b0;
    defparam \pid_side.error_cry_3_c_RNIVVTQ6_LC_21_16_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_3_c_RNIVVTQ6_LC_21_16_5 .LUT_INIT=16'b1011000110100001;
    LogicCell40 \pid_side.error_cry_3_c_RNIVVTQ6_LC_21_16_5  (
            .in0(N__84100),
            .in1(N__80755),
            .in2(N__80740),
            .in3(N__80737),
            .lcout(\pid_side.m7_2_01 ),
            .ltout(\pid_side.m7_2_01_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_3_c_RNIET557_LC_21_16_6 .C_ON=1'b0;
    defparam \pid_side.error_cry_3_c_RNIET557_LC_21_16_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_3_c_RNIET557_LC_21_16_6 .LUT_INIT=16'b0011000000000000;
    LogicCell40 \pid_side.error_cry_3_c_RNIET557_LC_21_16_6  (
            .in0(_gnd_net_),
            .in1(N__89232),
            .in2(N__80707),
            .in3(N__84500),
            .lcout(\pid_side.un4_error_i_reg_29_ns_rn_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_2_21_LC_21_17_0 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_2_21_LC_21_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_2_21_LC_21_17_0 .LUT_INIT=16'b0000000001011101;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_2_21_LC_21_17_0  (
            .in0(N__85068),
            .in1(N__87667),
            .in2(N__89531),
            .in3(N__80690),
            .lcout(\pid_front.error_i_reg_9_N_5L8_0_sx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.m17_2_03_4_o3_LC_21_17_1 .C_ON=1'b0;
    defparam \pid_side.m17_2_03_4_o3_LC_21_17_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.m17_2_03_4_o3_LC_21_17_1 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \pid_side.m17_2_03_4_o3_LC_21_17_1  (
            .in0(_gnd_net_),
            .in1(N__83174),
            .in2(_gnd_net_),
            .in3(N__82998),
            .lcout(pid_side_N_164),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_5_c_RNI2TTE2_LC_21_17_2 .C_ON=1'b0;
    defparam \pid_side.error_cry_5_c_RNI2TTE2_LC_21_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_5_c_RNI2TTE2_LC_21_17_2 .LUT_INIT=16'b0000001010100010;
    LogicCell40 \pid_side.error_cry_5_c_RNI2TTE2_LC_21_17_2  (
            .in0(N__85066),
            .in1(N__81576),
            .in2(N__89530),
            .in3(N__81487),
            .lcout(\pid_side.N_225 ),
            .ltout(\pid_side.N_225_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_2_21_LC_21_17_3 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_2_21_LC_21_17_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_2_21_LC_21_17_3 .LUT_INIT=16'b0001000111110000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_2_21_LC_21_17_3  (
            .in0(N__85842),
            .in1(N__89494),
            .in2(N__81448),
            .in3(N__87675),
            .lcout(),
            .ltout(\pid_side.m25_2_03_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_21_LC_21_17_4 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_21_LC_21_17_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_21_LC_21_17_4 .LUT_INIT=16'b0000001000000011;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_21_LC_21_17_4  (
            .in0(N__81445),
            .in1(N__87593),
            .in2(N__81373),
            .in3(N__81370),
            .lcout(),
            .ltout(\pid_side.error_i_reg_esr_RNO_0_0_21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_21_LC_21_17_5 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_21_LC_21_17_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_21_LC_21_17_5 .LUT_INIT=16'b1100100001000000;
    LogicCell40 \pid_side.error_i_reg_esr_21_LC_21_17_5  (
            .in0(N__84504),
            .in1(N__87088),
            .in2(N__81364),
            .in3(N__81361),
            .lcout(\pid_side.error_i_regZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94332),
            .ce(N__86785),
            .sr(N__86376));
    defparam \pid_side.error_cry_10_c_RNIHBAF1_LC_21_17_6 .C_ON=1'b0;
    defparam \pid_side.error_cry_10_c_RNIHBAF1_LC_21_17_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_10_c_RNIHBAF1_LC_21_17_6 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \pid_side.error_cry_10_c_RNIHBAF1_LC_21_17_6  (
            .in0(N__85067),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85841),
            .lcout(\pid_side.N_589 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_2_0_c_RNIKHPR1_LC_21_18_1 .C_ON=1'b0;
    defparam \pid_side.error_cry_2_0_c_RNIKHPR1_LC_21_18_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_2_0_c_RNIKHPR1_LC_21_18_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \pid_side.error_cry_2_0_c_RNIKHPR1_LC_21_18_1  (
            .in0(N__89502),
            .in1(N__83628),
            .in2(_gnd_net_),
            .in3(N__87540),
            .lcout(\pid_side.N_254 ),
            .ltout(\pid_side.N_254_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_5_16_LC_21_18_2 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_5_16_LC_21_18_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_5_16_LC_21_18_2 .LUT_INIT=16'b1010111000001100;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_5_16_LC_21_18_2  (
            .in0(N__85599),
            .in1(N__81126),
            .in2(N__81337),
            .in3(N__81292),
            .lcout(\pid_side.m20_2_03_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.m22_2_03_0_a2_0_0_LC_21_18_3 .C_ON=1'b0;
    defparam \pid_front.m22_2_03_0_a2_0_0_LC_21_18_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.m22_2_03_0_a2_0_0_LC_21_18_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \pid_front.m22_2_03_0_a2_0_0_LC_21_18_3  (
            .in0(N__82999),
            .in1(N__90181),
            .in2(_gnd_net_),
            .in3(N__90667),
            .lcout(pid_side_m22_2_03_0_a2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.m20_2_03_0_a2_0_0_LC_21_18_4 .C_ON=1'b0;
    defparam \pid_front.m20_2_03_0_a2_0_0_LC_21_18_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.m20_2_03_0_a2_0_0_LC_21_18_4 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \pid_front.m20_2_03_0_a2_0_0_LC_21_18_4  (
            .in0(N__90668),
            .in1(_gnd_net_),
            .in2(N__90220),
            .in3(N__83000),
            .lcout(pid_side_m20_2_03_0_a2_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.m5_0_a3_LC_21_18_5 .C_ON=1'b0;
    defparam \pid_front.m5_0_a3_LC_21_18_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.m5_0_a3_LC_21_18_5 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \pid_front.m5_0_a3_LC_21_18_5  (
            .in0(N__83001),
            .in1(_gnd_net_),
            .in2(N__84678),
            .in3(N__90669),
            .lcout(\pid_front.m0_0_03 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.N_40_0_i_i_a2_2_LC_21_18_6 .C_ON=1'b0;
    defparam \pid_front.N_40_0_i_i_a2_2_LC_21_18_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.N_40_0_i_i_a2_2_LC_21_18_6 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \pid_front.N_40_0_i_i_a2_2_LC_21_18_6  (
            .in0(N__83175),
            .in1(N__84671),
            .in2(_gnd_net_),
            .in3(N__82216),
            .lcout(\pid_front.N_574 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_3_LC_21_19_2 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_3_LC_21_19_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_3_LC_21_19_2 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \pid_front.error_i_reg_3_LC_21_19_2  (
            .in0(N__82138),
            .in1(N__82077),
            .in2(N__81990),
            .in3(N__81997),
            .lcout(\pid_front.error_i_regZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94362),
            .ce(),
            .sr(N__86368));
    defparam \pid_front.error_d_reg_esr_18_LC_21_23_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_18_LC_21_23_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_18_LC_21_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_18_LC_21_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81970),
            .lcout(\pid_front.error_d_regZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94392),
            .ce(N__93399),
            .sr(N__93010));
    defparam \pid_front.error_d_reg_esr_2_LC_21_23_5 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_2_LC_21_23_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_2_LC_21_23_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_2_LC_21_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81934),
            .lcout(\pid_front.error_d_regZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94392),
            .ce(N__93399),
            .sr(N__93010));
    defparam \pid_front.error_d_reg_esr_10_LC_21_24_0 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_10_LC_21_24_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_10_LC_21_24_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_10_LC_21_24_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81907),
            .lcout(\pid_front.error_d_regZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94396),
            .ce(N__93367),
            .sr(N__93011));
    defparam \pid_front.error_d_reg_esr_12_LC_21_25_0 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_12_LC_21_25_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_12_LC_21_25_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_12_LC_21_25_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81852),
            .lcout(\pid_front.error_d_regZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94401),
            .ce(N__93369),
            .sr(N__93012));
    defparam \pid_front.error_d_reg_esr_6_LC_21_26_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_6_LC_21_26_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_6_LC_21_26_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_6_LC_21_26_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81766),
            .lcout(\pid_front.error_d_regZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94406),
            .ce(N__93368),
            .sr(N__93014));
    defparam \pid_side.error_d_reg_esr_8_LC_22_8_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_8_LC_22_8_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_8_LC_22_8_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_8_LC_22_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81703),
            .lcout(\pid_side.error_d_regZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94201),
            .ce(N__92651),
            .sr(N__92985));
    defparam \pid_side.error_p_reg_esr_4_LC_22_8_6 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_4_LC_22_8_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_4_LC_22_8_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_4_LC_22_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82558),
            .lcout(\pid_side.error_p_regZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94201),
            .ce(N__92651),
            .sr(N__92985));
    defparam \pid_side.error_d_reg_prev_esr_RNIIFEI_1_LC_22_9_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIIFEI_1_LC_22_9_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIIFEI_1_LC_22_9_3 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIIFEI_1_LC_22_9_3  (
            .in0(_gnd_net_),
            .in1(N__82531),
            .in2(_gnd_net_),
            .in3(N__82490),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIIFEIZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIH7JO_18_LC_22_10_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIH7JO_18_LC_22_10_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIH7JO_18_LC_22_10_0 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIH7JO_18_LC_22_10_0  (
            .in0(N__90748),
            .in1(N__87868),
            .in2(_gnd_net_),
            .in3(N__92754),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIH7JOZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_19_LC_22_10_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_19_LC_22_10_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_19_LC_22_10_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_19_LC_22_10_3  (
            .in0(N__91127),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94235),
            .ce(N__88079),
            .sr(N__87949));
    defparam \pid_side.error_d_reg_prev_esr_RNISHIO_0_11_LC_22_10_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNISHIO_0_11_LC_22_10_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNISHIO_0_11_LC_22_10_5 .LUT_INIT=16'b1000100010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNISHIO_0_11_LC_22_10_5  (
            .in0(N__83721),
            .in1(N__91020),
            .in2(_gnd_net_),
            .in3(N__82368),
            .lcout(\pid_side.un1_pid_prereg_135_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNISHIO_11_LC_22_10_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNISHIO_11_LC_22_10_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNISHIO_11_LC_22_10_6 .LUT_INIT=16'b1111010101010000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNISHIO_11_LC_22_10_6  (
            .in0(N__82370),
            .in1(_gnd_net_),
            .in2(N__91027),
            .in3(N__83723),
            .lcout(\pid_side.g0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNISHIO_1_11_LC_22_10_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNISHIO_1_11_LC_22_10_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNISHIO_1_11_LC_22_10_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNISHIO_1_11_LC_22_10_7  (
            .in0(N__83722),
            .in1(N__91021),
            .in2(_gnd_net_),
            .in3(N__82369),
            .lcout(\pid_side.error_d_reg_prev_esr_RNISHIO_1Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_fast_esr_13_LC_22_11_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_fast_esr_13_LC_22_11_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_fast_esr_13_LC_22_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_fast_esr_13_LC_22_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__91522),
            .lcout(\pid_side.error_d_reg_fastZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94250),
            .ce(N__92678),
            .sr(N__92992));
    defparam \pid_side.error_d_reg_esr_11_LC_22_11_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_11_LC_22_11_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_11_LC_22_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_11_LC_22_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83740),
            .lcout(\pid_side.error_d_regZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94250),
            .ce(N__92678),
            .sr(N__92992));
    defparam \pid_side.error_i_reg_esr_20_LC_22_12_0 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_20_LC_22_12_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_20_LC_22_12_0 .LUT_INIT=16'b1011000000010000;
    LogicCell40 \pid_side.error_i_reg_esr_20_LC_22_12_0  (
            .in0(N__84538),
            .in1(N__83704),
            .in2(N__87145),
            .in3(N__83557),
            .lcout(\pid_side.error_i_regZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94268),
            .ce(N__86761),
            .sr(N__86430));
    defparam \pid_side.error_cry_2_0_c_RNI4KAG3_LC_22_12_1 .C_ON=1'b0;
    defparam \pid_side.error_cry_2_0_c_RNI4KAG3_LC_22_12_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_2_0_c_RNI4KAG3_LC_22_12_1 .LUT_INIT=16'b0000111000000100;
    LogicCell40 \pid_side.error_cry_2_0_c_RNI4KAG3_LC_22_12_1  (
            .in0(N__82765),
            .in1(N__83680),
            .in2(N__84850),
            .in3(N__83635),
            .lcout(\pid_side.N_551 ),
            .ltout(\pid_side.N_551_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_20_LC_22_12_2 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_20_LC_22_12_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_20_LC_22_12_2 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_20_LC_22_12_2  (
            .in0(N__82774),
            .in1(N__83492),
            .in2(N__83560),
            .in3(N__83550),
            .lcout(\pid_side.m8_2_03_3_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_4_LC_22_12_3 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_4_LC_22_12_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_4_LC_22_12_3 .LUT_INIT=16'b1111111110100000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_4_LC_22_12_3  (
            .in0(N__83551),
            .in1(_gnd_net_),
            .in2(N__83510),
            .in3(N__82773),
            .lcout(),
            .ltout(\pid_side.error_i_reg_esr_RNO_0Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_4_LC_22_12_4 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_4_LC_22_12_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_4_LC_22_12_4 .LUT_INIT=16'b1111110000000000;
    LogicCell40 \pid_side.error_i_reg_esr_4_LC_22_12_4  (
            .in0(_gnd_net_),
            .in1(N__83389),
            .in2(N__83383),
            .in3(N__83366),
            .lcout(\pid_side.error_i_regZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94268),
            .ce(N__86761),
            .sr(N__86430));
    defparam \pid_side.error_cry_0_c_RNI0Q6A2_LC_22_12_5 .C_ON=1'b0;
    defparam \pid_side.error_cry_0_c_RNI0Q6A2_LC_22_12_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_c_RNI0Q6A2_LC_22_12_5 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \pid_side.error_cry_0_c_RNI0Q6A2_LC_22_12_5  (
            .in0(N__83177),
            .in1(N__83012),
            .in2(N__85156),
            .in3(N__82878),
            .lcout(),
            .ltout(\pid_side.N_538_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_1_0_c_RNISB0C4_LC_22_12_6 .C_ON=1'b0;
    defparam \pid_side.error_cry_1_0_c_RNISB0C4_LC_22_12_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_1_0_c_RNISB0C4_LC_22_12_6 .LUT_INIT=16'b1111001011110000;
    LogicCell40 \pid_side.error_cry_1_0_c_RNISB0C4_LC_22_12_6  (
            .in0(N__85733),
            .in1(N__84826),
            .in2(N__82864),
            .in3(N__82852),
            .lcout(\pid_side.m58_0_o2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.m58_0_a2_1_sx_LC_22_13_0 .C_ON=1'b0;
    defparam \pid_side.m58_0_a2_1_sx_LC_22_13_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.m58_0_a2_1_sx_LC_22_13_0 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \pid_side.m58_0_a2_1_sx_LC_22_13_0  (
            .in0(N__87271),
            .in1(N__85034),
            .in2(N__84027),
            .in3(N__82751),
            .lcout(\pid_side.m58_0_a2_1_sxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_0_12_LC_22_13_5 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_12_LC_22_13_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_12_LC_22_13_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_12_LC_22_13_5  (
            .in0(N__89787),
            .in1(N__84831),
            .in2(N__84682),
            .in3(N__87272),
            .lcout(\pid_front.m0_2_03 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_1_18_LC_22_13_6 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_1_18_LC_22_13_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_1_18_LC_22_13_6 .LUT_INIT=16'b0101111101001111;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_1_18_LC_22_13_6  (
            .in0(N__84537),
            .in1(N__87600),
            .in2(N__87142),
            .in3(N__85543),
            .lcout(\pid_side.error_i_reg_9_sx_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_ki_1_rep2_esr_LC_22_14_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_1_rep2_esr_LC_22_14_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_1_rep2_esr_LC_22_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_1_rep2_esr_LC_22_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85530),
            .lcout(xy_ki_1_rep2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94300),
            .ce(N__83899),
            .sr(N__86411));
    defparam \Commands_frame_decoder.source_xy_ki_2_rep2_esr_LC_22_14_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_2_rep2_esr_LC_22_14_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_2_rep2_esr_LC_22_14_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_2_rep2_esr_LC_22_14_1  (
            .in0(N__92517),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(xy_ki_2_rep2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94300),
            .ce(N__83899),
            .sr(N__86411));
    defparam \Commands_frame_decoder.source_xy_ki_esr_2_LC_22_14_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_esr_2_LC_22_14_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_esr_2_LC_22_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_esr_2_LC_22_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__92516),
            .lcout(xy_ki_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94300),
            .ce(N__83899),
            .sr(N__86411));
    defparam \Commands_frame_decoder.source_xy_ki_3_rep1_esr_LC_22_14_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_3_rep1_esr_LC_22_14_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_3_rep1_esr_LC_22_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_3_rep1_esr_LC_22_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__92320),
            .lcout(xy_ki_3_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94300),
            .ce(N__83899),
            .sr(N__86411));
    defparam \Commands_frame_decoder.source_xy_ki_3_rep2_esr_LC_22_14_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_3_rep2_esr_LC_22_14_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_3_rep2_esr_LC_22_14_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_3_rep2_esr_LC_22_14_4  (
            .in0(N__92319),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(xy_ki_3_rep2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94300),
            .ce(N__83899),
            .sr(N__86411));
    defparam \Commands_frame_decoder.source_xy_ki_esr_3_LC_22_14_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_esr_3_LC_22_14_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_esr_3_LC_22_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_esr_3_LC_22_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__92321),
            .lcout(xy_ki_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94300),
            .ce(N__83899),
            .sr(N__86411));
    defparam \Commands_frame_decoder.source_CH2data_esr_0_LC_22_15_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_0_LC_22_15_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_0_LC_22_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_0_LC_22_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88324),
            .lcout(side_command_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94317),
            .ce(N__85264),
            .sr(N__86402));
    defparam \Commands_frame_decoder.source_CH2data_esr_1_LC_22_15_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_1_LC_22_15_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_1_LC_22_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_1_LC_22_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85529),
            .lcout(side_command_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94317),
            .ce(N__85264),
            .sr(N__86402));
    defparam \Commands_frame_decoder.source_CH2data_esr_2_LC_22_15_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_2_LC_22_15_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_2_LC_22_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_2_LC_22_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__92518),
            .lcout(side_command_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94317),
            .ce(N__85264),
            .sr(N__86402));
    defparam \Commands_frame_decoder.source_CH2data_esr_3_LC_22_15_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_3_LC_22_15_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_3_LC_22_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_3_LC_22_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__92322),
            .lcout(side_command_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94317),
            .ce(N__85264),
            .sr(N__86402));
    defparam \Commands_frame_decoder.source_CH2data_esr_4_LC_22_15_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_4_LC_22_15_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_4_LC_22_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_4_LC_22_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88854),
            .lcout(side_command_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94317),
            .ce(N__85264),
            .sr(N__86402));
    defparam \Commands_frame_decoder.source_CH2data_esr_5_LC_22_15_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_5_LC_22_15_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_5_LC_22_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_5_LC_22_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88700),
            .lcout(side_command_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94317),
            .ce(N__85264),
            .sr(N__86402));
    defparam \Commands_frame_decoder.source_CH2data_esr_6_LC_22_15_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_6_LC_22_15_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_6_LC_22_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_6_LC_22_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88507),
            .lcout(side_command_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94317),
            .ce(N__85264),
            .sr(N__86402));
    defparam \Commands_frame_decoder.source_CH2data_ess_7_LC_22_15_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_ess_7_LC_22_15_7 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_CH2data_ess_7_LC_22_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_ess_7_LC_22_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__92126),
            .lcout(side_command_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94317),
            .ce(N__85264),
            .sr(N__86402));
    defparam \pid_side.error_cry_3_0_c_RNIS6493_LC_22_16_0 .C_ON=1'b0;
    defparam \pid_side.error_cry_3_0_c_RNIS6493_LC_22_16_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_3_0_c_RNIS6493_LC_22_16_0 .LUT_INIT=16'b0100000001001100;
    LogicCell40 \pid_side.error_cry_3_0_c_RNIS6493_LC_22_16_0  (
            .in0(N__85232),
            .in1(N__85069),
            .in2(N__89508),
            .in3(N__84911),
            .lcout(\pid_side.N_226 ),
            .ltout(\pid_side.N_226_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_3_19_LC_22_16_1 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_3_19_LC_22_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_3_19_LC_22_16_1 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_3_19_LC_22_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__84853),
            .in3(N__87674),
            .lcout(),
            .ltout(\pid_side.N_459_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_19_LC_22_16_2 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_19_LC_22_16_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_19_LC_22_16_2 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_19_LC_22_16_2  (
            .in0(N__88881),
            .in1(N__87601),
            .in2(N__87565),
            .in3(N__87550),
            .lcout(\pid_side.m23_2_03_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_4_19_LC_22_16_3 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_4_19_LC_22_16_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_4_19_LC_22_16_3 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_4_19_LC_22_16_3  (
            .in0(N__89818),
            .in1(N__87461),
            .in2(N__87404),
            .in3(N__85783),
            .lcout(),
            .ltout(\pid_side.m23_2_03_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_1_19_LC_22_16_4 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_1_19_LC_22_16_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_1_19_LC_22_16_4 .LUT_INIT=16'b0010101000001000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_1_19_LC_22_16_4  (
            .in0(N__87105),
            .in1(N__87165),
            .in2(N__87169),
            .in3(N__87153),
            .lcout(\pid_side.error_i_reg_esr_RNO_1Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_2_19_LC_22_16_5 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_2_19_LC_22_16_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_2_19_LC_22_16_5 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_2_19_LC_22_16_5  (
            .in0(N__87166),
            .in1(_gnd_net_),
            .in2(N__87157),
            .in3(N__87106),
            .lcout(),
            .ltout(\pid_side.error_i_reg_esr_RNO_2Z0Z_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_19_LC_22_16_6 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_19_LC_22_16_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_19_LC_22_16_6 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \pid_side.error_i_reg_esr_19_LC_22_16_6  (
            .in0(_gnd_net_),
            .in1(N__86812),
            .in2(N__86806),
            .in3(N__86803),
            .lcout(\pid_side.error_i_regZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94333),
            .ce(N__86778),
            .sr(N__86392));
    defparam \pid_side.error_i_reg_esr_RNO_5_19_LC_22_16_7 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_5_19_LC_22_16_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_5_19_LC_22_16_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_5_19_LC_22_16_7  (
            .in0(_gnd_net_),
            .in1(N__89468),
            .in2(_gnd_net_),
            .in3(N__85860),
            .lcout(\pid_side.N_622 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_3_18_LC_22_17_7 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_3_18_LC_22_17_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_3_18_LC_22_17_7 .LUT_INIT=16'b1000100011111000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_3_18_LC_22_17_7  (
            .in0(N__85771),
            .in1(N__85592),
            .in2(N__85566),
            .in3(N__85549),
            .lcout(\pid_side.m22_2_03_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.m23_2_03_0_a2_3_1_LC_22_18_7 .C_ON=1'b0;
    defparam \pid_front.m23_2_03_0_a2_3_1_LC_22_18_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.m23_2_03_0_a2_3_1_LC_22_18_7 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \pid_front.m23_2_03_0_a2_3_1_LC_22_18_7  (
            .in0(N__89817),
            .in1(N__89495),
            .in2(N__89311),
            .in3(N__88972),
            .lcout(pid_front_N_463_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kd_4_LC_22_19_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kd_4_LC_22_19_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kd_4_LC_22_19_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_xy_kd_4_LC_22_19_2  (
            .in0(_gnd_net_),
            .in1(N__88859),
            .in2(_gnd_net_),
            .in3(N__93157),
            .lcout(xy_kd_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94370),
            .ce(N__91917),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kd_5_LC_22_20_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kd_5_LC_22_20_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kd_5_LC_22_20_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \Commands_frame_decoder.source_xy_kd_5_LC_22_20_2  (
            .in0(N__88699),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__93158),
            .lcout(xy_kd_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94378),
            .ce(N__91924),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kd_6_LC_22_21_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kd_6_LC_22_21_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kd_6_LC_22_21_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_xy_kd_6_LC_22_21_2  (
            .in0(_gnd_net_),
            .in1(N__88508),
            .in2(_gnd_net_),
            .in3(N__93160),
            .lcout(xy_kd_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94387),
            .ce(N__91936),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kd_0_LC_22_21_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kd_0_LC_22_21_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kd_0_LC_22_21_4 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \Commands_frame_decoder.source_xy_kd_0_LC_22_21_4  (
            .in0(N__88320),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__93159),
            .lcout(xy_kd_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94387),
            .ce(N__91936),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_18_LC_23_7_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_18_LC_23_7_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_18_LC_23_7_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_18_LC_23_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__92755),
            .lcout(\pid_side.error_d_reg_prevZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94202),
            .ce(N__88091),
            .sr(N__87954));
    defparam \pid_side.error_d_reg_esr_4_LC_23_8_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_4_LC_23_8_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_4_LC_23_8_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_4_LC_23_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__87898),
            .lcout(\pid_side.error_d_regZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94219),
            .ce(N__92682),
            .sr(N__92986));
    defparam \pid_side.error_d_reg_prev_esr_RNIH7JO_0_18_LC_23_9_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIH7JO_0_18_LC_23_9_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIH7JO_0_18_LC_23_9_4 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIH7JO_0_18_LC_23_9_4  (
            .in0(N__90744),
            .in1(N__87867),
            .in2(_gnd_net_),
            .in3(N__92747),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIH7JO_0Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_8_LC_23_10_2 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_8_LC_23_10_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_8_LC_23_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_8_LC_23_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__87835),
            .lcout(\pid_side.error_p_regZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94251),
            .ce(N__92661),
            .sr(N__92993));
    defparam \pid_side.error_p_reg_esr_1_LC_23_11_0 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_1_LC_23_11_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_1_LC_23_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_1_LC_23_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__90727),
            .lcout(\pid_side.error_p_regZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94269),
            .ce(N__92672),
            .sr(N__92996));
    defparam \pid_front.m24_2_03_0_a2_0_0_LC_23_14_4 .C_ON=1'b0;
    defparam \pid_front.m24_2_03_0_a2_0_0_LC_23_14_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.m24_2_03_0_a2_0_0_LC_23_14_4 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \pid_front.m24_2_03_0_a2_0_0_LC_23_14_4  (
            .in0(N__90663),
            .in1(N__90433),
            .in2(_gnd_net_),
            .in3(N__90126),
            .lcout(pid_side_m24_2_03_0_a2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_16_LC_24_9_0 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_16_LC_24_9_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_16_LC_24_9_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_p_reg_esr_16_LC_24_9_0  (
            .in0(N__90055),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_p_regZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94252),
            .ce(N__92683),
            .sr(N__92994));
    defparam \pid_side.error_p_reg_esr_6_LC_24_9_1 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_6_LC_24_9_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_6_LC_24_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_6_LC_24_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__90025),
            .lcout(\pid_side.error_p_regZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94252),
            .ce(N__92683),
            .sr(N__92994));
    defparam \pid_side.error_p_reg_esr_7_LC_24_9_2 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_7_LC_24_9_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_7_LC_24_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_7_LC_24_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__89980),
            .lcout(\pid_side.error_p_regZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94252),
            .ce(N__92683),
            .sr(N__92994));
    defparam \pid_side.error_p_reg_esr_9_LC_24_9_4 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_9_LC_24_9_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_9_LC_24_9_4 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \pid_side.error_p_reg_esr_9_LC_24_9_4  (
            .in0(_gnd_net_),
            .in1(N__89950),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_p_regZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94252),
            .ce(N__92683),
            .sr(N__92994));
    defparam \pid_side.error_p_reg_esr_5_LC_24_9_6 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_5_LC_24_9_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_5_LC_24_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_5_LC_24_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__89917),
            .lcout(\pid_side.error_p_regZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94252),
            .ce(N__92683),
            .sr(N__92994));
    defparam \pid_side.error_p_reg_esr_0_LC_24_10_0 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_0_LC_24_10_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_0_LC_24_10_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_p_reg_esr_0_LC_24_10_0  (
            .in0(N__89884),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_p_regZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94270),
            .ce(N__92677),
            .sr(N__92997));
    defparam \pid_side.error_p_reg_esr_19_LC_24_10_1 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_19_LC_24_10_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_19_LC_24_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_19_LC_24_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__91060),
            .lcout(\pid_side.error_p_regZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94270),
            .ce(N__92677),
            .sr(N__92997));
    defparam \pid_side.error_p_reg_esr_11_LC_24_10_3 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_11_LC_24_10_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_11_LC_24_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_11_LC_24_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__91033),
            .lcout(\pid_side.error_p_regZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94270),
            .ce(N__92677),
            .sr(N__92997));
    defparam \pid_side.error_p_reg_esr_12_LC_24_10_4 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_12_LC_24_10_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_12_LC_24_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_12_LC_24_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__90991),
            .lcout(\pid_side.error_p_regZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94270),
            .ce(N__92677),
            .sr(N__92997));
    defparam \pid_side.error_p_reg_esr_13_LC_24_10_5 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_13_LC_24_10_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_13_LC_24_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_13_LC_24_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__90931),
            .lcout(\pid_side.error_p_regZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94270),
            .ce(N__92677),
            .sr(N__92997));
    defparam \pid_side.error_p_reg_esr_14_LC_24_10_6 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_14_LC_24_10_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_14_LC_24_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_14_LC_24_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__90865),
            .lcout(\pid_side.error_p_regZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94270),
            .ce(N__92677),
            .sr(N__92997));
    defparam \pid_side.error_p_reg_esr_15_LC_24_10_7 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_15_LC_24_10_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_15_LC_24_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_15_LC_24_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__90823),
            .lcout(\pid_side.error_p_regZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94270),
            .ce(N__92677),
            .sr(N__92997));
    defparam \pid_side.error_p_reg_esr_17_LC_24_11_1 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_17_LC_24_11_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_17_LC_24_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_17_LC_24_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__90796),
            .lcout(\pid_side.error_p_regZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94286),
            .ce(N__92649),
            .sr(N__92998));
    defparam \pid_side.error_p_reg_esr_18_LC_24_11_2 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_18_LC_24_11_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_18_LC_24_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_18_LC_24_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__90754),
            .lcout(\pid_side.error_p_regZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94286),
            .ce(N__92649),
            .sr(N__92998));
    defparam \pid_side.error_p_reg_esr_20_LC_24_11_5 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_20_LC_24_11_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_20_LC_24_11_5 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \pid_side.error_p_reg_esr_20_LC_24_11_5  (
            .in0(_gnd_net_),
            .in1(N__91660),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_p_regZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94286),
            .ce(N__92649),
            .sr(N__92998));
    defparam \pid_side.error_d_reg_esr_15_LC_24_13_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_15_LC_24_13_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_15_LC_24_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_15_LC_24_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__91552),
            .lcout(\pid_side.error_d_regZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94318),
            .ce(N__92665),
            .sr(N__93000));
    defparam \pid_side.error_d_reg_esr_13_LC_24_13_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_13_LC_24_13_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_13_LC_24_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_13_LC_24_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__91518),
            .lcout(\pid_side.error_d_regZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94318),
            .ce(N__92665),
            .sr(N__93000));
    defparam \pid_side.error_d_reg_esr_14_LC_24_14_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_14_LC_24_14_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_14_LC_24_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_14_LC_24_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__91453),
            .lcout(\pid_side.error_d_regZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94334),
            .ce(N__92676),
            .sr(N__93001));
    defparam \pid_side.error_d_reg_esr_21_LC_24_14_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_21_LC_24_14_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_21_LC_24_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_21_LC_24_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__91396),
            .lcout(\pid_side.error_d_regZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94334),
            .ce(N__92676),
            .sr(N__93001));
    defparam \pid_side.error_d_reg_esr_12_LC_24_14_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_12_LC_24_14_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_12_LC_24_14_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_esr_12_LC_24_14_2  (
            .in0(N__91263),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_regZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94334),
            .ce(N__92676),
            .sr(N__93001));
    defparam \pid_side.error_d_reg_esr_17_LC_24_14_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_17_LC_24_14_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_17_LC_24_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_17_LC_24_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__91183),
            .lcout(\pid_side.error_d_regZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94334),
            .ce(N__92676),
            .sr(N__93001));
    defparam \pid_side.error_d_reg_esr_19_LC_24_14_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_19_LC_24_14_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_19_LC_24_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_19_LC_24_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__91141),
            .lcout(\pid_side.error_d_regZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94334),
            .ce(N__92676),
            .sr(N__93001));
    defparam \pid_side.error_d_reg_esr_20_LC_24_14_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_20_LC_24_14_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_20_LC_24_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_20_LC_24_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__91099),
            .lcout(\pid_side.error_d_regZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94334),
            .ce(N__92676),
            .sr(N__93001));
    defparam \pid_side.error_d_reg_esr_18_LC_24_15_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_18_LC_24_15_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_18_LC_24_15_2 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \pid_side.error_d_reg_esr_18_LC_24_15_2  (
            .in0(_gnd_net_),
            .in1(N__92764),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_regZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94348),
            .ce(N__92650),
            .sr(N__93002));
    defparam \pid_side.error_d_reg_esr_16_LC_24_15_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_16_LC_24_15_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_16_LC_24_15_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_esr_16_LC_24_15_7  (
            .in0(N__92719),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_regZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94348),
            .ce(N__92650),
            .sr(N__93002));
    defparam \Commands_frame_decoder.source_xy_kd_2_LC_24_20_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kd_2_LC_24_20_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kd_2_LC_24_20_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_xy_kd_2_LC_24_20_1  (
            .in0(_gnd_net_),
            .in1(N__92519),
            .in2(_gnd_net_),
            .in3(N__93161),
            .lcout(xy_kd_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94393),
            .ce(N__91932),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kd_3_LC_24_20_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kd_3_LC_24_20_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kd_3_LC_24_20_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_xy_kd_3_LC_24_20_3  (
            .in0(_gnd_net_),
            .in1(N__92332),
            .in2(_gnd_net_),
            .in3(N__93162),
            .lcout(xy_kd_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94393),
            .ce(N__91932),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kd_7_LC_24_20_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kd_7_LC_24_20_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kd_7_LC_24_20_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_kd_7_LC_24_20_4  (
            .in0(N__93163),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__92125),
            .lcout(xy_kd_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94393),
            .ce(N__91932),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_esr_20_LC_24_22_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_20_LC_24_22_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_20_LC_24_22_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_20_LC_24_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__91870),
            .lcout(\pid_front.error_d_regZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94402),
            .ce(N__93332),
            .sr(N__93013));
    defparam \pid_front.error_d_reg_esr_19_LC_24_23_0 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_19_LC_24_23_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_19_LC_24_23_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_19_LC_24_23_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__91828),
            .lcout(\pid_front.error_d_regZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94407),
            .ce(N__93407),
            .sr(N__93015));
    defparam \pid_front.error_d_reg_esr_21_LC_24_23_2 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_21_LC_24_23_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_21_LC_24_23_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_21_LC_24_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__91789),
            .lcout(\pid_front.error_d_regZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94407),
            .ce(N__93407),
            .sr(N__93015));
    defparam \pid_front.error_d_reg_esr_5_LC_24_23_4 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_5_LC_24_23_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_5_LC_24_23_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_5_LC_24_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__94687),
            .lcout(\pid_front.error_d_regZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94407),
            .ce(N__93407),
            .sr(N__93015));
    defparam \pid_front.error_d_reg_esr_7_LC_24_23_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_7_LC_24_23_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_7_LC_24_23_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_7_LC_24_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__94624),
            .lcout(\pid_front.error_d_regZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94407),
            .ce(N__93407),
            .sr(N__93015));
    defparam \pid_front.error_d_reg_esr_11_LC_24_24_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_11_LC_24_24_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_11_LC_24_24_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_11_LC_24_24_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__94597),
            .lcout(\pid_front.error_d_regZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94410),
            .ce(N__93408),
            .sr(N__93016));
    defparam \pid_front.error_d_reg_esr_14_LC_24_24_4 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_14_LC_24_24_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_14_LC_24_24_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_14_LC_24_24_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__94546),
            .lcout(\pid_front.error_d_regZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94410),
            .ce(N__93408),
            .sr(N__93016));
    defparam \pid_front.error_d_reg_esr_15_LC_24_24_5 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_15_LC_24_24_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_15_LC_24_24_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_15_LC_24_24_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__94501),
            .lcout(\pid_front.error_d_regZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94410),
            .ce(N__93408),
            .sr(N__93016));
    defparam \pid_front.error_d_reg_esr_16_LC_24_24_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_16_LC_24_24_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_16_LC_24_24_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_16_LC_24_24_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__94471),
            .lcout(\pid_front.error_d_regZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94410),
            .ce(N__93408),
            .sr(N__93016));
    defparam \pid_front.error_d_reg_esr_17_LC_24_24_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_17_LC_24_24_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_17_LC_24_24_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_17_LC_24_24_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__94441),
            .lcout(\pid_front.error_d_regZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__94410),
            .ce(N__93408),
            .sr(N__93016));
endmodule // Pc2drone
