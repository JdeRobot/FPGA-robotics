-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     Mar 13 2019 00:12:36

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "Pc2Drone" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of Pc2Drone
entity Pc2Drone is
port (
    debug_state_output : out std_logic_vector(4 downto 0);
    uart_input : in std_logic;
    uart_data_rdy : out std_logic;
    debug_sinkdatavalid_output : out std_logic;
    uart_input_debug : out std_logic;
    frame_decoder_dv : out std_logic;
    clk_system : in std_logic);
end Pc2Drone;

-- Architecture of Pc2Drone
-- View name is \INTERFACE\
architecture \INTERFACE\ of Pc2Drone is

signal \N__5663\ : std_logic;
signal \N__5662\ : std_logic;
signal \N__5661\ : std_logic;
signal \N__5652\ : std_logic;
signal \N__5651\ : std_logic;
signal \N__5650\ : std_logic;
signal \N__5643\ : std_logic;
signal \N__5642\ : std_logic;
signal \N__5641\ : std_logic;
signal \N__5634\ : std_logic;
signal \N__5633\ : std_logic;
signal \N__5632\ : std_logic;
signal \N__5625\ : std_logic;
signal \N__5624\ : std_logic;
signal \N__5623\ : std_logic;
signal \N__5616\ : std_logic;
signal \N__5615\ : std_logic;
signal \N__5614\ : std_logic;
signal \N__5607\ : std_logic;
signal \N__5606\ : std_logic;
signal \N__5605\ : std_logic;
signal \N__5598\ : std_logic;
signal \N__5597\ : std_logic;
signal \N__5596\ : std_logic;
signal \N__5589\ : std_logic;
signal \N__5588\ : std_logic;
signal \N__5587\ : std_logic;
signal \N__5580\ : std_logic;
signal \N__5579\ : std_logic;
signal \N__5578\ : std_logic;
signal \N__5571\ : std_logic;
signal \N__5570\ : std_logic;
signal \N__5569\ : std_logic;
signal \N__5552\ : std_logic;
signal \N__5551\ : std_logic;
signal \N__5550\ : std_logic;
signal \N__5549\ : std_logic;
signal \N__5546\ : std_logic;
signal \N__5543\ : std_logic;
signal \N__5540\ : std_logic;
signal \N__5537\ : std_logic;
signal \N__5536\ : std_logic;
signal \N__5533\ : std_logic;
signal \N__5530\ : std_logic;
signal \N__5527\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5521\ : std_logic;
signal \N__5518\ : std_logic;
signal \N__5511\ : std_logic;
signal \N__5504\ : std_logic;
signal \N__5503\ : std_logic;
signal \N__5502\ : std_logic;
signal \N__5501\ : std_logic;
signal \N__5498\ : std_logic;
signal \N__5497\ : std_logic;
signal \N__5496\ : std_logic;
signal \N__5495\ : std_logic;
signal \N__5494\ : std_logic;
signal \N__5493\ : std_logic;
signal \N__5492\ : std_logic;
signal \N__5491\ : std_logic;
signal \N__5488\ : std_logic;
signal \N__5485\ : std_logic;
signal \N__5482\ : std_logic;
signal \N__5479\ : std_logic;
signal \N__5464\ : std_logic;
signal \N__5461\ : std_logic;
signal \N__5460\ : std_logic;
signal \N__5459\ : std_logic;
signal \N__5458\ : std_logic;
signal \N__5457\ : std_logic;
signal \N__5456\ : std_logic;
signal \N__5455\ : std_logic;
signal \N__5450\ : std_logic;
signal \N__5445\ : std_logic;
signal \N__5444\ : std_logic;
signal \N__5443\ : std_logic;
signal \N__5440\ : std_logic;
signal \N__5437\ : std_logic;
signal \N__5432\ : std_logic;
signal \N__5427\ : std_logic;
signal \N__5424\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5422\ : std_logic;
signal \N__5419\ : std_logic;
signal \N__5416\ : std_logic;
signal \N__5411\ : std_logic;
signal \N__5406\ : std_logic;
signal \N__5401\ : std_logic;
signal \N__5398\ : std_logic;
signal \N__5393\ : std_logic;
signal \N__5378\ : std_logic;
signal \N__5377\ : std_logic;
signal \N__5376\ : std_logic;
signal \N__5373\ : std_logic;
signal \N__5372\ : std_logic;
signal \N__5369\ : std_logic;
signal \N__5368\ : std_logic;
signal \N__5365\ : std_logic;
signal \N__5364\ : std_logic;
signal \N__5363\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5361\ : std_logic;
signal \N__5360\ : std_logic;
signal \N__5359\ : std_logic;
signal \N__5358\ : std_logic;
signal \N__5355\ : std_logic;
signal \N__5352\ : std_logic;
signal \N__5349\ : std_logic;
signal \N__5346\ : std_logic;
signal \N__5343\ : std_logic;
signal \N__5338\ : std_logic;
signal \N__5331\ : std_logic;
signal \N__5328\ : std_logic;
signal \N__5325\ : std_logic;
signal \N__5318\ : std_logic;
signal \N__5309\ : std_logic;
signal \N__5300\ : std_logic;
signal \N__5297\ : std_logic;
signal \N__5296\ : std_logic;
signal \N__5293\ : std_logic;
signal \N__5290\ : std_logic;
signal \N__5287\ : std_logic;
signal \N__5284\ : std_logic;
signal \N__5279\ : std_logic;
signal \N__5278\ : std_logic;
signal \N__5275\ : std_logic;
signal \N__5274\ : std_logic;
signal \N__5271\ : std_logic;
signal \N__5266\ : std_logic;
signal \N__5261\ : std_logic;
signal \N__5258\ : std_logic;
signal \N__5255\ : std_logic;
signal \N__5252\ : std_logic;
signal \N__5249\ : std_logic;
signal \N__5246\ : std_logic;
signal \N__5245\ : std_logic;
signal \N__5244\ : std_logic;
signal \N__5241\ : std_logic;
signal \N__5238\ : std_logic;
signal \N__5233\ : std_logic;
signal \N__5228\ : std_logic;
signal \N__5225\ : std_logic;
signal \N__5222\ : std_logic;
signal \N__5219\ : std_logic;
signal \N__5216\ : std_logic;
signal \N__5215\ : std_logic;
signal \N__5212\ : std_logic;
signal \N__5211\ : std_logic;
signal \N__5208\ : std_logic;
signal \N__5207\ : std_logic;
signal \N__5206\ : std_logic;
signal \N__5203\ : std_logic;
signal \N__5200\ : std_logic;
signal \N__5197\ : std_logic;
signal \N__5192\ : std_logic;
signal \N__5183\ : std_logic;
signal \N__5182\ : std_logic;
signal \N__5181\ : std_logic;
signal \N__5180\ : std_logic;
signal \N__5177\ : std_logic;
signal \N__5172\ : std_logic;
signal \N__5167\ : std_logic;
signal \N__5162\ : std_logic;
signal \N__5159\ : std_logic;
signal \N__5158\ : std_logic;
signal \N__5157\ : std_logic;
signal \N__5154\ : std_logic;
signal \N__5153\ : std_logic;
signal \N__5148\ : std_logic;
signal \N__5143\ : std_logic;
signal \N__5138\ : std_logic;
signal \N__5135\ : std_logic;
signal \N__5132\ : std_logic;
signal \N__5129\ : std_logic;
signal \N__5126\ : std_logic;
signal \N__5123\ : std_logic;
signal \N__5122\ : std_logic;
signal \N__5119\ : std_logic;
signal \N__5118\ : std_logic;
signal \N__5115\ : std_logic;
signal \N__5110\ : std_logic;
signal \N__5105\ : std_logic;
signal \N__5104\ : std_logic;
signal \N__5103\ : std_logic;
signal \N__5102\ : std_logic;
signal \N__5099\ : std_logic;
signal \N__5094\ : std_logic;
signal \N__5089\ : std_logic;
signal \N__5084\ : std_logic;
signal \N__5081\ : std_logic;
signal \N__5078\ : std_logic;
signal \N__5075\ : std_logic;
signal \N__5074\ : std_logic;
signal \N__5073\ : std_logic;
signal \N__5070\ : std_logic;
signal \N__5067\ : std_logic;
signal \N__5064\ : std_logic;
signal \N__5057\ : std_logic;
signal \N__5056\ : std_logic;
signal \N__5055\ : std_logic;
signal \N__5052\ : std_logic;
signal \N__5051\ : std_logic;
signal \N__5046\ : std_logic;
signal \N__5041\ : std_logic;
signal \N__5036\ : std_logic;
signal \N__5033\ : std_logic;
signal \N__5032\ : std_logic;
signal \N__5031\ : std_logic;
signal \N__5030\ : std_logic;
signal \N__5027\ : std_logic;
signal \N__5026\ : std_logic;
signal \N__5021\ : std_logic;
signal \N__5018\ : std_logic;
signal \N__5017\ : std_logic;
signal \N__5014\ : std_logic;
signal \N__5011\ : std_logic;
signal \N__5010\ : std_logic;
signal \N__5009\ : std_logic;
signal \N__5008\ : std_logic;
signal \N__5003\ : std_logic;
signal \N__5000\ : std_logic;
signal \N__4995\ : std_logic;
signal \N__4990\ : std_logic;
signal \N__4987\ : std_logic;
signal \N__4982\ : std_logic;
signal \N__4979\ : std_logic;
signal \N__4970\ : std_logic;
signal \N__4967\ : std_logic;
signal \N__4964\ : std_logic;
signal \N__4961\ : std_logic;
signal \N__4958\ : std_logic;
signal \N__4955\ : std_logic;
signal \N__4954\ : std_logic;
signal \N__4953\ : std_logic;
signal \N__4950\ : std_logic;
signal \N__4947\ : std_logic;
signal \N__4942\ : std_logic;
signal \N__4937\ : std_logic;
signal \N__4934\ : std_logic;
signal \N__4931\ : std_logic;
signal \N__4928\ : std_logic;
signal \N__4927\ : std_logic;
signal \N__4924\ : std_logic;
signal \N__4921\ : std_logic;
signal \N__4916\ : std_logic;
signal \N__4915\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4913\ : std_logic;
signal \N__4912\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4910\ : std_logic;
signal \N__4909\ : std_logic;
signal \N__4908\ : std_logic;
signal \N__4893\ : std_logic;
signal \N__4888\ : std_logic;
signal \N__4883\ : std_logic;
signal \N__4882\ : std_logic;
signal \N__4881\ : std_logic;
signal \N__4880\ : std_logic;
signal \N__4879\ : std_logic;
signal \N__4878\ : std_logic;
signal \N__4877\ : std_logic;
signal \N__4876\ : std_logic;
signal \N__4875\ : std_logic;
signal \N__4874\ : std_logic;
signal \N__4873\ : std_logic;
signal \N__4872\ : std_logic;
signal \N__4871\ : std_logic;
signal \N__4870\ : std_logic;
signal \N__4869\ : std_logic;
signal \N__4868\ : std_logic;
signal \N__4867\ : std_logic;
signal \N__4866\ : std_logic;
signal \N__4865\ : std_logic;
signal \N__4864\ : std_logic;
signal \N__4863\ : std_logic;
signal \N__4862\ : std_logic;
signal \N__4861\ : std_logic;
signal \N__4860\ : std_logic;
signal \N__4859\ : std_logic;
signal \N__4808\ : std_logic;
signal \N__4805\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4801\ : std_logic;
signal \N__4800\ : std_logic;
signal \N__4797\ : std_logic;
signal \N__4794\ : std_logic;
signal \N__4791\ : std_logic;
signal \N__4784\ : std_logic;
signal \N__4781\ : std_logic;
signal \N__4780\ : std_logic;
signal \N__4779\ : std_logic;
signal \N__4776\ : std_logic;
signal \N__4773\ : std_logic;
signal \N__4770\ : std_logic;
signal \N__4767\ : std_logic;
signal \N__4764\ : std_logic;
signal \N__4757\ : std_logic;
signal \N__4754\ : std_logic;
signal \N__4753\ : std_logic;
signal \N__4752\ : std_logic;
signal \N__4749\ : std_logic;
signal \N__4746\ : std_logic;
signal \N__4743\ : std_logic;
signal \N__4736\ : std_logic;
signal \N__4733\ : std_logic;
signal \N__4732\ : std_logic;
signal \N__4731\ : std_logic;
signal \N__4728\ : std_logic;
signal \N__4727\ : std_logic;
signal \N__4724\ : std_logic;
signal \N__4719\ : std_logic;
signal \N__4716\ : std_logic;
signal \N__4709\ : std_logic;
signal \N__4706\ : std_logic;
signal \N__4705\ : std_logic;
signal \N__4704\ : std_logic;
signal \N__4701\ : std_logic;
signal \N__4698\ : std_logic;
signal \N__4695\ : std_logic;
signal \N__4688\ : std_logic;
signal \N__4685\ : std_logic;
signal \N__4684\ : std_logic;
signal \N__4683\ : std_logic;
signal \N__4680\ : std_logic;
signal \N__4677\ : std_logic;
signal \N__4674\ : std_logic;
signal \N__4667\ : std_logic;
signal \N__4664\ : std_logic;
signal \N__4663\ : std_logic;
signal \N__4662\ : std_logic;
signal \N__4661\ : std_logic;
signal \N__4658\ : std_logic;
signal \N__4655\ : std_logic;
signal \N__4648\ : std_logic;
signal \N__4643\ : std_logic;
signal \N__4640\ : std_logic;
signal \N__4639\ : std_logic;
signal \N__4634\ : std_logic;
signal \N__4633\ : std_logic;
signal \N__4632\ : std_logic;
signal \N__4631\ : std_logic;
signal \N__4630\ : std_logic;
signal \N__4627\ : std_logic;
signal \N__4624\ : std_logic;
signal \N__4617\ : std_logic;
signal \N__4614\ : std_logic;
signal \N__4607\ : std_logic;
signal \N__4604\ : std_logic;
signal \N__4601\ : std_logic;
signal \N__4600\ : std_logic;
signal \N__4597\ : std_logic;
signal \N__4594\ : std_logic;
signal \N__4591\ : std_logic;
signal \N__4588\ : std_logic;
signal \N__4583\ : std_logic;
signal \N__4580\ : std_logic;
signal \N__4577\ : std_logic;
signal \N__4574\ : std_logic;
signal \N__4571\ : std_logic;
signal \N__4570\ : std_logic;
signal \N__4567\ : std_logic;
signal \N__4564\ : std_logic;
signal \N__4559\ : std_logic;
signal \N__4556\ : std_logic;
signal \N__4553\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4547\ : std_logic;
signal \N__4546\ : std_logic;
signal \N__4543\ : std_logic;
signal \N__4540\ : std_logic;
signal \N__4537\ : std_logic;
signal \N__4534\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4528\ : std_logic;
signal \N__4525\ : std_logic;
signal \N__4522\ : std_logic;
signal \N__4519\ : std_logic;
signal \N__4516\ : std_logic;
signal \N__4515\ : std_logic;
signal \N__4512\ : std_logic;
signal \N__4509\ : std_logic;
signal \N__4506\ : std_logic;
signal \N__4499\ : std_logic;
signal \N__4498\ : std_logic;
signal \N__4495\ : std_logic;
signal \N__4492\ : std_logic;
signal \N__4489\ : std_logic;
signal \N__4486\ : std_logic;
signal \N__4481\ : std_logic;
signal \N__4478\ : std_logic;
signal \N__4475\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4469\ : std_logic;
signal \N__4466\ : std_logic;
signal \N__4463\ : std_logic;
signal \N__4460\ : std_logic;
signal \N__4457\ : std_logic;
signal \N__4454\ : std_logic;
signal \N__4451\ : std_logic;
signal \N__4448\ : std_logic;
signal \N__4447\ : std_logic;
signal \N__4446\ : std_logic;
signal \N__4443\ : std_logic;
signal \N__4438\ : std_logic;
signal \N__4433\ : std_logic;
signal \N__4430\ : std_logic;
signal \N__4427\ : std_logic;
signal \N__4426\ : std_logic;
signal \N__4425\ : std_logic;
signal \N__4422\ : std_logic;
signal \N__4419\ : std_logic;
signal \N__4416\ : std_logic;
signal \N__4413\ : std_logic;
signal \N__4406\ : std_logic;
signal \N__4403\ : std_logic;
signal \N__4402\ : std_logic;
signal \N__4401\ : std_logic;
signal \N__4398\ : std_logic;
signal \N__4395\ : std_logic;
signal \N__4392\ : std_logic;
signal \N__4389\ : std_logic;
signal \N__4382\ : std_logic;
signal \N__4379\ : std_logic;
signal \N__4376\ : std_logic;
signal \N__4373\ : std_logic;
signal \N__4370\ : std_logic;
signal \N__4367\ : std_logic;
signal \N__4364\ : std_logic;
signal \N__4361\ : std_logic;
signal \N__4358\ : std_logic;
signal \N__4357\ : std_logic;
signal \N__4352\ : std_logic;
signal \N__4349\ : std_logic;
signal \N__4346\ : std_logic;
signal \N__4345\ : std_logic;
signal \N__4342\ : std_logic;
signal \N__4339\ : std_logic;
signal \N__4334\ : std_logic;
signal \N__4331\ : std_logic;
signal \N__4328\ : std_logic;
signal \N__4325\ : std_logic;
signal \N__4324\ : std_logic;
signal \N__4321\ : std_logic;
signal \N__4320\ : std_logic;
signal \N__4319\ : std_logic;
signal \N__4316\ : std_logic;
signal \N__4313\ : std_logic;
signal \N__4308\ : std_logic;
signal \N__4305\ : std_logic;
signal \N__4302\ : std_logic;
signal \N__4295\ : std_logic;
signal \N__4294\ : std_logic;
signal \N__4291\ : std_logic;
signal \N__4288\ : std_logic;
signal \N__4283\ : std_logic;
signal \N__4280\ : std_logic;
signal \N__4277\ : std_logic;
signal \N__4274\ : std_logic;
signal \N__4271\ : std_logic;
signal \N__4270\ : std_logic;
signal \N__4269\ : std_logic;
signal \N__4264\ : std_logic;
signal \N__4261\ : std_logic;
signal \N__4256\ : std_logic;
signal \N__4255\ : std_logic;
signal \N__4252\ : std_logic;
signal \N__4249\ : std_logic;
signal \N__4244\ : std_logic;
signal \N__4241\ : std_logic;
signal \N__4240\ : std_logic;
signal \N__4237\ : std_logic;
signal \N__4234\ : std_logic;
signal \N__4231\ : std_logic;
signal \N__4228\ : std_logic;
signal \N__4223\ : std_logic;
signal \N__4220\ : std_logic;
signal \N__4217\ : std_logic;
signal \N__4214\ : std_logic;
signal \N__4211\ : std_logic;
signal \N__4208\ : std_logic;
signal \N__4205\ : std_logic;
signal \N__4202\ : std_logic;
signal \N__4199\ : std_logic;
signal \N__4196\ : std_logic;
signal \N__4193\ : std_logic;
signal \N__4190\ : std_logic;
signal \N__4187\ : std_logic;
signal \N__4184\ : std_logic;
signal \N__4183\ : std_logic;
signal \N__4182\ : std_logic;
signal \N__4179\ : std_logic;
signal \N__4174\ : std_logic;
signal \N__4169\ : std_logic;
signal \N__4166\ : std_logic;
signal \N__4163\ : std_logic;
signal \N__4160\ : std_logic;
signal \N__4157\ : std_logic;
signal \N__4156\ : std_logic;
signal \N__4155\ : std_logic;
signal \N__4152\ : std_logic;
signal \N__4149\ : std_logic;
signal \N__4148\ : std_logic;
signal \N__4145\ : std_logic;
signal \N__4142\ : std_logic;
signal \N__4139\ : std_logic;
signal \N__4136\ : std_logic;
signal \N__4127\ : std_logic;
signal \N__4124\ : std_logic;
signal \N__4121\ : std_logic;
signal \N__4118\ : std_logic;
signal \N__4115\ : std_logic;
signal \N__4112\ : std_logic;
signal \N__4109\ : std_logic;
signal \N__4106\ : std_logic;
signal \N__4103\ : std_logic;
signal \N__4100\ : std_logic;
signal \N__4097\ : std_logic;
signal \N__4094\ : std_logic;
signal \N__4093\ : std_logic;
signal \N__4088\ : std_logic;
signal \N__4085\ : std_logic;
signal \N__4082\ : std_logic;
signal \N__4081\ : std_logic;
signal \N__4080\ : std_logic;
signal \N__4077\ : std_logic;
signal \N__4076\ : std_logic;
signal \N__4071\ : std_logic;
signal \N__4066\ : std_logic;
signal \N__4061\ : std_logic;
signal \N__4060\ : std_logic;
signal \N__4059\ : std_logic;
signal \N__4056\ : std_logic;
signal \N__4051\ : std_logic;
signal \N__4046\ : std_logic;
signal \N__4045\ : std_logic;
signal \N__4040\ : std_logic;
signal \N__4037\ : std_logic;
signal \N__4036\ : std_logic;
signal \N__4035\ : std_logic;
signal \N__4034\ : std_logic;
signal \N__4031\ : std_logic;
signal \N__4024\ : std_logic;
signal \N__4019\ : std_logic;
signal \N__4018\ : std_logic;
signal \N__4015\ : std_logic;
signal \N__4010\ : std_logic;
signal \N__4007\ : std_logic;
signal \N__4004\ : std_logic;
signal \N__4003\ : std_logic;
signal \N__4002\ : std_logic;
signal \N__4001\ : std_logic;
signal \N__4000\ : std_logic;
signal \N__3997\ : std_logic;
signal \N__3994\ : std_logic;
signal \N__3987\ : std_logic;
signal \N__3980\ : std_logic;
signal \N__3977\ : std_logic;
signal \N__3974\ : std_logic;
signal \N__3971\ : std_logic;
signal \N__3968\ : std_logic;
signal \N__3967\ : std_logic;
signal \N__3966\ : std_logic;
signal \N__3965\ : std_logic;
signal \N__3964\ : std_logic;
signal \N__3961\ : std_logic;
signal \N__3958\ : std_logic;
signal \N__3955\ : std_logic;
signal \N__3952\ : std_logic;
signal \N__3949\ : std_logic;
signal \N__3946\ : std_logic;
signal \N__3941\ : std_logic;
signal \N__3932\ : std_logic;
signal \N__3929\ : std_logic;
signal \N__3926\ : std_logic;
signal \N__3925\ : std_logic;
signal \N__3924\ : std_logic;
signal \N__3921\ : std_logic;
signal \N__3920\ : std_logic;
signal \N__3919\ : std_logic;
signal \N__3916\ : std_logic;
signal \N__3913\ : std_logic;
signal \N__3910\ : std_logic;
signal \N__3907\ : std_logic;
signal \N__3904\ : std_logic;
signal \N__3893\ : std_logic;
signal \N__3890\ : std_logic;
signal \N__3887\ : std_logic;
signal \N__3886\ : std_logic;
signal \N__3885\ : std_logic;
signal \N__3884\ : std_logic;
signal \N__3881\ : std_logic;
signal \N__3880\ : std_logic;
signal \N__3877\ : std_logic;
signal \N__3874\ : std_logic;
signal \N__3871\ : std_logic;
signal \N__3868\ : std_logic;
signal \N__3865\ : std_logic;
signal \N__3862\ : std_logic;
signal \N__3851\ : std_logic;
signal \N__3848\ : std_logic;
signal \N__3847\ : std_logic;
signal \N__3844\ : std_logic;
signal \N__3843\ : std_logic;
signal \N__3842\ : std_logic;
signal \N__3841\ : std_logic;
signal \N__3838\ : std_logic;
signal \N__3835\ : std_logic;
signal \N__3828\ : std_logic;
signal \N__3821\ : std_logic;
signal \N__3818\ : std_logic;
signal \N__3817\ : std_logic;
signal \N__3814\ : std_logic;
signal \N__3813\ : std_logic;
signal \N__3812\ : std_logic;
signal \N__3809\ : std_logic;
signal \N__3806\ : std_logic;
signal \N__3801\ : std_logic;
signal \N__3794\ : std_logic;
signal \N__3791\ : std_logic;
signal \N__3788\ : std_logic;
signal \N__3787\ : std_logic;
signal \N__3784\ : std_logic;
signal \N__3781\ : std_logic;
signal \N__3780\ : std_logic;
signal \N__3779\ : std_logic;
signal \N__3774\ : std_logic;
signal \N__3773\ : std_logic;
signal \N__3772\ : std_logic;
signal \N__3771\ : std_logic;
signal \N__3770\ : std_logic;
signal \N__3767\ : std_logic;
signal \N__3764\ : std_logic;
signal \N__3761\ : std_logic;
signal \N__3754\ : std_logic;
signal \N__3749\ : std_logic;
signal \N__3740\ : std_logic;
signal \N__3737\ : std_logic;
signal \N__3734\ : std_logic;
signal \N__3731\ : std_logic;
signal \N__3730\ : std_logic;
signal \N__3725\ : std_logic;
signal \N__3722\ : std_logic;
signal \N__3721\ : std_logic;
signal \N__3716\ : std_logic;
signal \N__3713\ : std_logic;
signal \N__3710\ : std_logic;
signal \N__3709\ : std_logic;
signal \N__3704\ : std_logic;
signal \N__3701\ : std_logic;
signal \N__3700\ : std_logic;
signal \N__3695\ : std_logic;
signal \N__3692\ : std_logic;
signal \N__3689\ : std_logic;
signal \N__3686\ : std_logic;
signal \N__3683\ : std_logic;
signal \N__3682\ : std_logic;
signal \N__3681\ : std_logic;
signal \N__3678\ : std_logic;
signal \N__3677\ : std_logic;
signal \N__3676\ : std_logic;
signal \N__3673\ : std_logic;
signal \N__3672\ : std_logic;
signal \N__3671\ : std_logic;
signal \N__3670\ : std_logic;
signal \N__3669\ : std_logic;
signal \N__3668\ : std_logic;
signal \N__3665\ : std_logic;
signal \N__3662\ : std_logic;
signal \N__3659\ : std_logic;
signal \N__3656\ : std_logic;
signal \N__3653\ : std_logic;
signal \N__3652\ : std_logic;
signal \N__3651\ : std_logic;
signal \N__3650\ : std_logic;
signal \N__3647\ : std_logic;
signal \N__3638\ : std_logic;
signal \N__3635\ : std_logic;
signal \N__3626\ : std_logic;
signal \N__3619\ : std_logic;
signal \N__3616\ : std_logic;
signal \N__3613\ : std_logic;
signal \N__3608\ : std_logic;
signal \N__3599\ : std_logic;
signal \N__3596\ : std_logic;
signal \N__3593\ : std_logic;
signal \N__3590\ : std_logic;
signal \N__3587\ : std_logic;
signal \N__3584\ : std_logic;
signal \N__3581\ : std_logic;
signal \N__3578\ : std_logic;
signal \N__3575\ : std_logic;
signal \N__3572\ : std_logic;
signal \N__3571\ : std_logic;
signal \N__3568\ : std_logic;
signal \N__3567\ : std_logic;
signal \N__3566\ : std_logic;
signal \N__3565\ : std_logic;
signal \N__3562\ : std_logic;
signal \N__3559\ : std_logic;
signal \N__3556\ : std_logic;
signal \N__3553\ : std_logic;
signal \N__3550\ : std_logic;
signal \N__3539\ : std_logic;
signal \N__3536\ : std_logic;
signal \N__3535\ : std_logic;
signal \N__3534\ : std_logic;
signal \N__3531\ : std_logic;
signal \N__3526\ : std_logic;
signal \N__3521\ : std_logic;
signal \N__3520\ : std_logic;
signal \N__3517\ : std_logic;
signal \N__3514\ : std_logic;
signal \N__3513\ : std_logic;
signal \N__3512\ : std_logic;
signal \N__3511\ : std_logic;
signal \N__3506\ : std_logic;
signal \N__3505\ : std_logic;
signal \N__3502\ : std_logic;
signal \N__3501\ : std_logic;
signal \N__3500\ : std_logic;
signal \N__3497\ : std_logic;
signal \N__3494\ : std_logic;
signal \N__3491\ : std_logic;
signal \N__3488\ : std_logic;
signal \N__3483\ : std_logic;
signal \N__3480\ : std_logic;
signal \N__3467\ : std_logic;
signal \N__3464\ : std_logic;
signal \N__3461\ : std_logic;
signal \N__3458\ : std_logic;
signal \N__3455\ : std_logic;
signal \N__3454\ : std_logic;
signal \N__3453\ : std_logic;
signal \N__3450\ : std_logic;
signal \N__3447\ : std_logic;
signal \N__3444\ : std_logic;
signal \N__3439\ : std_logic;
signal \N__3436\ : std_logic;
signal \N__3433\ : std_logic;
signal \N__3430\ : std_logic;
signal \N__3427\ : std_logic;
signal \N__3422\ : std_logic;
signal \N__3421\ : std_logic;
signal \N__3420\ : std_logic;
signal \N__3417\ : std_logic;
signal \N__3412\ : std_logic;
signal \N__3407\ : std_logic;
signal \N__3404\ : std_logic;
signal \N__3403\ : std_logic;
signal \N__3400\ : std_logic;
signal \N__3397\ : std_logic;
signal \N__3396\ : std_logic;
signal \N__3393\ : std_logic;
signal \N__3392\ : std_logic;
signal \N__3389\ : std_logic;
signal \N__3386\ : std_logic;
signal \N__3383\ : std_logic;
signal \N__3380\ : std_logic;
signal \N__3371\ : std_logic;
signal \N__3370\ : std_logic;
signal \N__3369\ : std_logic;
signal \N__3366\ : std_logic;
signal \N__3363\ : std_logic;
signal \N__3362\ : std_logic;
signal \N__3361\ : std_logic;
signal \N__3360\ : std_logic;
signal \N__3357\ : std_logic;
signal \N__3356\ : std_logic;
signal \N__3353\ : std_logic;
signal \N__3352\ : std_logic;
signal \N__3349\ : std_logic;
signal \N__3346\ : std_logic;
signal \N__3343\ : std_logic;
signal \N__3338\ : std_logic;
signal \N__3335\ : std_logic;
signal \N__3334\ : std_logic;
signal \N__3331\ : std_logic;
signal \N__3328\ : std_logic;
signal \N__3317\ : std_logic;
signal \N__3314\ : std_logic;
signal \N__3305\ : std_logic;
signal \N__3302\ : std_logic;
signal \N__3299\ : std_logic;
signal \N__3296\ : std_logic;
signal \N__3293\ : std_logic;
signal \N__3290\ : std_logic;
signal \N__3287\ : std_logic;
signal \N__3284\ : std_logic;
signal \N__3283\ : std_logic;
signal \N__3280\ : std_logic;
signal \N__3277\ : std_logic;
signal \N__3272\ : std_logic;
signal \N__3269\ : std_logic;
signal \N__3266\ : std_logic;
signal \N__3263\ : std_logic;
signal \N__3260\ : std_logic;
signal \N__3259\ : std_logic;
signal \N__3256\ : std_logic;
signal \N__3253\ : std_logic;
signal \N__3250\ : std_logic;
signal \N__3247\ : std_logic;
signal \N__3242\ : std_logic;
signal \N__3239\ : std_logic;
signal \N__3238\ : std_logic;
signal \N__3237\ : std_logic;
signal \N__3234\ : std_logic;
signal \N__3231\ : std_logic;
signal \N__3228\ : std_logic;
signal \N__3221\ : std_logic;
signal \N__3218\ : std_logic;
signal \N__3217\ : std_logic;
signal \N__3214\ : std_logic;
signal \N__3211\ : std_logic;
signal \N__3206\ : std_logic;
signal \N__3205\ : std_logic;
signal \N__3202\ : std_logic;
signal \N__3199\ : std_logic;
signal \N__3194\ : std_logic;
signal \N__3191\ : std_logic;
signal \N__3188\ : std_logic;
signal \N__3185\ : std_logic;
signal \N__3184\ : std_logic;
signal \N__3181\ : std_logic;
signal \N__3178\ : std_logic;
signal \N__3173\ : std_logic;
signal \N__3172\ : std_logic;
signal \N__3171\ : std_logic;
signal \N__3170\ : std_logic;
signal \N__3167\ : std_logic;
signal \N__3164\ : std_logic;
signal \N__3161\ : std_logic;
signal \N__3158\ : std_logic;
signal \N__3155\ : std_logic;
signal \N__3152\ : std_logic;
signal \N__3143\ : std_logic;
signal \N__3140\ : std_logic;
signal \N__3137\ : std_logic;
signal \N__3134\ : std_logic;
signal \N__3133\ : std_logic;
signal \N__3132\ : std_logic;
signal \N__3131\ : std_logic;
signal \N__3130\ : std_logic;
signal \N__3119\ : std_logic;
signal \N__3116\ : std_logic;
signal \N__3113\ : std_logic;
signal \N__3110\ : std_logic;
signal \N__3109\ : std_logic;
signal \N__3106\ : std_logic;
signal \N__3103\ : std_logic;
signal \N__3098\ : std_logic;
signal \N__3097\ : std_logic;
signal \N__3094\ : std_logic;
signal \N__3091\ : std_logic;
signal \N__3088\ : std_logic;
signal \N__3085\ : std_logic;
signal \N__3080\ : std_logic;
signal \N__3079\ : std_logic;
signal \N__3076\ : std_logic;
signal \N__3073\ : std_logic;
signal \N__3070\ : std_logic;
signal \N__3065\ : std_logic;
signal \N__3062\ : std_logic;
signal \N__3061\ : std_logic;
signal \N__3058\ : std_logic;
signal \N__3055\ : std_logic;
signal \N__3050\ : std_logic;
signal \N__3047\ : std_logic;
signal \N__3046\ : std_logic;
signal \N__3043\ : std_logic;
signal \N__3040\ : std_logic;
signal \N__3035\ : std_logic;
signal \N__3034\ : std_logic;
signal \N__3031\ : std_logic;
signal \N__3028\ : std_logic;
signal \N__3023\ : std_logic;
signal \N__3020\ : std_logic;
signal \N__3019\ : std_logic;
signal \N__3016\ : std_logic;
signal \N__3013\ : std_logic;
signal \N__3010\ : std_logic;
signal \N__3005\ : std_logic;
signal \N__3002\ : std_logic;
signal \N__3001\ : std_logic;
signal \N__2998\ : std_logic;
signal \N__2995\ : std_logic;
signal \N__2990\ : std_logic;
signal \N__2989\ : std_logic;
signal \N__2986\ : std_logic;
signal \N__2983\ : std_logic;
signal \N__2978\ : std_logic;
signal \N__2975\ : std_logic;
signal \N__2974\ : std_logic;
signal \N__2971\ : std_logic;
signal \N__2968\ : std_logic;
signal \N__2965\ : std_logic;
signal \N__2960\ : std_logic;
signal \N__2959\ : std_logic;
signal \N__2956\ : std_logic;
signal \N__2953\ : std_logic;
signal \N__2948\ : std_logic;
signal \N__2947\ : std_logic;
signal \N__2944\ : std_logic;
signal \N__2941\ : std_logic;
signal \N__2936\ : std_logic;
signal \N__2935\ : std_logic;
signal \N__2932\ : std_logic;
signal \N__2929\ : std_logic;
signal \N__2926\ : std_logic;
signal \N__2921\ : std_logic;
signal \N__2920\ : std_logic;
signal \N__2917\ : std_logic;
signal \N__2914\ : std_logic;
signal \N__2909\ : std_logic;
signal \N__2906\ : std_logic;
signal \N__2903\ : std_logic;
signal \N__2900\ : std_logic;
signal \N__2897\ : std_logic;
signal \N__2894\ : std_logic;
signal \N__2893\ : std_logic;
signal \N__2892\ : std_logic;
signal \N__2889\ : std_logic;
signal \N__2886\ : std_logic;
signal \N__2883\ : std_logic;
signal \N__2876\ : std_logic;
signal \N__2875\ : std_logic;
signal \N__2872\ : std_logic;
signal \N__2869\ : std_logic;
signal \N__2868\ : std_logic;
signal \N__2867\ : std_logic;
signal \N__2866\ : std_logic;
signal \N__2855\ : std_logic;
signal \N__2852\ : std_logic;
signal \N__2849\ : std_logic;
signal \N__2846\ : std_logic;
signal \N__2843\ : std_logic;
signal \N__2842\ : std_logic;
signal \N__2841\ : std_logic;
signal \N__2840\ : std_logic;
signal \N__2831\ : std_logic;
signal \N__2828\ : std_logic;
signal \N__2825\ : std_logic;
signal \N__2822\ : std_logic;
signal \N__2819\ : std_logic;
signal \N__2818\ : std_logic;
signal \N__2815\ : std_logic;
signal \N__2812\ : std_logic;
signal \N__2807\ : std_logic;
signal \N__2806\ : std_logic;
signal \N__2803\ : std_logic;
signal \N__2800\ : std_logic;
signal \N__2795\ : std_logic;
signal \N__2794\ : std_logic;
signal \N__2791\ : std_logic;
signal \N__2788\ : std_logic;
signal \N__2783\ : std_logic;
signal \N__2782\ : std_logic;
signal \N__2781\ : std_logic;
signal \N__2778\ : std_logic;
signal \N__2777\ : std_logic;
signal \N__2776\ : std_logic;
signal \N__2775\ : std_logic;
signal \N__2774\ : std_logic;
signal \N__2771\ : std_logic;
signal \N__2764\ : std_logic;
signal \N__2757\ : std_logic;
signal \N__2750\ : std_logic;
signal \N__2747\ : std_logic;
signal \N__2744\ : std_logic;
signal \N__2741\ : std_logic;
signal \N__2738\ : std_logic;
signal \N__2735\ : std_logic;
signal \N__2732\ : std_logic;
signal \N__2729\ : std_logic;
signal \N__2726\ : std_logic;
signal \N__2723\ : std_logic;
signal \N__2722\ : std_logic;
signal \N__2721\ : std_logic;
signal \N__2714\ : std_logic;
signal \N__2711\ : std_logic;
signal \N__2710\ : std_logic;
signal \N__2709\ : std_logic;
signal \N__2708\ : std_logic;
signal \N__2707\ : std_logic;
signal \N__2706\ : std_logic;
signal \N__2705\ : std_logic;
signal \N__2704\ : std_logic;
signal \N__2701\ : std_logic;
signal \N__2698\ : std_logic;
signal \N__2697\ : std_logic;
signal \N__2696\ : std_logic;
signal \N__2693\ : std_logic;
signal \N__2682\ : std_logic;
signal \N__2677\ : std_logic;
signal \N__2672\ : std_logic;
signal \N__2663\ : std_logic;
signal \N__2662\ : std_logic;
signal \N__2661\ : std_logic;
signal \N__2658\ : std_logic;
signal \N__2657\ : std_logic;
signal \N__2656\ : std_logic;
signal \N__2653\ : std_logic;
signal \N__2652\ : std_logic;
signal \N__2651\ : std_logic;
signal \N__2650\ : std_logic;
signal \N__2649\ : std_logic;
signal \N__2648\ : std_logic;
signal \N__2645\ : std_logic;
signal \N__2644\ : std_logic;
signal \N__2633\ : std_logic;
signal \N__2628\ : std_logic;
signal \N__2623\ : std_logic;
signal \N__2618\ : std_logic;
signal \N__2609\ : std_logic;
signal \N__2608\ : std_logic;
signal \N__2607\ : std_logic;
signal \N__2606\ : std_logic;
signal \N__2605\ : std_logic;
signal \N__2604\ : std_logic;
signal \N__2603\ : std_logic;
signal \N__2602\ : std_logic;
signal \N__2601\ : std_logic;
signal \N__2600\ : std_logic;
signal \N__2599\ : std_logic;
signal \N__2598\ : std_logic;
signal \N__2587\ : std_logic;
signal \N__2582\ : std_logic;
signal \N__2575\ : std_logic;
signal \N__2570\ : std_logic;
signal \N__2561\ : std_logic;
signal \N__2558\ : std_logic;
signal \N__2555\ : std_logic;
signal \N__2552\ : std_logic;
signal \N__2549\ : std_logic;
signal \N__2546\ : std_logic;
signal \N__2543\ : std_logic;
signal \N__2542\ : std_logic;
signal \N__2539\ : std_logic;
signal \N__2536\ : std_logic;
signal \N__2533\ : std_logic;
signal \N__2528\ : std_logic;
signal \N__2525\ : std_logic;
signal \N__2522\ : std_logic;
signal \N__2519\ : std_logic;
signal \N__2516\ : std_logic;
signal \N__2513\ : std_logic;
signal \N__2510\ : std_logic;
signal \N__2507\ : std_logic;
signal \N__2504\ : std_logic;
signal \N__2501\ : std_logic;
signal \N__2500\ : std_logic;
signal \N__2497\ : std_logic;
signal \N__2494\ : std_logic;
signal \N__2489\ : std_logic;
signal \N__2486\ : std_logic;
signal \N__2483\ : std_logic;
signal \N__2482\ : std_logic;
signal \N__2479\ : std_logic;
signal \N__2476\ : std_logic;
signal \N__2471\ : std_logic;
signal \N__2468\ : std_logic;
signal \N__2465\ : std_logic;
signal \N__2462\ : std_logic;
signal \N__2459\ : std_logic;
signal \N__2458\ : std_logic;
signal \N__2455\ : std_logic;
signal \N__2452\ : std_logic;
signal \N__2447\ : std_logic;
signal \N__2444\ : std_logic;
signal \N__2441\ : std_logic;
signal \N__2438\ : std_logic;
signal \N__2435\ : std_logic;
signal \N__2432\ : std_logic;
signal \N__2429\ : std_logic;
signal \N__2426\ : std_logic;
signal \N__2423\ : std_logic;
signal \N__2420\ : std_logic;
signal \N__2417\ : std_logic;
signal \N__2416\ : std_logic;
signal \N__2413\ : std_logic;
signal \N__2410\ : std_logic;
signal \N__2405\ : std_logic;
signal \N__2402\ : std_logic;
signal \N__2399\ : std_logic;
signal \N__2396\ : std_logic;
signal \N__2393\ : std_logic;
signal \N__2390\ : std_logic;
signal \N__2387\ : std_logic;
signal \N__2384\ : std_logic;
signal \N__2383\ : std_logic;
signal \N__2380\ : std_logic;
signal \N__2377\ : std_logic;
signal \N__2374\ : std_logic;
signal \N__2371\ : std_logic;
signal \N__2366\ : std_logic;
signal \N__2365\ : std_logic;
signal \N__2362\ : std_logic;
signal \N__2359\ : std_logic;
signal \N__2356\ : std_logic;
signal \N__2353\ : std_logic;
signal \N__2350\ : std_logic;
signal \N__2347\ : std_logic;
signal \N__2342\ : std_logic;
signal \N__2339\ : std_logic;
signal \N__2336\ : std_logic;
signal \N__2333\ : std_logic;
signal \N__2330\ : std_logic;
signal \N__2327\ : std_logic;
signal \N__2324\ : std_logic;
signal \N__2321\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal frame_decoder_dv_c : std_logic;
signal uart_input_c : std_logic;
signal \uart_sync.aux_0__0_Z0Z_0\ : std_logic;
signal \uart_sync.aux_1__0_Z0Z_0\ : std_logic;
signal \uart_sync.aux_2__0_Z0Z_0\ : std_logic;
signal \uart_sync.aux_3__0_Z0Z_0\ : std_logic;
signal \uart.N_133_0_cascade_\ : std_logic;
signal \uart.N_133_0\ : std_logic;
signal \uart.data_Auxce_0_6_cascade_\ : std_logic;
signal \uart.CO1_0\ : std_logic;
signal \bfn_8_1_0_\ : std_logic;
signal \reset_module_System.count_1_cry_1\ : std_logic;
signal \reset_module_System.count_1_cry_2\ : std_logic;
signal \reset_module_System.count_1_cry_3\ : std_logic;
signal \reset_module_System.count_1_cry_4\ : std_logic;
signal \reset_module_System.count_1_cry_5\ : std_logic;
signal \reset_module_System.count_1_cry_6\ : std_logic;
signal \reset_module_System.count_1_cry_7\ : std_logic;
signal \reset_module_System.count_1_cry_8\ : std_logic;
signal \bfn_8_2_0_\ : std_logic;
signal \reset_module_System.count_1_cry_9\ : std_logic;
signal \reset_module_System.count_1_cry_10\ : std_logic;
signal \reset_module_System.count_1_cry_11\ : std_logic;
signal \reset_module_System.countZ0Z_13\ : std_logic;
signal \reset_module_System.count_1_cry_12\ : std_logic;
signal \reset_module_System.count_1_cry_13\ : std_logic;
signal \reset_module_System.countZ0Z_15\ : std_logic;
signal \reset_module_System.count_1_cry_14\ : std_logic;
signal \reset_module_System.count_1_cry_15\ : std_logic;
signal \reset_module_System.count_1_cry_16\ : std_logic;
signal \bfn_8_3_0_\ : std_logic;
signal \reset_module_System.count_1_cry_17\ : std_logic;
signal \reset_module_System.countZ0Z_19\ : std_logic;
signal \reset_module_System.count_1_cry_18\ : std_logic;
signal \reset_module_System.count_1_cry_19\ : std_logic;
signal \reset_module_System.count_1_cry_20\ : std_logic;
signal \reset_module_System.countZ0Z_21\ : std_logic;
signal \uart.data_Auxce_0_5\ : std_logic;
signal \uart.timer_Count_RNI9M0NZ0Z_1\ : std_logic;
signal \uart.timer_Count_RNILKMA1Z0Z_0_cascade_\ : std_logic;
signal \uart.un1_state_2_0_cascade_\ : std_logic;
signal \uart.un1_state_2_0\ : std_logic;
signal \uart.data_Auxce_0_0_4\ : std_logic;
signal \uart.data_Auxce_0_0_0\ : std_logic;
signal \uart.data_Auxce_0_1\ : std_logic;
signal \uart.data_Auxce_0_0_2\ : std_logic;
signal \uart.un1_state_5_0\ : std_logic;
signal \uart.bit_CountZ0Z_2\ : std_logic;
signal \uart.bit_CountZ0Z_1\ : std_logic;
signal \uart.bit_CountZ0Z_0\ : std_logic;
signal \uart.data_Auxce_0_3\ : std_logic;
signal \reset_module_System.countZ0Z_16\ : std_logic;
signal \reset_module_System.countZ0Z_4\ : std_logic;
signal \reset_module_System.countZ0Z_18\ : std_logic;
signal \reset_module_System.reset6_14_cascade_\ : std_logic;
signal \reset_module_System.countZ0Z_6\ : std_logic;
signal \reset_module_System.countZ0Z_3\ : std_logic;
signal \reset_module_System.countZ0Z_20\ : std_logic;
signal \reset_module_System.countZ0Z_8\ : std_logic;
signal \reset_module_System.countZ0Z_7\ : std_logic;
signal \reset_module_System.countZ0Z_9\ : std_logic;
signal \reset_module_System.countZ0Z_5\ : std_logic;
signal \reset_module_System.count_1_1\ : std_logic;
signal \reset_module_System.countZ0Z_1\ : std_logic;
signal \reset_module_System.reset6_15\ : std_logic;
signal \reset_module_System.reset6_14\ : std_logic;
signal \reset_module_System.count_1_2\ : std_logic;
signal \reset_module_System.countZ0Z_2\ : std_logic;
signal \reset_module_System.countZ0Z_11\ : std_logic;
signal \reset_module_System.countZ0Z_10\ : std_logic;
signal \reset_module_System.countZ0Z_14\ : std_logic;
signal \reset_module_System.countZ0Z_17\ : std_logic;
signal \reset_module_System.reset6_3_cascade_\ : std_logic;
signal \reset_module_System.reset6_13\ : std_logic;
signal \reset_module_System.countZ0Z_12\ : std_logic;
signal \reset_module_System.countZ0Z_0\ : std_logic;
signal \reset_module_System.reset6_17_cascade_\ : std_logic;
signal \reset_module_System.reset6_11\ : std_logic;
signal \reset_module_System.reset6_19\ : std_logic;
signal \uart.N_169_cascade_\ : std_logic;
signal \uart.state_srsts_i_1_3_cascade_\ : std_logic;
signal \uart.data_AuxZ0Z_0\ : std_logic;
signal \uart.data_AuxZ0Z_2\ : std_logic;
signal \uart.data_AuxZ0Z_3\ : std_logic;
signal \uart.data_AuxZ0Z_5\ : std_logic;
signal \uart.data_AuxZ0Z_7\ : std_logic;
signal \uart.timer_Count10lto5_0_0_cascade_\ : std_logic;
signal \uart.N_177\ : std_logic;
signal \uart.N_168_cascade_\ : std_logic;
signal \uart.state_RNIAFHLZ0Z_4\ : std_logic;
signal \uart.stateZ0Z_1\ : std_logic;
signal \uart.N_151_cascade_\ : std_logic;
signal \uart.stateZ0Z_2\ : std_logic;
signal \uart.stateZ0Z_3\ : std_logic;
signal \uart.state_srsts_i_1_1_3\ : std_logic;
signal \uart.N_166_cascade_\ : std_logic;
signal \uart.state_srsts_0_1_0_cascade_\ : std_logic;
signal \uart.stateZ0Z_0\ : std_logic;
signal \uart_frame_decoder.N_43\ : std_logic;
signal \uart_frame_decoder.N_43_cascade_\ : std_logic;
signal \uart_frame_decoder.state_1_ns_i_i_a2_1_1_0_cascade_\ : std_logic;
signal \uart_frame_decoder.N_81_cascade_\ : std_logic;
signal \uart_frame_decoder.state_1_ns_0_i_a2_0_0_1Z0Z_2_cascade_\ : std_logic;
signal uart_data_3 : std_logic;
signal \uart_frame_decoder.state_1_ns_0_i_a2_1_0Z0Z_2_cascade_\ : std_logic;
signal uart_data_2 : std_logic;
signal uart_data_5 : std_logic;
signal uart_data_7 : std_logic;
signal uart_data_0 : std_logic;
signal \uart_frame_decoder.N_79_4\ : std_logic;
signal \uart_frame_decoder.N_79_4_cascade_\ : std_logic;
signal uart_input_sync : std_logic;
signal \uart.data_8_0_cascade_\ : std_logic;
signal \uart.state_srsts_0_a3_1_4\ : std_logic;
signal \uart.N_152_0_cascade_\ : std_logic;
signal \uart.N_167\ : std_logic;
signal \uart.N_159\ : std_logic;
signal \uart.N_167_cascade_\ : std_logic;
signal \uart.N_180\ : std_logic;
signal \uart.N_152_0\ : std_logic;
signal \uart.stateZ0Z_4\ : std_logic;
signal \uart.N_145_0\ : std_logic;
signal \uart.state_1_sqmuxa\ : std_logic;
signal \uart.state_1_sqmuxa_cascade_\ : std_logic;
signal \bfn_10_5_0_\ : std_logic;
signal \uart.timer_CountZ0Z_2\ : std_logic;
signal \uart.un4_timer_Count_1_cry_1\ : std_logic;
signal \uart.timer_CountZ0Z_3\ : std_logic;
signal \uart.un4_timer_Count_1_cry_2\ : std_logic;
signal \uart.timer_CountZ0Z_4\ : std_logic;
signal \uart.un4_timer_Count_1_cry_3\ : std_logic;
signal \uart.timer_CountZ0Z_5\ : std_logic;
signal \uart.un4_timer_Count_1_cry_4\ : std_logic;
signal \uart.timer_CountZ0Z_6\ : std_logic;
signal \uart.un4_timer_Count_1_cry_5\ : std_logic;
signal \uart.un4_timer_Count_1_cry_6\ : std_logic;
signal \uart.timer_CountZ0Z_7\ : std_logic;
signal \bfn_11_1_0_\ : std_logic;
signal \uart_frame_decoder.count8_axb_1\ : std_logic;
signal \uart_frame_decoder.count8_cry_0\ : std_logic;
signal \uart_frame_decoder.count_i_2\ : std_logic;
signal \uart_frame_decoder.count8_cry_1\ : std_logic;
signal \uart_frame_decoder.count8\ : std_logic;
signal \uart_frame_decoder.count8_THRU_CO\ : std_logic;
signal \uart_frame_decoder.count8_THRU_CO_cascade_\ : std_logic;
signal \uart_frame_decoder.N_37\ : std_logic;
signal \uart_frame_decoder.N_37_cascade_\ : std_logic;
signal \uart_frame_decoder.countZ0Z_1\ : std_logic;
signal \uart_frame_decoder.countZ0Z_2\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \uart_frame_decoder.count8_0\ : std_logic;
signal \uart_frame_decoder.count8_0_i\ : std_logic;
signal \uart_frame_decoder.N_4_0_cascade_\ : std_logic;
signal \uart_frame_decoder.g0_1_0_1\ : std_logic;
signal \uart_frame_decoder.g0_1_a3_3\ : std_logic;
signal \uart_frame_decoder.WDT8lto15_cascade_\ : std_logic;
signal \uart_frame_decoder.state_1_ns_0_i_o2_0_tz_10\ : std_logic;
signal \uart_frame_decoder.state_1_ns_i_i_a2_1_1_0\ : std_logic;
signal \uart_frame_decoder.state_1Z0Z_0\ : std_logic;
signal \uart_frame_decoder.state_1_ns_0_i_a2_0_0_0_10_cascade_\ : std_logic;
signal \uart_frame_decoder.N_35_i_1\ : std_logic;
signal \uart.timer_CountZ0Z_1\ : std_logic;
signal \uart_frame_decoder.WDT_RNIQAB11Z0Z_4\ : std_logic;
signal \uart_frame_decoder.WDT_RNISS5HZ0Z_11_cascade_\ : std_logic;
signal \uart_frame_decoder.WDT8lt13_cascade_\ : std_logic;
signal \uart_frame_decoder.state_1_ns_i_i_a2_0_0\ : std_logic;
signal \uart_frame_decoder.WDT8lt13\ : std_logic;
signal \uart_frame_decoder.WDT8lto15\ : std_logic;
signal \uart_frame_decoder.N_80\ : std_logic;
signal \uart.timer_CountZ0Z_0\ : std_logic;
signal \uart.timer_Count_1_sqmuxa_i\ : std_logic;
signal \uart_frame_decoder.state_1_ns_0_i_a2_0_0_1\ : std_logic;
signal \uart_frame_decoder.N_99\ : std_logic;
signal \uart_frame_decoder.N_92\ : std_logic;
signal \uart.data_AuxZ0Z_1\ : std_logic;
signal uart_data_1 : std_logic;
signal \uart.data_AuxZ0Z_4\ : std_logic;
signal uart_data_4 : std_logic;
signal \uart.data_AuxZ0Z_6\ : std_logic;
signal uart_data_6 : std_logic;
signal \uart.state_1_sqmuxa_0\ : std_logic;
signal \uart.timer_Count_RNIS4183Z0Z_7\ : std_logic;
signal \uart_frame_decoder.WDT8_0_i\ : std_logic;
signal \uart_frame_decoder.WDTZ0Z_0\ : std_logic;
signal \bfn_12_2_0_\ : std_logic;
signal \uart_frame_decoder.WDTZ0Z_1\ : std_logic;
signal \uart_frame_decoder.un1_WDT_cry_0\ : std_logic;
signal \uart_frame_decoder.WDTZ0Z_2\ : std_logic;
signal \uart_frame_decoder.un1_WDT_cry_1\ : std_logic;
signal \uart_frame_decoder.WDTZ0Z_3\ : std_logic;
signal \uart_frame_decoder.un1_WDT_cry_2\ : std_logic;
signal \uart_frame_decoder.WDTZ0Z_4\ : std_logic;
signal \uart_frame_decoder.un1_WDT_cry_3\ : std_logic;
signal \uart_frame_decoder.WDTZ0Z_5\ : std_logic;
signal \uart_frame_decoder.un1_WDT_cry_4\ : std_logic;
signal \uart_frame_decoder.WDTZ0Z_6\ : std_logic;
signal \uart_frame_decoder.un1_WDT_cry_5\ : std_logic;
signal \uart_frame_decoder.WDTZ0Z_7\ : std_logic;
signal \uart_frame_decoder.un1_WDT_cry_6\ : std_logic;
signal \uart_frame_decoder.un1_WDT_cry_7\ : std_logic;
signal \uart_frame_decoder.WDTZ0Z_8\ : std_logic;
signal \bfn_12_3_0_\ : std_logic;
signal \uart_frame_decoder.WDTZ0Z_9\ : std_logic;
signal \uart_frame_decoder.un1_WDT_cry_8\ : std_logic;
signal \uart_frame_decoder.WDTZ0Z_10\ : std_logic;
signal \uart_frame_decoder.un1_WDT_cry_9\ : std_logic;
signal \uart_frame_decoder.WDTZ0Z_11\ : std_logic;
signal \uart_frame_decoder.un1_WDT_cry_10\ : std_logic;
signal \uart_frame_decoder.WDTZ0Z_12\ : std_logic;
signal \uart_frame_decoder.un1_WDT_cry_11\ : std_logic;
signal \uart_frame_decoder.WDTZ0Z_13\ : std_logic;
signal \uart_frame_decoder.un1_WDT_cry_12\ : std_logic;
signal \uart_frame_decoder.WDTZ0Z_14\ : std_logic;
signal \uart_frame_decoder.un1_WDT_cry_13\ : std_logic;
signal \uart_frame_decoder.un1_WDT_cry_14\ : std_logic;
signal \uart_frame_decoder.WDTZ0Z_15\ : std_logic;
signal \uart_frame_decoder.state_1_ns_0_i_a2_0_0_0_10\ : std_logic;
signal \uart_frame_decoder.state_1_ns_0_i_a2_0_d_10\ : std_logic;
signal \uart_frame_decoder.N_85\ : std_logic;
signal clk_system_c_g : std_logic;
signal \reset_module_System_reset_iso\ : std_logic;
signal uart_data_rdy_c : std_logic;
signal reset_system : std_logic;
signal \uart_frame_decoder.source_data_valid_2_sqmuxa_iZ0\ : std_logic;
signal \uart_frame_decoder.state_1Z0Z_4\ : std_logic;
signal \uart_frame_decoder_N_307_i\ : std_logic;
signal \uart_frame_decoder.state_1Z0Z_8\ : std_logic;
signal \uart_frame_decoder_N_308_i\ : std_logic;
signal \uart_frame_decoder.state_1Z0Z_1\ : std_logic;
signal \uart_frame_decoder.state_1Z0Z_9\ : std_logic;
signal \uart_frame_decoder.un14_i_a2_0_a2_1_0_cascade_\ : std_logic;
signal \uart_frame_decoder.state_1Z0Z_5\ : std_logic;
signal \uart_frame_decoder_N_305_i\ : std_logic;
signal \uart_frame_decoder.state_1Z0Z_6\ : std_logic;
signal \uart_frame_decoder.state_1Z0Z_7\ : std_logic;
signal \uart_frame_decoder.N_306_1\ : std_logic;
signal \uart_frame_decoder.state_1Z0Z_2\ : std_logic;
signal \uart_frame_decoder.state_1Z0Z_3\ : std_logic;
signal \uart_frame_decoder.N_306_1_cascade_\ : std_logic;
signal \uart_frame_decoder.state_1Z0Z_10\ : std_logic;
signal \uart_frame_decoder_N_306_i\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal clk_system_wire : std_logic;
signal debug_state_output_wire : std_logic_vector(4 downto 0);
signal uart_data_rdy_wire : std_logic;
signal debug_sinkdatavalid_output_wire : std_logic;
signal frame_decoder_dv_wire : std_logic;
signal uart_input_wire : std_logic;
signal uart_input_debug_wire : std_logic;

begin
    clk_system_wire <= clk_system;
    debug_state_output <= debug_state_output_wire;
    uart_data_rdy <= uart_data_rdy_wire;
    debug_sinkdatavalid_output <= debug_sinkdatavalid_output_wire;
    frame_decoder_dv <= frame_decoder_dv_wire;
    uart_input_wire <= uart_input;
    uart_input_debug <= uart_input_debug_wire;

    \clk_system_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__5661\,
            GLOBALBUFFEROUTPUT => clk_system_c_g
        );

    \clk_system_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5663\,
            DIN => \N__5662\,
            DOUT => \N__5661\,
            PACKAGEPIN => clk_system_wire
        );

    \clk_system_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5663\,
            PADOUT => \N__5662\,
            PADIN => \N__5661\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \debug_state_output_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5652\,
            DIN => \N__5651\,
            DOUT => \N__5650\,
            PACKAGEPIN => debug_state_output_wire(4)
        );

    \debug_state_output_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5652\,
            PADOUT => \N__5651\,
            PADIN => \N__5650\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \debug_state_output_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5643\,
            DIN => \N__5642\,
            DOUT => \N__5641\,
            PACKAGEPIN => debug_state_output_wire(1)
        );

    \debug_state_output_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5643\,
            PADOUT => \N__5642\,
            PADIN => \N__5641\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4970\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \uart_data_rdy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5634\,
            DIN => \N__5633\,
            DOUT => \N__5632\,
            PACKAGEPIN => uart_data_rdy_wire
        );

    \uart_data_rdy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5634\,
            PADOUT => \N__5633\,
            PADIN => \N__5632\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5503\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \debug_state_output_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5625\,
            DIN => \N__5624\,
            DOUT => \N__5623\,
            PACKAGEPIN => debug_state_output_wire(3)
        );

    \debug_state_output_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5625\,
            PADOUT => \N__5624\,
            PADIN => \N__5623\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5228\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \debug_sinkdatavalid_output_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5616\,
            DIN => \N__5615\,
            DOUT => \N__5614\,
            PACKAGEPIN => debug_sinkdatavalid_output_wire
        );

    \debug_sinkdatavalid_output_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5616\,
            PADOUT => \N__5615\,
            PADIN => \N__5614\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5502\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \frame_decoder_dv_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5607\,
            DIN => \N__5606\,
            DOUT => \N__5605\,
            PACKAGEPIN => frame_decoder_dv_wire
        );

    \frame_decoder_dv_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5607\,
            PADOUT => \N__5606\,
            PADIN => \N__5605\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2393\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \uart_input_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5598\,
            DIN => \N__5597\,
            DOUT => \N__5596\,
            PACKAGEPIN => uart_input_wire
        );

    \uart_input_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5598\,
            PADOUT => \N__5597\,
            PADIN => \N__5596\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => uart_input_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \debug_state_output_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5589\,
            DIN => \N__5588\,
            DOUT => \N__5587\,
            PACKAGEPIN => debug_state_output_wire(0)
        );

    \debug_state_output_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5589\,
            PADOUT => \N__5588\,
            PADIN => \N__5587\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5138\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \debug_state_output_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5580\,
            DIN => \N__5579\,
            DOUT => \N__5578\,
            PACKAGEPIN => debug_state_output_wire(2)
        );

    \debug_state_output_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5580\,
            PADOUT => \N__5579\,
            PADIN => \N__5578\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5261\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \uart_input_debug_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5571\,
            DIN => \N__5570\,
            DOUT => \N__5569\,
            PACKAGEPIN => uart_input_debug_wire
        );

    \uart_input_debug_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5571\,
            PADOUT => \N__5570\,
            PADIN => \N__5569\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2365\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__1274\ : SRMux
    port map (
            O => \N__5552\,
            I => \N__5546\
        );

    \I__1273\ : SRMux
    port map (
            O => \N__5551\,
            I => \N__5543\
        );

    \I__1272\ : SRMux
    port map (
            O => \N__5550\,
            I => \N__5540\
        );

    \I__1271\ : SRMux
    port map (
            O => \N__5549\,
            I => \N__5537\
        );

    \I__1270\ : LocalMux
    port map (
            O => \N__5546\,
            I => \N__5533\
        );

    \I__1269\ : LocalMux
    port map (
            O => \N__5543\,
            I => \N__5530\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__5540\,
            I => \N__5527\
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__5537\,
            I => \N__5524\
        );

    \I__1266\ : SRMux
    port map (
            O => \N__5536\,
            I => \N__5521\
        );

    \I__1265\ : Span4Mux_v
    port map (
            O => \N__5533\,
            I => \N__5518\
        );

    \I__1264\ : Span4Mux_s0_v
    port map (
            O => \N__5530\,
            I => \N__5511\
        );

    \I__1263\ : Span4Mux_v
    port map (
            O => \N__5527\,
            I => \N__5511\
        );

    \I__1262\ : Span4Mux_v
    port map (
            O => \N__5524\,
            I => \N__5511\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__5521\,
            I => \reset_module_System_reset_iso\
        );

    \I__1260\ : Odrv4
    port map (
            O => \N__5518\,
            I => \reset_module_System_reset_iso\
        );

    \I__1259\ : Odrv4
    port map (
            O => \N__5511\,
            I => \reset_module_System_reset_iso\
        );

    \I__1258\ : CascadeMux
    port map (
            O => \N__5504\,
            I => \N__5498\
        );

    \I__1257\ : IoInMux
    port map (
            O => \N__5503\,
            I => \N__5488\
        );

    \I__1256\ : IoInMux
    port map (
            O => \N__5502\,
            I => \N__5485\
        );

    \I__1255\ : InMux
    port map (
            O => \N__5501\,
            I => \N__5482\
        );

    \I__1254\ : InMux
    port map (
            O => \N__5498\,
            I => \N__5479\
        );

    \I__1253\ : InMux
    port map (
            O => \N__5497\,
            I => \N__5464\
        );

    \I__1252\ : InMux
    port map (
            O => \N__5496\,
            I => \N__5464\
        );

    \I__1251\ : InMux
    port map (
            O => \N__5495\,
            I => \N__5464\
        );

    \I__1250\ : InMux
    port map (
            O => \N__5494\,
            I => \N__5464\
        );

    \I__1249\ : InMux
    port map (
            O => \N__5493\,
            I => \N__5464\
        );

    \I__1248\ : InMux
    port map (
            O => \N__5492\,
            I => \N__5464\
        );

    \I__1247\ : InMux
    port map (
            O => \N__5491\,
            I => \N__5464\
        );

    \I__1246\ : LocalMux
    port map (
            O => \N__5488\,
            I => \N__5461\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__5485\,
            I => \N__5450\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__5482\,
            I => \N__5450\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__5479\,
            I => \N__5445\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__5464\,
            I => \N__5445\
        );

    \I__1241\ : Span4Mux_s2_v
    port map (
            O => \N__5461\,
            I => \N__5440\
        );

    \I__1240\ : InMux
    port map (
            O => \N__5460\,
            I => \N__5437\
        );

    \I__1239\ : InMux
    port map (
            O => \N__5459\,
            I => \N__5432\
        );

    \I__1238\ : InMux
    port map (
            O => \N__5458\,
            I => \N__5432\
        );

    \I__1237\ : InMux
    port map (
            O => \N__5457\,
            I => \N__5427\
        );

    \I__1236\ : InMux
    port map (
            O => \N__5456\,
            I => \N__5427\
        );

    \I__1235\ : InMux
    port map (
            O => \N__5455\,
            I => \N__5424\
        );

    \I__1234\ : Span4Mux_s2_v
    port map (
            O => \N__5450\,
            I => \N__5419\
        );

    \I__1233\ : Span4Mux_h
    port map (
            O => \N__5445\,
            I => \N__5416\
        );

    \I__1232\ : InMux
    port map (
            O => \N__5444\,
            I => \N__5411\
        );

    \I__1231\ : InMux
    port map (
            O => \N__5443\,
            I => \N__5411\
        );

    \I__1230\ : Span4Mux_h
    port map (
            O => \N__5440\,
            I => \N__5406\
        );

    \I__1229\ : LocalMux
    port map (
            O => \N__5437\,
            I => \N__5406\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__5432\,
            I => \N__5401\
        );

    \I__1227\ : LocalMux
    port map (
            O => \N__5427\,
            I => \N__5401\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__5424\,
            I => \N__5398\
        );

    \I__1225\ : InMux
    port map (
            O => \N__5423\,
            I => \N__5393\
        );

    \I__1224\ : InMux
    port map (
            O => \N__5422\,
            I => \N__5393\
        );

    \I__1223\ : Odrv4
    port map (
            O => \N__5419\,
            I => uart_data_rdy_c
        );

    \I__1222\ : Odrv4
    port map (
            O => \N__5416\,
            I => uart_data_rdy_c
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__5411\,
            I => uart_data_rdy_c
        );

    \I__1220\ : Odrv4
    port map (
            O => \N__5406\,
            I => uart_data_rdy_c
        );

    \I__1219\ : Odrv4
    port map (
            O => \N__5401\,
            I => uart_data_rdy_c
        );

    \I__1218\ : Odrv4
    port map (
            O => \N__5398\,
            I => uart_data_rdy_c
        );

    \I__1217\ : LocalMux
    port map (
            O => \N__5393\,
            I => uart_data_rdy_c
        );

    \I__1216\ : InMux
    port map (
            O => \N__5378\,
            I => \N__5373\
        );

    \I__1215\ : InMux
    port map (
            O => \N__5377\,
            I => \N__5369\
        );

    \I__1214\ : InMux
    port map (
            O => \N__5376\,
            I => \N__5365\
        );

    \I__1213\ : LocalMux
    port map (
            O => \N__5373\,
            I => \N__5355\
        );

    \I__1212\ : InMux
    port map (
            O => \N__5372\,
            I => \N__5352\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__5369\,
            I => \N__5349\
        );

    \I__1210\ : InMux
    port map (
            O => \N__5368\,
            I => \N__5346\
        );

    \I__1209\ : LocalMux
    port map (
            O => \N__5365\,
            I => \N__5343\
        );

    \I__1208\ : InMux
    port map (
            O => \N__5364\,
            I => \N__5338\
        );

    \I__1207\ : InMux
    port map (
            O => \N__5363\,
            I => \N__5338\
        );

    \I__1206\ : InMux
    port map (
            O => \N__5362\,
            I => \N__5331\
        );

    \I__1205\ : InMux
    port map (
            O => \N__5361\,
            I => \N__5331\
        );

    \I__1204\ : InMux
    port map (
            O => \N__5360\,
            I => \N__5331\
        );

    \I__1203\ : InMux
    port map (
            O => \N__5359\,
            I => \N__5328\
        );

    \I__1202\ : InMux
    port map (
            O => \N__5358\,
            I => \N__5325\
        );

    \I__1201\ : Span4Mux_v
    port map (
            O => \N__5355\,
            I => \N__5318\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__5352\,
            I => \N__5318\
        );

    \I__1199\ : Span4Mux_v
    port map (
            O => \N__5349\,
            I => \N__5318\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__5346\,
            I => \N__5309\
        );

    \I__1197\ : Span4Mux_v
    port map (
            O => \N__5343\,
            I => \N__5309\
        );

    \I__1196\ : LocalMux
    port map (
            O => \N__5338\,
            I => \N__5309\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__5331\,
            I => \N__5309\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__5328\,
            I => reset_system
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__5325\,
            I => reset_system
        );

    \I__1192\ : Odrv4
    port map (
            O => \N__5318\,
            I => reset_system
        );

    \I__1191\ : Odrv4
    port map (
            O => \N__5309\,
            I => reset_system
        );

    \I__1190\ : SRMux
    port map (
            O => \N__5300\,
            I => \N__5297\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__5297\,
            I => \N__5293\
        );

    \I__1188\ : SRMux
    port map (
            O => \N__5296\,
            I => \N__5290\
        );

    \I__1187\ : Span4Mux_s2_v
    port map (
            O => \N__5293\,
            I => \N__5287\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__5290\,
            I => \N__5284\
        );

    \I__1185\ : Odrv4
    port map (
            O => \N__5287\,
            I => \uart_frame_decoder.source_data_valid_2_sqmuxa_iZ0\
        );

    \I__1184\ : Odrv4
    port map (
            O => \N__5284\,
            I => \uart_frame_decoder.source_data_valid_2_sqmuxa_iZ0\
        );

    \I__1183\ : CascadeMux
    port map (
            O => \N__5279\,
            I => \N__5275\
        );

    \I__1182\ : InMux
    port map (
            O => \N__5278\,
            I => \N__5271\
        );

    \I__1181\ : InMux
    port map (
            O => \N__5275\,
            I => \N__5266\
        );

    \I__1180\ : InMux
    port map (
            O => \N__5274\,
            I => \N__5266\
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__5271\,
            I => \uart_frame_decoder.state_1Z0Z_4\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__5266\,
            I => \uart_frame_decoder.state_1Z0Z_4\
        );

    \I__1177\ : IoInMux
    port map (
            O => \N__5261\,
            I => \N__5258\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__5258\,
            I => \N__5255\
        );

    \I__1175\ : IoSpan4Mux
    port map (
            O => \N__5255\,
            I => \N__5252\
        );

    \I__1174\ : IoSpan4Mux
    port map (
            O => \N__5252\,
            I => \N__5249\
        );

    \I__1173\ : Odrv4
    port map (
            O => \N__5249\,
            I => \uart_frame_decoder_N_307_i\
        );

    \I__1172\ : CascadeMux
    port map (
            O => \N__5246\,
            I => \N__5241\
        );

    \I__1171\ : InMux
    port map (
            O => \N__5245\,
            I => \N__5238\
        );

    \I__1170\ : InMux
    port map (
            O => \N__5244\,
            I => \N__5233\
        );

    \I__1169\ : InMux
    port map (
            O => \N__5241\,
            I => \N__5233\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__5238\,
            I => \uart_frame_decoder.state_1Z0Z_8\
        );

    \I__1167\ : LocalMux
    port map (
            O => \N__5233\,
            I => \uart_frame_decoder.state_1Z0Z_8\
        );

    \I__1166\ : IoInMux
    port map (
            O => \N__5228\,
            I => \N__5225\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__5225\,
            I => \N__5222\
        );

    \I__1164\ : Span4Mux_s3_v
    port map (
            O => \N__5222\,
            I => \N__5219\
        );

    \I__1163\ : Odrv4
    port map (
            O => \N__5219\,
            I => \uart_frame_decoder_N_308_i\
        );

    \I__1162\ : InMux
    port map (
            O => \N__5216\,
            I => \N__5212\
        );

    \I__1161\ : InMux
    port map (
            O => \N__5215\,
            I => \N__5208\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__5212\,
            I => \N__5203\
        );

    \I__1159\ : InMux
    port map (
            O => \N__5211\,
            I => \N__5200\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__5208\,
            I => \N__5197\
        );

    \I__1157\ : InMux
    port map (
            O => \N__5207\,
            I => \N__5192\
        );

    \I__1156\ : InMux
    port map (
            O => \N__5206\,
            I => \N__5192\
        );

    \I__1155\ : Odrv4
    port map (
            O => \N__5203\,
            I => \uart_frame_decoder.state_1Z0Z_1\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__5200\,
            I => \uart_frame_decoder.state_1Z0Z_1\
        );

    \I__1153\ : Odrv4
    port map (
            O => \N__5197\,
            I => \uart_frame_decoder.state_1Z0Z_1\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__5192\,
            I => \uart_frame_decoder.state_1Z0Z_1\
        );

    \I__1151\ : CascadeMux
    port map (
            O => \N__5183\,
            I => \N__5177\
        );

    \I__1150\ : InMux
    port map (
            O => \N__5182\,
            I => \N__5172\
        );

    \I__1149\ : InMux
    port map (
            O => \N__5181\,
            I => \N__5172\
        );

    \I__1148\ : InMux
    port map (
            O => \N__5180\,
            I => \N__5167\
        );

    \I__1147\ : InMux
    port map (
            O => \N__5177\,
            I => \N__5167\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__5172\,
            I => \uart_frame_decoder.state_1Z0Z_9\
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__5167\,
            I => \uart_frame_decoder.state_1Z0Z_9\
        );

    \I__1144\ : CascadeMux
    port map (
            O => \N__5162\,
            I => \uart_frame_decoder.un14_i_a2_0_a2_1_0_cascade_\
        );

    \I__1143\ : CascadeMux
    port map (
            O => \N__5159\,
            I => \N__5154\
        );

    \I__1142\ : InMux
    port map (
            O => \N__5158\,
            I => \N__5148\
        );

    \I__1141\ : InMux
    port map (
            O => \N__5157\,
            I => \N__5148\
        );

    \I__1140\ : InMux
    port map (
            O => \N__5154\,
            I => \N__5143\
        );

    \I__1139\ : InMux
    port map (
            O => \N__5153\,
            I => \N__5143\
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__5148\,
            I => \uart_frame_decoder.state_1Z0Z_5\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__5143\,
            I => \uart_frame_decoder.state_1Z0Z_5\
        );

    \I__1136\ : IoInMux
    port map (
            O => \N__5138\,
            I => \N__5135\
        );

    \I__1135\ : LocalMux
    port map (
            O => \N__5135\,
            I => \N__5132\
        );

    \I__1134\ : IoSpan4Mux
    port map (
            O => \N__5132\,
            I => \N__5129\
        );

    \I__1133\ : Span4Mux_s3_v
    port map (
            O => \N__5129\,
            I => \N__5126\
        );

    \I__1132\ : Odrv4
    port map (
            O => \N__5126\,
            I => \uart_frame_decoder_N_305_i\
        );

    \I__1131\ : CascadeMux
    port map (
            O => \N__5123\,
            I => \N__5119\
        );

    \I__1130\ : InMux
    port map (
            O => \N__5122\,
            I => \N__5115\
        );

    \I__1129\ : InMux
    port map (
            O => \N__5119\,
            I => \N__5110\
        );

    \I__1128\ : InMux
    port map (
            O => \N__5118\,
            I => \N__5110\
        );

    \I__1127\ : LocalMux
    port map (
            O => \N__5115\,
            I => \uart_frame_decoder.state_1Z0Z_6\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__5110\,
            I => \uart_frame_decoder.state_1Z0Z_6\
        );

    \I__1125\ : CascadeMux
    port map (
            O => \N__5105\,
            I => \N__5099\
        );

    \I__1124\ : InMux
    port map (
            O => \N__5104\,
            I => \N__5094\
        );

    \I__1123\ : InMux
    port map (
            O => \N__5103\,
            I => \N__5094\
        );

    \I__1122\ : InMux
    port map (
            O => \N__5102\,
            I => \N__5089\
        );

    \I__1121\ : InMux
    port map (
            O => \N__5099\,
            I => \N__5089\
        );

    \I__1120\ : LocalMux
    port map (
            O => \N__5094\,
            I => \uart_frame_decoder.state_1Z0Z_7\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__5089\,
            I => \uart_frame_decoder.state_1Z0Z_7\
        );

    \I__1118\ : InMux
    port map (
            O => \N__5084\,
            I => \N__5081\
        );

    \I__1117\ : LocalMux
    port map (
            O => \N__5081\,
            I => \uart_frame_decoder.N_306_1\
        );

    \I__1116\ : InMux
    port map (
            O => \N__5078\,
            I => \N__5075\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__5075\,
            I => \N__5070\
        );

    \I__1114\ : InMux
    port map (
            O => \N__5074\,
            I => \N__5067\
        );

    \I__1113\ : InMux
    port map (
            O => \N__5073\,
            I => \N__5064\
        );

    \I__1112\ : Odrv4
    port map (
            O => \N__5070\,
            I => \uart_frame_decoder.state_1Z0Z_2\
        );

    \I__1111\ : LocalMux
    port map (
            O => \N__5067\,
            I => \uart_frame_decoder.state_1Z0Z_2\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__5064\,
            I => \uart_frame_decoder.state_1Z0Z_2\
        );

    \I__1109\ : CascadeMux
    port map (
            O => \N__5057\,
            I => \N__5052\
        );

    \I__1108\ : InMux
    port map (
            O => \N__5056\,
            I => \N__5046\
        );

    \I__1107\ : InMux
    port map (
            O => \N__5055\,
            I => \N__5046\
        );

    \I__1106\ : InMux
    port map (
            O => \N__5052\,
            I => \N__5041\
        );

    \I__1105\ : InMux
    port map (
            O => \N__5051\,
            I => \N__5041\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__5046\,
            I => \uart_frame_decoder.state_1Z0Z_3\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__5041\,
            I => \uart_frame_decoder.state_1Z0Z_3\
        );

    \I__1102\ : CascadeMux
    port map (
            O => \N__5036\,
            I => \uart_frame_decoder.N_306_1_cascade_\
        );

    \I__1101\ : InMux
    port map (
            O => \N__5033\,
            I => \N__5027\
        );

    \I__1100\ : InMux
    port map (
            O => \N__5032\,
            I => \N__5021\
        );

    \I__1099\ : InMux
    port map (
            O => \N__5031\,
            I => \N__5021\
        );

    \I__1098\ : InMux
    port map (
            O => \N__5030\,
            I => \N__5018\
        );

    \I__1097\ : LocalMux
    port map (
            O => \N__5027\,
            I => \N__5014\
        );

    \I__1096\ : InMux
    port map (
            O => \N__5026\,
            I => \N__5011\
        );

    \I__1095\ : LocalMux
    port map (
            O => \N__5021\,
            I => \N__5003\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__5018\,
            I => \N__5003\
        );

    \I__1093\ : InMux
    port map (
            O => \N__5017\,
            I => \N__5000\
        );

    \I__1092\ : Span4Mux_s1_v
    port map (
            O => \N__5014\,
            I => \N__4995\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__5011\,
            I => \N__4995\
        );

    \I__1090\ : InMux
    port map (
            O => \N__5010\,
            I => \N__4990\
        );

    \I__1089\ : InMux
    port map (
            O => \N__5009\,
            I => \N__4990\
        );

    \I__1088\ : InMux
    port map (
            O => \N__5008\,
            I => \N__4987\
        );

    \I__1087\ : Span4Mux_h
    port map (
            O => \N__5003\,
            I => \N__4982\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__5000\,
            I => \N__4982\
        );

    \I__1085\ : Span4Mux_h
    port map (
            O => \N__4995\,
            I => \N__4979\
        );

    \I__1084\ : LocalMux
    port map (
            O => \N__4990\,
            I => \uart_frame_decoder.state_1Z0Z_10\
        );

    \I__1083\ : LocalMux
    port map (
            O => \N__4987\,
            I => \uart_frame_decoder.state_1Z0Z_10\
        );

    \I__1082\ : Odrv4
    port map (
            O => \N__4982\,
            I => \uart_frame_decoder.state_1Z0Z_10\
        );

    \I__1081\ : Odrv4
    port map (
            O => \N__4979\,
            I => \uart_frame_decoder.state_1Z0Z_10\
        );

    \I__1080\ : IoInMux
    port map (
            O => \N__4970\,
            I => \N__4967\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__4967\,
            I => \N__4964\
        );

    \I__1078\ : Span12Mux_s3_v
    port map (
            O => \N__4964\,
            I => \N__4961\
        );

    \I__1077\ : Odrv12
    port map (
            O => \N__4961\,
            I => \uart_frame_decoder_N_306_i\
        );

    \I__1076\ : InMux
    port map (
            O => \N__4958\,
            I => \uart_frame_decoder.un1_WDT_cry_14\
        );

    \I__1075\ : CascadeMux
    port map (
            O => \N__4955\,
            I => \N__4950\
        );

    \I__1074\ : InMux
    port map (
            O => \N__4954\,
            I => \N__4947\
        );

    \I__1073\ : InMux
    port map (
            O => \N__4953\,
            I => \N__4942\
        );

    \I__1072\ : InMux
    port map (
            O => \N__4950\,
            I => \N__4942\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__4947\,
            I => \uart_frame_decoder.WDTZ0Z_15\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__4942\,
            I => \uart_frame_decoder.WDTZ0Z_15\
        );

    \I__1069\ : InMux
    port map (
            O => \N__4937\,
            I => \N__4934\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__4934\,
            I => \N__4931\
        );

    \I__1067\ : Odrv4
    port map (
            O => \N__4931\,
            I => \uart_frame_decoder.state_1_ns_0_i_a2_0_0_0_10\
        );

    \I__1066\ : InMux
    port map (
            O => \N__4928\,
            I => \N__4924\
        );

    \I__1065\ : InMux
    port map (
            O => \N__4927\,
            I => \N__4921\
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__4924\,
            I => \uart_frame_decoder.state_1_ns_0_i_a2_0_d_10\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__4921\,
            I => \uart_frame_decoder.state_1_ns_0_i_a2_0_d_10\
        );

    \I__1062\ : InMux
    port map (
            O => \N__4916\,
            I => \N__4893\
        );

    \I__1061\ : InMux
    port map (
            O => \N__4915\,
            I => \N__4893\
        );

    \I__1060\ : InMux
    port map (
            O => \N__4914\,
            I => \N__4893\
        );

    \I__1059\ : InMux
    port map (
            O => \N__4913\,
            I => \N__4893\
        );

    \I__1058\ : InMux
    port map (
            O => \N__4912\,
            I => \N__4893\
        );

    \I__1057\ : InMux
    port map (
            O => \N__4911\,
            I => \N__4893\
        );

    \I__1056\ : InMux
    port map (
            O => \N__4910\,
            I => \N__4893\
        );

    \I__1055\ : InMux
    port map (
            O => \N__4909\,
            I => \N__4888\
        );

    \I__1054\ : InMux
    port map (
            O => \N__4908\,
            I => \N__4888\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__4893\,
            I => \uart_frame_decoder.N_85\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__4888\,
            I => \uart_frame_decoder.N_85\
        );

    \I__1051\ : ClkMux
    port map (
            O => \N__4883\,
            I => \N__4808\
        );

    \I__1050\ : ClkMux
    port map (
            O => \N__4882\,
            I => \N__4808\
        );

    \I__1049\ : ClkMux
    port map (
            O => \N__4881\,
            I => \N__4808\
        );

    \I__1048\ : ClkMux
    port map (
            O => \N__4880\,
            I => \N__4808\
        );

    \I__1047\ : ClkMux
    port map (
            O => \N__4879\,
            I => \N__4808\
        );

    \I__1046\ : ClkMux
    port map (
            O => \N__4878\,
            I => \N__4808\
        );

    \I__1045\ : ClkMux
    port map (
            O => \N__4877\,
            I => \N__4808\
        );

    \I__1044\ : ClkMux
    port map (
            O => \N__4876\,
            I => \N__4808\
        );

    \I__1043\ : ClkMux
    port map (
            O => \N__4875\,
            I => \N__4808\
        );

    \I__1042\ : ClkMux
    port map (
            O => \N__4874\,
            I => \N__4808\
        );

    \I__1041\ : ClkMux
    port map (
            O => \N__4873\,
            I => \N__4808\
        );

    \I__1040\ : ClkMux
    port map (
            O => \N__4872\,
            I => \N__4808\
        );

    \I__1039\ : ClkMux
    port map (
            O => \N__4871\,
            I => \N__4808\
        );

    \I__1038\ : ClkMux
    port map (
            O => \N__4870\,
            I => \N__4808\
        );

    \I__1037\ : ClkMux
    port map (
            O => \N__4869\,
            I => \N__4808\
        );

    \I__1036\ : ClkMux
    port map (
            O => \N__4868\,
            I => \N__4808\
        );

    \I__1035\ : ClkMux
    port map (
            O => \N__4867\,
            I => \N__4808\
        );

    \I__1034\ : ClkMux
    port map (
            O => \N__4866\,
            I => \N__4808\
        );

    \I__1033\ : ClkMux
    port map (
            O => \N__4865\,
            I => \N__4808\
        );

    \I__1032\ : ClkMux
    port map (
            O => \N__4864\,
            I => \N__4808\
        );

    \I__1031\ : ClkMux
    port map (
            O => \N__4863\,
            I => \N__4808\
        );

    \I__1030\ : ClkMux
    port map (
            O => \N__4862\,
            I => \N__4808\
        );

    \I__1029\ : ClkMux
    port map (
            O => \N__4861\,
            I => \N__4808\
        );

    \I__1028\ : ClkMux
    port map (
            O => \N__4860\,
            I => \N__4808\
        );

    \I__1027\ : ClkMux
    port map (
            O => \N__4859\,
            I => \N__4808\
        );

    \I__1026\ : GlobalMux
    port map (
            O => \N__4808\,
            I => \N__4805\
        );

    \I__1025\ : gio2CtrlBuf
    port map (
            O => \N__4805\,
            I => clk_system_c_g
        );

    \I__1024\ : InMux
    port map (
            O => \N__4802\,
            I => \N__4797\
        );

    \I__1023\ : InMux
    port map (
            O => \N__4801\,
            I => \N__4794\
        );

    \I__1022\ : InMux
    port map (
            O => \N__4800\,
            I => \N__4791\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__4797\,
            I => \uart_frame_decoder.WDTZ0Z_7\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__4794\,
            I => \uart_frame_decoder.WDTZ0Z_7\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__4791\,
            I => \uart_frame_decoder.WDTZ0Z_7\
        );

    \I__1018\ : InMux
    port map (
            O => \N__4784\,
            I => \uart_frame_decoder.un1_WDT_cry_6\
        );

    \I__1017\ : CascadeMux
    port map (
            O => \N__4781\,
            I => \N__4776\
        );

    \I__1016\ : InMux
    port map (
            O => \N__4780\,
            I => \N__4773\
        );

    \I__1015\ : InMux
    port map (
            O => \N__4779\,
            I => \N__4770\
        );

    \I__1014\ : InMux
    port map (
            O => \N__4776\,
            I => \N__4767\
        );

    \I__1013\ : LocalMux
    port map (
            O => \N__4773\,
            I => \N__4764\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__4770\,
            I => \uart_frame_decoder.WDTZ0Z_8\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__4767\,
            I => \uart_frame_decoder.WDTZ0Z_8\
        );

    \I__1010\ : Odrv4
    port map (
            O => \N__4764\,
            I => \uart_frame_decoder.WDTZ0Z_8\
        );

    \I__1009\ : InMux
    port map (
            O => \N__4757\,
            I => \bfn_12_3_0_\
        );

    \I__1008\ : InMux
    port map (
            O => \N__4754\,
            I => \N__4749\
        );

    \I__1007\ : InMux
    port map (
            O => \N__4753\,
            I => \N__4746\
        );

    \I__1006\ : InMux
    port map (
            O => \N__4752\,
            I => \N__4743\
        );

    \I__1005\ : LocalMux
    port map (
            O => \N__4749\,
            I => \uart_frame_decoder.WDTZ0Z_9\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__4746\,
            I => \uart_frame_decoder.WDTZ0Z_9\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__4743\,
            I => \uart_frame_decoder.WDTZ0Z_9\
        );

    \I__1002\ : InMux
    port map (
            O => \N__4736\,
            I => \uart_frame_decoder.un1_WDT_cry_8\
        );

    \I__1001\ : CascadeMux
    port map (
            O => \N__4733\,
            I => \N__4728\
        );

    \I__1000\ : InMux
    port map (
            O => \N__4732\,
            I => \N__4724\
        );

    \I__999\ : InMux
    port map (
            O => \N__4731\,
            I => \N__4719\
        );

    \I__998\ : InMux
    port map (
            O => \N__4728\,
            I => \N__4719\
        );

    \I__997\ : InMux
    port map (
            O => \N__4727\,
            I => \N__4716\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__4724\,
            I => \uart_frame_decoder.WDTZ0Z_10\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__4719\,
            I => \uart_frame_decoder.WDTZ0Z_10\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__4716\,
            I => \uart_frame_decoder.WDTZ0Z_10\
        );

    \I__993\ : InMux
    port map (
            O => \N__4709\,
            I => \uart_frame_decoder.un1_WDT_cry_9\
        );

    \I__992\ : InMux
    port map (
            O => \N__4706\,
            I => \N__4701\
        );

    \I__991\ : InMux
    port map (
            O => \N__4705\,
            I => \N__4698\
        );

    \I__990\ : InMux
    port map (
            O => \N__4704\,
            I => \N__4695\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__4701\,
            I => \uart_frame_decoder.WDTZ0Z_11\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__4698\,
            I => \uart_frame_decoder.WDTZ0Z_11\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__4695\,
            I => \uart_frame_decoder.WDTZ0Z_11\
        );

    \I__986\ : InMux
    port map (
            O => \N__4688\,
            I => \uart_frame_decoder.un1_WDT_cry_10\
        );

    \I__985\ : InMux
    port map (
            O => \N__4685\,
            I => \N__4680\
        );

    \I__984\ : InMux
    port map (
            O => \N__4684\,
            I => \N__4677\
        );

    \I__983\ : InMux
    port map (
            O => \N__4683\,
            I => \N__4674\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__4680\,
            I => \uart_frame_decoder.WDTZ0Z_12\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__4677\,
            I => \uart_frame_decoder.WDTZ0Z_12\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__4674\,
            I => \uart_frame_decoder.WDTZ0Z_12\
        );

    \I__979\ : InMux
    port map (
            O => \N__4667\,
            I => \uart_frame_decoder.un1_WDT_cry_11\
        );

    \I__978\ : CascadeMux
    port map (
            O => \N__4664\,
            I => \N__4658\
        );

    \I__977\ : InMux
    port map (
            O => \N__4663\,
            I => \N__4655\
        );

    \I__976\ : InMux
    port map (
            O => \N__4662\,
            I => \N__4648\
        );

    \I__975\ : InMux
    port map (
            O => \N__4661\,
            I => \N__4648\
        );

    \I__974\ : InMux
    port map (
            O => \N__4658\,
            I => \N__4648\
        );

    \I__973\ : LocalMux
    port map (
            O => \N__4655\,
            I => \uart_frame_decoder.WDTZ0Z_13\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__4648\,
            I => \uart_frame_decoder.WDTZ0Z_13\
        );

    \I__971\ : InMux
    port map (
            O => \N__4643\,
            I => \uart_frame_decoder.un1_WDT_cry_12\
        );

    \I__970\ : InMux
    port map (
            O => \N__4640\,
            I => \N__4634\
        );

    \I__969\ : InMux
    port map (
            O => \N__4639\,
            I => \N__4634\
        );

    \I__968\ : LocalMux
    port map (
            O => \N__4634\,
            I => \N__4627\
        );

    \I__967\ : InMux
    port map (
            O => \N__4633\,
            I => \N__4624\
        );

    \I__966\ : InMux
    port map (
            O => \N__4632\,
            I => \N__4617\
        );

    \I__965\ : InMux
    port map (
            O => \N__4631\,
            I => \N__4617\
        );

    \I__964\ : InMux
    port map (
            O => \N__4630\,
            I => \N__4617\
        );

    \I__963\ : Span4Mux_s1_v
    port map (
            O => \N__4627\,
            I => \N__4614\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__4624\,
            I => \uart_frame_decoder.WDTZ0Z_14\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__4617\,
            I => \uart_frame_decoder.WDTZ0Z_14\
        );

    \I__960\ : Odrv4
    port map (
            O => \N__4614\,
            I => \uart_frame_decoder.WDTZ0Z_14\
        );

    \I__959\ : InMux
    port map (
            O => \N__4607\,
            I => \uart_frame_decoder.un1_WDT_cry_13\
        );

    \I__958\ : InMux
    port map (
            O => \N__4604\,
            I => \N__4601\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__4601\,
            I => \N__4597\
        );

    \I__956\ : CascadeMux
    port map (
            O => \N__4600\,
            I => \N__4594\
        );

    \I__955\ : Span4Mux_h
    port map (
            O => \N__4597\,
            I => \N__4591\
        );

    \I__954\ : InMux
    port map (
            O => \N__4594\,
            I => \N__4588\
        );

    \I__953\ : Odrv4
    port map (
            O => \N__4591\,
            I => \uart.data_AuxZ0Z_4\
        );

    \I__952\ : LocalMux
    port map (
            O => \N__4588\,
            I => \uart.data_AuxZ0Z_4\
        );

    \I__951\ : InMux
    port map (
            O => \N__4583\,
            I => \N__4580\
        );

    \I__950\ : LocalMux
    port map (
            O => \N__4580\,
            I => \N__4577\
        );

    \I__949\ : Odrv4
    port map (
            O => \N__4577\,
            I => uart_data_4
        );

    \I__948\ : InMux
    port map (
            O => \N__4574\,
            I => \N__4571\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__4571\,
            I => \N__4567\
        );

    \I__946\ : InMux
    port map (
            O => \N__4570\,
            I => \N__4564\
        );

    \I__945\ : Odrv12
    port map (
            O => \N__4567\,
            I => \uart.data_AuxZ0Z_6\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__4564\,
            I => \uart.data_AuxZ0Z_6\
        );

    \I__943\ : InMux
    port map (
            O => \N__4559\,
            I => \N__4556\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__4556\,
            I => \N__4553\
        );

    \I__941\ : Span4Mux_s2_v
    port map (
            O => \N__4553\,
            I => \N__4550\
        );

    \I__940\ : Odrv4
    port map (
            O => \N__4550\,
            I => uart_data_6
        );

    \I__939\ : CEMux
    port map (
            O => \N__4547\,
            I => \N__4543\
        );

    \I__938\ : CEMux
    port map (
            O => \N__4546\,
            I => \N__4540\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__4543\,
            I => \N__4537\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__4540\,
            I => \N__4534\
        );

    \I__935\ : Odrv4
    port map (
            O => \N__4537\,
            I => \uart.state_1_sqmuxa_0\
        );

    \I__934\ : Odrv4
    port map (
            O => \N__4534\,
            I => \uart.state_1_sqmuxa_0\
        );

    \I__933\ : SRMux
    port map (
            O => \N__4529\,
            I => \N__4525\
        );

    \I__932\ : SRMux
    port map (
            O => \N__4528\,
            I => \N__4522\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__4525\,
            I => \N__4519\
        );

    \I__930\ : LocalMux
    port map (
            O => \N__4522\,
            I => \N__4516\
        );

    \I__929\ : Span4Mux_s3_v
    port map (
            O => \N__4519\,
            I => \N__4512\
        );

    \I__928\ : Span4Mux_h
    port map (
            O => \N__4516\,
            I => \N__4509\
        );

    \I__927\ : InMux
    port map (
            O => \N__4515\,
            I => \N__4506\
        );

    \I__926\ : Odrv4
    port map (
            O => \N__4512\,
            I => \uart.timer_Count_RNIS4183Z0Z_7\
        );

    \I__925\ : Odrv4
    port map (
            O => \N__4509\,
            I => \uart.timer_Count_RNIS4183Z0Z_7\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__4506\,
            I => \uart.timer_Count_RNIS4183Z0Z_7\
        );

    \I__923\ : InMux
    port map (
            O => \N__4499\,
            I => \N__4495\
        );

    \I__922\ : CascadeMux
    port map (
            O => \N__4498\,
            I => \N__4492\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__4495\,
            I => \N__4489\
        );

    \I__920\ : InMux
    port map (
            O => \N__4492\,
            I => \N__4486\
        );

    \I__919\ : Odrv4
    port map (
            O => \N__4489\,
            I => \uart_frame_decoder.WDT8_0_i\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__4486\,
            I => \uart_frame_decoder.WDT8_0_i\
        );

    \I__917\ : InMux
    port map (
            O => \N__4481\,
            I => \N__4478\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__4478\,
            I => \uart_frame_decoder.WDTZ0Z_0\
        );

    \I__915\ : InMux
    port map (
            O => \N__4475\,
            I => \N__4472\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__4472\,
            I => \uart_frame_decoder.WDTZ0Z_1\
        );

    \I__913\ : InMux
    port map (
            O => \N__4469\,
            I => \uart_frame_decoder.un1_WDT_cry_0\
        );

    \I__912\ : InMux
    port map (
            O => \N__4466\,
            I => \N__4463\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__4463\,
            I => \uart_frame_decoder.WDTZ0Z_2\
        );

    \I__910\ : InMux
    port map (
            O => \N__4460\,
            I => \uart_frame_decoder.un1_WDT_cry_1\
        );

    \I__909\ : InMux
    port map (
            O => \N__4457\,
            I => \N__4454\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__4454\,
            I => \uart_frame_decoder.WDTZ0Z_3\
        );

    \I__907\ : InMux
    port map (
            O => \N__4451\,
            I => \uart_frame_decoder.un1_WDT_cry_2\
        );

    \I__906\ : InMux
    port map (
            O => \N__4448\,
            I => \N__4443\
        );

    \I__905\ : InMux
    port map (
            O => \N__4447\,
            I => \N__4438\
        );

    \I__904\ : InMux
    port map (
            O => \N__4446\,
            I => \N__4438\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__4443\,
            I => \uart_frame_decoder.WDTZ0Z_4\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__4438\,
            I => \uart_frame_decoder.WDTZ0Z_4\
        );

    \I__901\ : InMux
    port map (
            O => \N__4433\,
            I => \uart_frame_decoder.un1_WDT_cry_3\
        );

    \I__900\ : CascadeMux
    port map (
            O => \N__4430\,
            I => \N__4427\
        );

    \I__899\ : InMux
    port map (
            O => \N__4427\,
            I => \N__4422\
        );

    \I__898\ : InMux
    port map (
            O => \N__4426\,
            I => \N__4419\
        );

    \I__897\ : InMux
    port map (
            O => \N__4425\,
            I => \N__4416\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__4422\,
            I => \N__4413\
        );

    \I__895\ : LocalMux
    port map (
            O => \N__4419\,
            I => \uart_frame_decoder.WDTZ0Z_5\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__4416\,
            I => \uart_frame_decoder.WDTZ0Z_5\
        );

    \I__893\ : Odrv4
    port map (
            O => \N__4413\,
            I => \uart_frame_decoder.WDTZ0Z_5\
        );

    \I__892\ : InMux
    port map (
            O => \N__4406\,
            I => \uart_frame_decoder.un1_WDT_cry_4\
        );

    \I__891\ : CascadeMux
    port map (
            O => \N__4403\,
            I => \N__4398\
        );

    \I__890\ : InMux
    port map (
            O => \N__4402\,
            I => \N__4395\
        );

    \I__889\ : InMux
    port map (
            O => \N__4401\,
            I => \N__4392\
        );

    \I__888\ : InMux
    port map (
            O => \N__4398\,
            I => \N__4389\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__4395\,
            I => \uart_frame_decoder.WDTZ0Z_6\
        );

    \I__886\ : LocalMux
    port map (
            O => \N__4392\,
            I => \uart_frame_decoder.WDTZ0Z_6\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__4389\,
            I => \uart_frame_decoder.WDTZ0Z_6\
        );

    \I__884\ : InMux
    port map (
            O => \N__4382\,
            I => \uart_frame_decoder.un1_WDT_cry_5\
        );

    \I__883\ : InMux
    port map (
            O => \N__4379\,
            I => \N__4376\
        );

    \I__882\ : LocalMux
    port map (
            O => \N__4376\,
            I => \uart_frame_decoder.WDT_RNIQAB11Z0Z_4\
        );

    \I__881\ : CascadeMux
    port map (
            O => \N__4373\,
            I => \uart_frame_decoder.WDT_RNISS5HZ0Z_11_cascade_\
        );

    \I__880\ : CascadeMux
    port map (
            O => \N__4370\,
            I => \uart_frame_decoder.WDT8lt13_cascade_\
        );

    \I__879\ : InMux
    port map (
            O => \N__4367\,
            I => \N__4364\
        );

    \I__878\ : LocalMux
    port map (
            O => \N__4364\,
            I => \uart_frame_decoder.state_1_ns_i_i_a2_0_0\
        );

    \I__877\ : CascadeMux
    port map (
            O => \N__4361\,
            I => \N__4358\
        );

    \I__876\ : InMux
    port map (
            O => \N__4358\,
            I => \N__4352\
        );

    \I__875\ : InMux
    port map (
            O => \N__4357\,
            I => \N__4352\
        );

    \I__874\ : LocalMux
    port map (
            O => \N__4352\,
            I => \uart_frame_decoder.WDT8lt13\
        );

    \I__873\ : CascadeMux
    port map (
            O => \N__4349\,
            I => \N__4346\
        );

    \I__872\ : InMux
    port map (
            O => \N__4346\,
            I => \N__4342\
        );

    \I__871\ : InMux
    port map (
            O => \N__4345\,
            I => \N__4339\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__4342\,
            I => \uart_frame_decoder.WDT8lto15\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__4339\,
            I => \uart_frame_decoder.WDT8lto15\
        );

    \I__868\ : InMux
    port map (
            O => \N__4334\,
            I => \N__4331\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__4331\,
            I => \uart_frame_decoder.N_80\
        );

    \I__866\ : CascadeMux
    port map (
            O => \N__4328\,
            I => \N__4325\
        );

    \I__865\ : InMux
    port map (
            O => \N__4325\,
            I => \N__4321\
        );

    \I__864\ : InMux
    port map (
            O => \N__4324\,
            I => \N__4316\
        );

    \I__863\ : LocalMux
    port map (
            O => \N__4321\,
            I => \N__4313\
        );

    \I__862\ : InMux
    port map (
            O => \N__4320\,
            I => \N__4308\
        );

    \I__861\ : InMux
    port map (
            O => \N__4319\,
            I => \N__4308\
        );

    \I__860\ : LocalMux
    port map (
            O => \N__4316\,
            I => \N__4305\
        );

    \I__859\ : Span4Mux_h
    port map (
            O => \N__4313\,
            I => \N__4302\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__4308\,
            I => \uart.timer_CountZ0Z_0\
        );

    \I__857\ : Odrv4
    port map (
            O => \N__4305\,
            I => \uart.timer_CountZ0Z_0\
        );

    \I__856\ : Odrv4
    port map (
            O => \N__4302\,
            I => \uart.timer_CountZ0Z_0\
        );

    \I__855\ : SRMux
    port map (
            O => \N__4295\,
            I => \N__4291\
        );

    \I__854\ : SRMux
    port map (
            O => \N__4294\,
            I => \N__4288\
        );

    \I__853\ : LocalMux
    port map (
            O => \N__4291\,
            I => \uart.timer_Count_1_sqmuxa_i\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__4288\,
            I => \uart.timer_Count_1_sqmuxa_i\
        );

    \I__851\ : CascadeMux
    port map (
            O => \N__4283\,
            I => \N__4280\
        );

    \I__850\ : InMux
    port map (
            O => \N__4280\,
            I => \N__4277\
        );

    \I__849\ : LocalMux
    port map (
            O => \N__4277\,
            I => \uart_frame_decoder.state_1_ns_0_i_a2_0_0_1\
        );

    \I__848\ : CascadeMux
    port map (
            O => \N__4274\,
            I => \N__4271\
        );

    \I__847\ : InMux
    port map (
            O => \N__4271\,
            I => \N__4264\
        );

    \I__846\ : InMux
    port map (
            O => \N__4270\,
            I => \N__4264\
        );

    \I__845\ : InMux
    port map (
            O => \N__4269\,
            I => \N__4261\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__4264\,
            I => \uart_frame_decoder.N_99\
        );

    \I__843\ : LocalMux
    port map (
            O => \N__4261\,
            I => \uart_frame_decoder.N_99\
        );

    \I__842\ : InMux
    port map (
            O => \N__4256\,
            I => \N__4252\
        );

    \I__841\ : InMux
    port map (
            O => \N__4255\,
            I => \N__4249\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__4252\,
            I => \uart_frame_decoder.N_92\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__4249\,
            I => \uart_frame_decoder.N_92\
        );

    \I__838\ : InMux
    port map (
            O => \N__4244\,
            I => \N__4241\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__4241\,
            I => \N__4237\
        );

    \I__836\ : CascadeMux
    port map (
            O => \N__4240\,
            I => \N__4234\
        );

    \I__835\ : Span4Mux_v
    port map (
            O => \N__4237\,
            I => \N__4231\
        );

    \I__834\ : InMux
    port map (
            O => \N__4234\,
            I => \N__4228\
        );

    \I__833\ : Odrv4
    port map (
            O => \N__4231\,
            I => \uart.data_AuxZ0Z_1\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__4228\,
            I => \uart.data_AuxZ0Z_1\
        );

    \I__831\ : InMux
    port map (
            O => \N__4223\,
            I => \N__4220\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__4220\,
            I => \N__4217\
        );

    \I__829\ : Odrv4
    port map (
            O => \N__4217\,
            I => uart_data_1
        );

    \I__828\ : CascadeMux
    port map (
            O => \N__4214\,
            I => \uart_frame_decoder.N_4_0_cascade_\
        );

    \I__827\ : InMux
    port map (
            O => \N__4211\,
            I => \N__4208\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__4208\,
            I => \uart_frame_decoder.g0_1_0_1\
        );

    \I__825\ : InMux
    port map (
            O => \N__4205\,
            I => \N__4202\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__4202\,
            I => \uart_frame_decoder.g0_1_a3_3\
        );

    \I__823\ : CascadeMux
    port map (
            O => \N__4199\,
            I => \uart_frame_decoder.WDT8lto15_cascade_\
        );

    \I__822\ : InMux
    port map (
            O => \N__4196\,
            I => \N__4193\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__4193\,
            I => \uart_frame_decoder.state_1_ns_0_i_o2_0_tz_10\
        );

    \I__820\ : InMux
    port map (
            O => \N__4190\,
            I => \N__4187\
        );

    \I__819\ : LocalMux
    port map (
            O => \N__4187\,
            I => \uart_frame_decoder.state_1_ns_i_i_a2_1_1_0\
        );

    \I__818\ : InMux
    port map (
            O => \N__4184\,
            I => \N__4179\
        );

    \I__817\ : InMux
    port map (
            O => \N__4183\,
            I => \N__4174\
        );

    \I__816\ : InMux
    port map (
            O => \N__4182\,
            I => \N__4174\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__4179\,
            I => \uart_frame_decoder.state_1Z0Z_0\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__4174\,
            I => \uart_frame_decoder.state_1Z0Z_0\
        );

    \I__813\ : CascadeMux
    port map (
            O => \N__4169\,
            I => \uart_frame_decoder.state_1_ns_0_i_a2_0_0_0_10_cascade_\
        );

    \I__812\ : InMux
    port map (
            O => \N__4166\,
            I => \N__4163\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__4163\,
            I => \uart_frame_decoder.N_35_i_1\
        );

    \I__810\ : CascadeMux
    port map (
            O => \N__4160\,
            I => \N__4157\
        );

    \I__809\ : InMux
    port map (
            O => \N__4157\,
            I => \N__4152\
        );

    \I__808\ : InMux
    port map (
            O => \N__4156\,
            I => \N__4149\
        );

    \I__807\ : InMux
    port map (
            O => \N__4155\,
            I => \N__4145\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__4152\,
            I => \N__4142\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__4149\,
            I => \N__4139\
        );

    \I__804\ : InMux
    port map (
            O => \N__4148\,
            I => \N__4136\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__4145\,
            I => \uart.timer_CountZ0Z_1\
        );

    \I__802\ : Odrv4
    port map (
            O => \N__4142\,
            I => \uart.timer_CountZ0Z_1\
        );

    \I__801\ : Odrv12
    port map (
            O => \N__4139\,
            I => \uart.timer_CountZ0Z_1\
        );

    \I__800\ : LocalMux
    port map (
            O => \N__4136\,
            I => \uart.timer_CountZ0Z_1\
        );

    \I__799\ : CascadeMux
    port map (
            O => \N__4127\,
            I => \N__4124\
        );

    \I__798\ : InMux
    port map (
            O => \N__4124\,
            I => \N__4121\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__4121\,
            I => \uart_frame_decoder.count8_axb_1\
        );

    \I__796\ : CascadeMux
    port map (
            O => \N__4118\,
            I => \N__4115\
        );

    \I__795\ : InMux
    port map (
            O => \N__4115\,
            I => \N__4112\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__4112\,
            I => \uart_frame_decoder.count_i_2\
        );

    \I__793\ : InMux
    port map (
            O => \N__4109\,
            I => \uart_frame_decoder.count8\
        );

    \I__792\ : InMux
    port map (
            O => \N__4106\,
            I => \N__4103\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__4103\,
            I => \N__4100\
        );

    \I__790\ : Odrv12
    port map (
            O => \N__4100\,
            I => \uart_frame_decoder.count8_THRU_CO\
        );

    \I__789\ : CascadeMux
    port map (
            O => \N__4097\,
            I => \uart_frame_decoder.count8_THRU_CO_cascade_\
        );

    \I__788\ : InMux
    port map (
            O => \N__4094\,
            I => \N__4088\
        );

    \I__787\ : InMux
    port map (
            O => \N__4093\,
            I => \N__4088\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__4088\,
            I => \uart_frame_decoder.N_37\
        );

    \I__785\ : CascadeMux
    port map (
            O => \N__4085\,
            I => \uart_frame_decoder.N_37_cascade_\
        );

    \I__784\ : CascadeMux
    port map (
            O => \N__4082\,
            I => \N__4077\
        );

    \I__783\ : InMux
    port map (
            O => \N__4081\,
            I => \N__4071\
        );

    \I__782\ : InMux
    port map (
            O => \N__4080\,
            I => \N__4071\
        );

    \I__781\ : InMux
    port map (
            O => \N__4077\,
            I => \N__4066\
        );

    \I__780\ : InMux
    port map (
            O => \N__4076\,
            I => \N__4066\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__4071\,
            I => \uart_frame_decoder.countZ0Z_1\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__4066\,
            I => \uart_frame_decoder.countZ0Z_1\
        );

    \I__777\ : InMux
    port map (
            O => \N__4061\,
            I => \N__4056\
        );

    \I__776\ : InMux
    port map (
            O => \N__4060\,
            I => \N__4051\
        );

    \I__775\ : InMux
    port map (
            O => \N__4059\,
            I => \N__4051\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__4056\,
            I => \uart_frame_decoder.countZ0Z_2\
        );

    \I__773\ : LocalMux
    port map (
            O => \N__4051\,
            I => \uart_frame_decoder.countZ0Z_2\
        );

    \I__772\ : InMux
    port map (
            O => \N__4046\,
            I => \N__4040\
        );

    \I__771\ : InMux
    port map (
            O => \N__4045\,
            I => \N__4040\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__4040\,
            I => \CONSTANT_ONE_NET\
        );

    \I__769\ : InMux
    port map (
            O => \N__4037\,
            I => \N__4031\
        );

    \I__768\ : InMux
    port map (
            O => \N__4036\,
            I => \N__4024\
        );

    \I__767\ : InMux
    port map (
            O => \N__4035\,
            I => \N__4024\
        );

    \I__766\ : InMux
    port map (
            O => \N__4034\,
            I => \N__4024\
        );

    \I__765\ : LocalMux
    port map (
            O => \N__4031\,
            I => \uart_frame_decoder.count8_0\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__4024\,
            I => \uart_frame_decoder.count8_0\
        );

    \I__763\ : CascadeMux
    port map (
            O => \N__4019\,
            I => \N__4015\
        );

    \I__762\ : InMux
    port map (
            O => \N__4018\,
            I => \N__4010\
        );

    \I__761\ : InMux
    port map (
            O => \N__4015\,
            I => \N__4010\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__4010\,
            I => \uart_frame_decoder.count8_0_i\
        );

    \I__759\ : InMux
    port map (
            O => \N__4007\,
            I => \N__4004\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__4004\,
            I => \N__3997\
        );

    \I__757\ : InMux
    port map (
            O => \N__4003\,
            I => \N__3994\
        );

    \I__756\ : InMux
    port map (
            O => \N__4002\,
            I => \N__3987\
        );

    \I__755\ : InMux
    port map (
            O => \N__4001\,
            I => \N__3987\
        );

    \I__754\ : InMux
    port map (
            O => \N__4000\,
            I => \N__3987\
        );

    \I__753\ : Odrv4
    port map (
            O => \N__3997\,
            I => \uart.N_145_0\
        );

    \I__752\ : LocalMux
    port map (
            O => \N__3994\,
            I => \uart.N_145_0\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__3987\,
            I => \uart.N_145_0\
        );

    \I__750\ : InMux
    port map (
            O => \N__3980\,
            I => \N__3977\
        );

    \I__749\ : LocalMux
    port map (
            O => \N__3977\,
            I => \uart.state_1_sqmuxa\
        );

    \I__748\ : CascadeMux
    port map (
            O => \N__3974\,
            I => \uart.state_1_sqmuxa_cascade_\
        );

    \I__747\ : InMux
    port map (
            O => \N__3971\,
            I => \N__3968\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__3968\,
            I => \N__3961\
        );

    \I__745\ : InMux
    port map (
            O => \N__3967\,
            I => \N__3958\
        );

    \I__744\ : InMux
    port map (
            O => \N__3966\,
            I => \N__3955\
        );

    \I__743\ : InMux
    port map (
            O => \N__3965\,
            I => \N__3952\
        );

    \I__742\ : InMux
    port map (
            O => \N__3964\,
            I => \N__3949\
        );

    \I__741\ : Span4Mux_v
    port map (
            O => \N__3961\,
            I => \N__3946\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__3958\,
            I => \N__3941\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__3955\,
            I => \N__3941\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__3952\,
            I => \uart.timer_CountZ0Z_2\
        );

    \I__737\ : LocalMux
    port map (
            O => \N__3949\,
            I => \uart.timer_CountZ0Z_2\
        );

    \I__736\ : Odrv4
    port map (
            O => \N__3946\,
            I => \uart.timer_CountZ0Z_2\
        );

    \I__735\ : Odrv4
    port map (
            O => \N__3941\,
            I => \uart.timer_CountZ0Z_2\
        );

    \I__734\ : InMux
    port map (
            O => \N__3932\,
            I => \uart.un4_timer_Count_1_cry_1\
        );

    \I__733\ : InMux
    port map (
            O => \N__3929\,
            I => \N__3926\
        );

    \I__732\ : LocalMux
    port map (
            O => \N__3926\,
            I => \N__3921\
        );

    \I__731\ : InMux
    port map (
            O => \N__3925\,
            I => \N__3916\
        );

    \I__730\ : InMux
    port map (
            O => \N__3924\,
            I => \N__3913\
        );

    \I__729\ : Span4Mux_h
    port map (
            O => \N__3921\,
            I => \N__3910\
        );

    \I__728\ : InMux
    port map (
            O => \N__3920\,
            I => \N__3907\
        );

    \I__727\ : InMux
    port map (
            O => \N__3919\,
            I => \N__3904\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__3916\,
            I => \uart.timer_CountZ0Z_3\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__3913\,
            I => \uart.timer_CountZ0Z_3\
        );

    \I__724\ : Odrv4
    port map (
            O => \N__3910\,
            I => \uart.timer_CountZ0Z_3\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__3907\,
            I => \uart.timer_CountZ0Z_3\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__3904\,
            I => \uart.timer_CountZ0Z_3\
        );

    \I__721\ : InMux
    port map (
            O => \N__3893\,
            I => \uart.un4_timer_Count_1_cry_2\
        );

    \I__720\ : InMux
    port map (
            O => \N__3890\,
            I => \N__3887\
        );

    \I__719\ : LocalMux
    port map (
            O => \N__3887\,
            I => \N__3881\
        );

    \I__718\ : CascadeMux
    port map (
            O => \N__3886\,
            I => \N__3877\
        );

    \I__717\ : InMux
    port map (
            O => \N__3885\,
            I => \N__3874\
        );

    \I__716\ : InMux
    port map (
            O => \N__3884\,
            I => \N__3871\
        );

    \I__715\ : Span4Mux_h
    port map (
            O => \N__3881\,
            I => \N__3868\
        );

    \I__714\ : InMux
    port map (
            O => \N__3880\,
            I => \N__3865\
        );

    \I__713\ : InMux
    port map (
            O => \N__3877\,
            I => \N__3862\
        );

    \I__712\ : LocalMux
    port map (
            O => \N__3874\,
            I => \uart.timer_CountZ0Z_4\
        );

    \I__711\ : LocalMux
    port map (
            O => \N__3871\,
            I => \uart.timer_CountZ0Z_4\
        );

    \I__710\ : Odrv4
    port map (
            O => \N__3868\,
            I => \uart.timer_CountZ0Z_4\
        );

    \I__709\ : LocalMux
    port map (
            O => \N__3865\,
            I => \uart.timer_CountZ0Z_4\
        );

    \I__708\ : LocalMux
    port map (
            O => \N__3862\,
            I => \uart.timer_CountZ0Z_4\
        );

    \I__707\ : InMux
    port map (
            O => \N__3851\,
            I => \uart.un4_timer_Count_1_cry_3\
        );

    \I__706\ : InMux
    port map (
            O => \N__3848\,
            I => \N__3844\
        );

    \I__705\ : InMux
    port map (
            O => \N__3847\,
            I => \N__3838\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__3844\,
            I => \N__3835\
        );

    \I__703\ : InMux
    port map (
            O => \N__3843\,
            I => \N__3828\
        );

    \I__702\ : InMux
    port map (
            O => \N__3842\,
            I => \N__3828\
        );

    \I__701\ : InMux
    port map (
            O => \N__3841\,
            I => \N__3828\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__3838\,
            I => \uart.timer_CountZ0Z_5\
        );

    \I__699\ : Odrv4
    port map (
            O => \N__3835\,
            I => \uart.timer_CountZ0Z_5\
        );

    \I__698\ : LocalMux
    port map (
            O => \N__3828\,
            I => \uart.timer_CountZ0Z_5\
        );

    \I__697\ : InMux
    port map (
            O => \N__3821\,
            I => \uart.un4_timer_Count_1_cry_4\
        );

    \I__696\ : InMux
    port map (
            O => \N__3818\,
            I => \N__3814\
        );

    \I__695\ : InMux
    port map (
            O => \N__3817\,
            I => \N__3809\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__3814\,
            I => \N__3806\
        );

    \I__693\ : InMux
    port map (
            O => \N__3813\,
            I => \N__3801\
        );

    \I__692\ : InMux
    port map (
            O => \N__3812\,
            I => \N__3801\
        );

    \I__691\ : LocalMux
    port map (
            O => \N__3809\,
            I => \uart.timer_CountZ0Z_6\
        );

    \I__690\ : Odrv4
    port map (
            O => \N__3806\,
            I => \uart.timer_CountZ0Z_6\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__3801\,
            I => \uart.timer_CountZ0Z_6\
        );

    \I__688\ : InMux
    port map (
            O => \N__3794\,
            I => \uart.un4_timer_Count_1_cry_5\
        );

    \I__687\ : InMux
    port map (
            O => \N__3791\,
            I => \uart.un4_timer_Count_1_cry_6\
        );

    \I__686\ : InMux
    port map (
            O => \N__3788\,
            I => \N__3784\
        );

    \I__685\ : InMux
    port map (
            O => \N__3787\,
            I => \N__3781\
        );

    \I__684\ : LocalMux
    port map (
            O => \N__3784\,
            I => \N__3774\
        );

    \I__683\ : LocalMux
    port map (
            O => \N__3781\,
            I => \N__3774\
        );

    \I__682\ : CascadeMux
    port map (
            O => \N__3780\,
            I => \N__3767\
        );

    \I__681\ : InMux
    port map (
            O => \N__3779\,
            I => \N__3764\
        );

    \I__680\ : Span4Mux_s1_v
    port map (
            O => \N__3774\,
            I => \N__3761\
        );

    \I__679\ : InMux
    port map (
            O => \N__3773\,
            I => \N__3754\
        );

    \I__678\ : InMux
    port map (
            O => \N__3772\,
            I => \N__3754\
        );

    \I__677\ : InMux
    port map (
            O => \N__3771\,
            I => \N__3754\
        );

    \I__676\ : InMux
    port map (
            O => \N__3770\,
            I => \N__3749\
        );

    \I__675\ : InMux
    port map (
            O => \N__3767\,
            I => \N__3749\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__3764\,
            I => \uart.timer_CountZ0Z_7\
        );

    \I__673\ : Odrv4
    port map (
            O => \N__3761\,
            I => \uart.timer_CountZ0Z_7\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__3754\,
            I => \uart.timer_CountZ0Z_7\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__3749\,
            I => \uart.timer_CountZ0Z_7\
        );

    \I__670\ : InMux
    port map (
            O => \N__3740\,
            I => \N__3737\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__3737\,
            I => uart_data_3
        );

    \I__668\ : CascadeMux
    port map (
            O => \N__3734\,
            I => \uart_frame_decoder.state_1_ns_0_i_a2_1_0Z0Z_2_cascade_\
        );

    \I__667\ : InMux
    port map (
            O => \N__3731\,
            I => \N__3725\
        );

    \I__666\ : InMux
    port map (
            O => \N__3730\,
            I => \N__3725\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__3725\,
            I => uart_data_2
        );

    \I__664\ : InMux
    port map (
            O => \N__3722\,
            I => \N__3716\
        );

    \I__663\ : InMux
    port map (
            O => \N__3721\,
            I => \N__3716\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__3716\,
            I => uart_data_5
        );

    \I__661\ : CascadeMux
    port map (
            O => \N__3713\,
            I => \N__3710\
        );

    \I__660\ : InMux
    port map (
            O => \N__3710\,
            I => \N__3704\
        );

    \I__659\ : InMux
    port map (
            O => \N__3709\,
            I => \N__3704\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__3704\,
            I => uart_data_7
        );

    \I__657\ : InMux
    port map (
            O => \N__3701\,
            I => \N__3695\
        );

    \I__656\ : InMux
    port map (
            O => \N__3700\,
            I => \N__3695\
        );

    \I__655\ : LocalMux
    port map (
            O => \N__3695\,
            I => uart_data_0
        );

    \I__654\ : InMux
    port map (
            O => \N__3692\,
            I => \N__3689\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__3689\,
            I => \uart_frame_decoder.N_79_4\
        );

    \I__652\ : CascadeMux
    port map (
            O => \N__3686\,
            I => \uart_frame_decoder.N_79_4_cascade_\
        );

    \I__651\ : CascadeMux
    port map (
            O => \N__3683\,
            I => \N__3678\
        );

    \I__650\ : CascadeMux
    port map (
            O => \N__3682\,
            I => \N__3673\
        );

    \I__649\ : InMux
    port map (
            O => \N__3681\,
            I => \N__3665\
        );

    \I__648\ : InMux
    port map (
            O => \N__3678\,
            I => \N__3662\
        );

    \I__647\ : InMux
    port map (
            O => \N__3677\,
            I => \N__3659\
        );

    \I__646\ : InMux
    port map (
            O => \N__3676\,
            I => \N__3656\
        );

    \I__645\ : InMux
    port map (
            O => \N__3673\,
            I => \N__3653\
        );

    \I__644\ : InMux
    port map (
            O => \N__3672\,
            I => \N__3647\
        );

    \I__643\ : InMux
    port map (
            O => \N__3671\,
            I => \N__3638\
        );

    \I__642\ : InMux
    port map (
            O => \N__3670\,
            I => \N__3638\
        );

    \I__641\ : InMux
    port map (
            O => \N__3669\,
            I => \N__3638\
        );

    \I__640\ : InMux
    port map (
            O => \N__3668\,
            I => \N__3638\
        );

    \I__639\ : LocalMux
    port map (
            O => \N__3665\,
            I => \N__3635\
        );

    \I__638\ : LocalMux
    port map (
            O => \N__3662\,
            I => \N__3626\
        );

    \I__637\ : LocalMux
    port map (
            O => \N__3659\,
            I => \N__3626\
        );

    \I__636\ : LocalMux
    port map (
            O => \N__3656\,
            I => \N__3626\
        );

    \I__635\ : LocalMux
    port map (
            O => \N__3653\,
            I => \N__3626\
        );

    \I__634\ : InMux
    port map (
            O => \N__3652\,
            I => \N__3619\
        );

    \I__633\ : InMux
    port map (
            O => \N__3651\,
            I => \N__3619\
        );

    \I__632\ : InMux
    port map (
            O => \N__3650\,
            I => \N__3619\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__3647\,
            I => \N__3616\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__3638\,
            I => \N__3613\
        );

    \I__629\ : Span4Mux_s1_v
    port map (
            O => \N__3635\,
            I => \N__3608\
        );

    \I__628\ : Span4Mux_v
    port map (
            O => \N__3626\,
            I => \N__3608\
        );

    \I__627\ : LocalMux
    port map (
            O => \N__3619\,
            I => uart_input_sync
        );

    \I__626\ : Odrv4
    port map (
            O => \N__3616\,
            I => uart_input_sync
        );

    \I__625\ : Odrv4
    port map (
            O => \N__3613\,
            I => uart_input_sync
        );

    \I__624\ : Odrv4
    port map (
            O => \N__3608\,
            I => uart_input_sync
        );

    \I__623\ : CascadeMux
    port map (
            O => \N__3599\,
            I => \uart.data_8_0_cascade_\
        );

    \I__622\ : InMux
    port map (
            O => \N__3596\,
            I => \N__3593\
        );

    \I__621\ : LocalMux
    port map (
            O => \N__3593\,
            I => \uart.state_srsts_0_a3_1_4\
        );

    \I__620\ : CascadeMux
    port map (
            O => \N__3590\,
            I => \uart.N_152_0_cascade_\
        );

    \I__619\ : InMux
    port map (
            O => \N__3587\,
            I => \N__3584\
        );

    \I__618\ : LocalMux
    port map (
            O => \N__3584\,
            I => \uart.N_167\
        );

    \I__617\ : InMux
    port map (
            O => \N__3581\,
            I => \N__3578\
        );

    \I__616\ : LocalMux
    port map (
            O => \N__3578\,
            I => \uart.N_159\
        );

    \I__615\ : CascadeMux
    port map (
            O => \N__3575\,
            I => \uart.N_167_cascade_\
        );

    \I__614\ : InMux
    port map (
            O => \N__3572\,
            I => \N__3568\
        );

    \I__613\ : InMux
    port map (
            O => \N__3571\,
            I => \N__3562\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__3568\,
            I => \N__3559\
        );

    \I__611\ : InMux
    port map (
            O => \N__3567\,
            I => \N__3556\
        );

    \I__610\ : InMux
    port map (
            O => \N__3566\,
            I => \N__3553\
        );

    \I__609\ : InMux
    port map (
            O => \N__3565\,
            I => \N__3550\
        );

    \I__608\ : LocalMux
    port map (
            O => \N__3562\,
            I => \uart.N_180\
        );

    \I__607\ : Odrv4
    port map (
            O => \N__3559\,
            I => \uart.N_180\
        );

    \I__606\ : LocalMux
    port map (
            O => \N__3556\,
            I => \uart.N_180\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__3553\,
            I => \uart.N_180\
        );

    \I__604\ : LocalMux
    port map (
            O => \N__3550\,
            I => \uart.N_180\
        );

    \I__603\ : InMux
    port map (
            O => \N__3539\,
            I => \N__3536\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__3536\,
            I => \N__3531\
        );

    \I__601\ : InMux
    port map (
            O => \N__3535\,
            I => \N__3526\
        );

    \I__600\ : InMux
    port map (
            O => \N__3534\,
            I => \N__3526\
        );

    \I__599\ : Odrv4
    port map (
            O => \N__3531\,
            I => \uart.N_152_0\
        );

    \I__598\ : LocalMux
    port map (
            O => \N__3526\,
            I => \uart.N_152_0\
        );

    \I__597\ : InMux
    port map (
            O => \N__3521\,
            I => \N__3517\
        );

    \I__596\ : InMux
    port map (
            O => \N__3520\,
            I => \N__3514\
        );

    \I__595\ : LocalMux
    port map (
            O => \N__3517\,
            I => \N__3506\
        );

    \I__594\ : LocalMux
    port map (
            O => \N__3514\,
            I => \N__3506\
        );

    \I__593\ : CascadeMux
    port map (
            O => \N__3513\,
            I => \N__3502\
        );

    \I__592\ : InMux
    port map (
            O => \N__3512\,
            I => \N__3497\
        );

    \I__591\ : InMux
    port map (
            O => \N__3511\,
            I => \N__3494\
        );

    \I__590\ : Span4Mux_s1_v
    port map (
            O => \N__3506\,
            I => \N__3491\
        );

    \I__589\ : InMux
    port map (
            O => \N__3505\,
            I => \N__3488\
        );

    \I__588\ : InMux
    port map (
            O => \N__3502\,
            I => \N__3483\
        );

    \I__587\ : InMux
    port map (
            O => \N__3501\,
            I => \N__3483\
        );

    \I__586\ : InMux
    port map (
            O => \N__3500\,
            I => \N__3480\
        );

    \I__585\ : LocalMux
    port map (
            O => \N__3497\,
            I => \uart.stateZ0Z_4\
        );

    \I__584\ : LocalMux
    port map (
            O => \N__3494\,
            I => \uart.stateZ0Z_4\
        );

    \I__583\ : Odrv4
    port map (
            O => \N__3491\,
            I => \uart.stateZ0Z_4\
        );

    \I__582\ : LocalMux
    port map (
            O => \N__3488\,
            I => \uart.stateZ0Z_4\
        );

    \I__581\ : LocalMux
    port map (
            O => \N__3483\,
            I => \uart.stateZ0Z_4\
        );

    \I__580\ : LocalMux
    port map (
            O => \N__3480\,
            I => \uart.stateZ0Z_4\
        );

    \I__579\ : CascadeMux
    port map (
            O => \N__3467\,
            I => \uart_frame_decoder.N_43_cascade_\
        );

    \I__578\ : CascadeMux
    port map (
            O => \N__3464\,
            I => \uart_frame_decoder.state_1_ns_i_i_a2_1_1_0_cascade_\
        );

    \I__577\ : CascadeMux
    port map (
            O => \N__3461\,
            I => \uart_frame_decoder.N_81_cascade_\
        );

    \I__576\ : CascadeMux
    port map (
            O => \N__3458\,
            I => \uart_frame_decoder.state_1_ns_0_i_a2_0_0_1Z0Z_2_cascade_\
        );

    \I__575\ : SRMux
    port map (
            O => \N__3455\,
            I => \N__3450\
        );

    \I__574\ : SRMux
    port map (
            O => \N__3454\,
            I => \N__3447\
        );

    \I__573\ : SRMux
    port map (
            O => \N__3453\,
            I => \N__3444\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__3450\,
            I => \N__3439\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__3447\,
            I => \N__3439\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__3444\,
            I => \N__3436\
        );

    \I__569\ : Span4Mux_v
    port map (
            O => \N__3439\,
            I => \N__3433\
        );

    \I__568\ : Span4Mux_h
    port map (
            O => \N__3436\,
            I => \N__3430\
        );

    \I__567\ : Span4Mux_h
    port map (
            O => \N__3433\,
            I => \N__3427\
        );

    \I__566\ : Odrv4
    port map (
            O => \N__3430\,
            I => \uart.state_RNIAFHLZ0Z_4\
        );

    \I__565\ : Odrv4
    port map (
            O => \N__3427\,
            I => \uart.state_RNIAFHLZ0Z_4\
        );

    \I__564\ : InMux
    port map (
            O => \N__3422\,
            I => \N__3417\
        );

    \I__563\ : InMux
    port map (
            O => \N__3421\,
            I => \N__3412\
        );

    \I__562\ : InMux
    port map (
            O => \N__3420\,
            I => \N__3412\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__3417\,
            I => \uart.stateZ0Z_1\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__3412\,
            I => \uart.stateZ0Z_1\
        );

    \I__559\ : CascadeMux
    port map (
            O => \N__3407\,
            I => \uart.N_151_cascade_\
        );

    \I__558\ : CascadeMux
    port map (
            O => \N__3404\,
            I => \N__3400\
        );

    \I__557\ : InMux
    port map (
            O => \N__3403\,
            I => \N__3397\
        );

    \I__556\ : InMux
    port map (
            O => \N__3400\,
            I => \N__3393\
        );

    \I__555\ : LocalMux
    port map (
            O => \N__3397\,
            I => \N__3389\
        );

    \I__554\ : InMux
    port map (
            O => \N__3396\,
            I => \N__3386\
        );

    \I__553\ : LocalMux
    port map (
            O => \N__3393\,
            I => \N__3383\
        );

    \I__552\ : InMux
    port map (
            O => \N__3392\,
            I => \N__3380\
        );

    \I__551\ : Odrv12
    port map (
            O => \N__3389\,
            I => \uart.stateZ0Z_2\
        );

    \I__550\ : LocalMux
    port map (
            O => \N__3386\,
            I => \uart.stateZ0Z_2\
        );

    \I__549\ : Odrv4
    port map (
            O => \N__3383\,
            I => \uart.stateZ0Z_2\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__3380\,
            I => \uart.stateZ0Z_2\
        );

    \I__547\ : InMux
    port map (
            O => \N__3371\,
            I => \N__3366\
        );

    \I__546\ : CascadeMux
    port map (
            O => \N__3370\,
            I => \N__3363\
        );

    \I__545\ : CascadeMux
    port map (
            O => \N__3369\,
            I => \N__3357\
        );

    \I__544\ : LocalMux
    port map (
            O => \N__3366\,
            I => \N__3353\
        );

    \I__543\ : InMux
    port map (
            O => \N__3363\,
            I => \N__3349\
        );

    \I__542\ : InMux
    port map (
            O => \N__3362\,
            I => \N__3346\
        );

    \I__541\ : InMux
    port map (
            O => \N__3361\,
            I => \N__3343\
        );

    \I__540\ : InMux
    port map (
            O => \N__3360\,
            I => \N__3338\
        );

    \I__539\ : InMux
    port map (
            O => \N__3357\,
            I => \N__3338\
        );

    \I__538\ : InMux
    port map (
            O => \N__3356\,
            I => \N__3335\
        );

    \I__537\ : Span4Mux_h
    port map (
            O => \N__3353\,
            I => \N__3331\
        );

    \I__536\ : InMux
    port map (
            O => \N__3352\,
            I => \N__3328\
        );

    \I__535\ : LocalMux
    port map (
            O => \N__3349\,
            I => \N__3317\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__3346\,
            I => \N__3317\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__3343\,
            I => \N__3317\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__3338\,
            I => \N__3317\
        );

    \I__531\ : LocalMux
    port map (
            O => \N__3335\,
            I => \N__3317\
        );

    \I__530\ : InMux
    port map (
            O => \N__3334\,
            I => \N__3314\
        );

    \I__529\ : Odrv4
    port map (
            O => \N__3331\,
            I => \uart.stateZ0Z_3\
        );

    \I__528\ : LocalMux
    port map (
            O => \N__3328\,
            I => \uart.stateZ0Z_3\
        );

    \I__527\ : Odrv4
    port map (
            O => \N__3317\,
            I => \uart.stateZ0Z_3\
        );

    \I__526\ : LocalMux
    port map (
            O => \N__3314\,
            I => \uart.stateZ0Z_3\
        );

    \I__525\ : InMux
    port map (
            O => \N__3305\,
            I => \N__3302\
        );

    \I__524\ : LocalMux
    port map (
            O => \N__3302\,
            I => \N__3299\
        );

    \I__523\ : Span4Mux_s1_v
    port map (
            O => \N__3299\,
            I => \N__3296\
        );

    \I__522\ : Odrv4
    port map (
            O => \N__3296\,
            I => \uart.state_srsts_i_1_1_3\
        );

    \I__521\ : CascadeMux
    port map (
            O => \N__3293\,
            I => \uart.N_166_cascade_\
        );

    \I__520\ : CascadeMux
    port map (
            O => \N__3290\,
            I => \uart.state_srsts_0_1_0_cascade_\
        );

    \I__519\ : InMux
    port map (
            O => \N__3287\,
            I => \N__3284\
        );

    \I__518\ : LocalMux
    port map (
            O => \N__3284\,
            I => \N__3280\
        );

    \I__517\ : InMux
    port map (
            O => \N__3283\,
            I => \N__3277\
        );

    \I__516\ : Odrv4
    port map (
            O => \N__3280\,
            I => \uart.stateZ0Z_0\
        );

    \I__515\ : LocalMux
    port map (
            O => \N__3277\,
            I => \uart.stateZ0Z_0\
        );

    \I__514\ : CascadeMux
    port map (
            O => \N__3272\,
            I => \N__3269\
        );

    \I__513\ : InMux
    port map (
            O => \N__3269\,
            I => \N__3266\
        );

    \I__512\ : LocalMux
    port map (
            O => \N__3266\,
            I => \N__3263\
        );

    \I__511\ : Odrv4
    port map (
            O => \N__3263\,
            I => \uart_frame_decoder.N_43\
        );

    \I__510\ : InMux
    port map (
            O => \N__3260\,
            I => \N__3256\
        );

    \I__509\ : CascadeMux
    port map (
            O => \N__3259\,
            I => \N__3253\
        );

    \I__508\ : LocalMux
    port map (
            O => \N__3256\,
            I => \N__3250\
        );

    \I__507\ : InMux
    port map (
            O => \N__3253\,
            I => \N__3247\
        );

    \I__506\ : Odrv4
    port map (
            O => \N__3250\,
            I => \uart.data_AuxZ0Z_7\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__3247\,
            I => \uart.data_AuxZ0Z_7\
        );

    \I__504\ : CascadeMux
    port map (
            O => \N__3242\,
            I => \uart.timer_Count10lto5_0_0_cascade_\
        );

    \I__503\ : InMux
    port map (
            O => \N__3239\,
            I => \N__3234\
        );

    \I__502\ : InMux
    port map (
            O => \N__3238\,
            I => \N__3231\
        );

    \I__501\ : InMux
    port map (
            O => \N__3237\,
            I => \N__3228\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__3234\,
            I => \uart.N_177\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__3231\,
            I => \uart.N_177\
        );

    \I__498\ : LocalMux
    port map (
            O => \N__3228\,
            I => \uart.N_177\
        );

    \I__497\ : CascadeMux
    port map (
            O => \N__3221\,
            I => \uart.N_168_cascade_\
        );

    \I__496\ : InMux
    port map (
            O => \N__3218\,
            I => \N__3214\
        );

    \I__495\ : InMux
    port map (
            O => \N__3217\,
            I => \N__3211\
        );

    \I__494\ : LocalMux
    port map (
            O => \N__3214\,
            I => \reset_module_System.countZ0Z_14\
        );

    \I__493\ : LocalMux
    port map (
            O => \N__3211\,
            I => \reset_module_System.countZ0Z_14\
        );

    \I__492\ : InMux
    port map (
            O => \N__3206\,
            I => \N__3202\
        );

    \I__491\ : InMux
    port map (
            O => \N__3205\,
            I => \N__3199\
        );

    \I__490\ : LocalMux
    port map (
            O => \N__3202\,
            I => \reset_module_System.countZ0Z_17\
        );

    \I__489\ : LocalMux
    port map (
            O => \N__3199\,
            I => \reset_module_System.countZ0Z_17\
        );

    \I__488\ : CascadeMux
    port map (
            O => \N__3194\,
            I => \reset_module_System.reset6_3_cascade_\
        );

    \I__487\ : InMux
    port map (
            O => \N__3191\,
            I => \N__3188\
        );

    \I__486\ : LocalMux
    port map (
            O => \N__3188\,
            I => \reset_module_System.reset6_13\
        );

    \I__485\ : InMux
    port map (
            O => \N__3185\,
            I => \N__3181\
        );

    \I__484\ : InMux
    port map (
            O => \N__3184\,
            I => \N__3178\
        );

    \I__483\ : LocalMux
    port map (
            O => \N__3181\,
            I => \reset_module_System.countZ0Z_12\
        );

    \I__482\ : LocalMux
    port map (
            O => \N__3178\,
            I => \reset_module_System.countZ0Z_12\
        );

    \I__481\ : InMux
    port map (
            O => \N__3173\,
            I => \N__3167\
        );

    \I__480\ : CascadeMux
    port map (
            O => \N__3172\,
            I => \N__3164\
        );

    \I__479\ : InMux
    port map (
            O => \N__3171\,
            I => \N__3161\
        );

    \I__478\ : InMux
    port map (
            O => \N__3170\,
            I => \N__3158\
        );

    \I__477\ : LocalMux
    port map (
            O => \N__3167\,
            I => \N__3155\
        );

    \I__476\ : InMux
    port map (
            O => \N__3164\,
            I => \N__3152\
        );

    \I__475\ : LocalMux
    port map (
            O => \N__3161\,
            I => \reset_module_System.countZ0Z_0\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__3158\,
            I => \reset_module_System.countZ0Z_0\
        );

    \I__473\ : Odrv12
    port map (
            O => \N__3155\,
            I => \reset_module_System.countZ0Z_0\
        );

    \I__472\ : LocalMux
    port map (
            O => \N__3152\,
            I => \reset_module_System.countZ0Z_0\
        );

    \I__471\ : CascadeMux
    port map (
            O => \N__3143\,
            I => \reset_module_System.reset6_17_cascade_\
        );

    \I__470\ : InMux
    port map (
            O => \N__3140\,
            I => \N__3137\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__3137\,
            I => \reset_module_System.reset6_11\
        );

    \I__468\ : InMux
    port map (
            O => \N__3134\,
            I => \N__3119\
        );

    \I__467\ : InMux
    port map (
            O => \N__3133\,
            I => \N__3119\
        );

    \I__466\ : InMux
    port map (
            O => \N__3132\,
            I => \N__3119\
        );

    \I__465\ : InMux
    port map (
            O => \N__3131\,
            I => \N__3119\
        );

    \I__464\ : InMux
    port map (
            O => \N__3130\,
            I => \N__3119\
        );

    \I__463\ : LocalMux
    port map (
            O => \N__3119\,
            I => \reset_module_System.reset6_19\
        );

    \I__462\ : CascadeMux
    port map (
            O => \N__3116\,
            I => \uart.N_169_cascade_\
        );

    \I__461\ : CascadeMux
    port map (
            O => \N__3113\,
            I => \uart.state_srsts_i_1_3_cascade_\
        );

    \I__460\ : InMux
    port map (
            O => \N__3110\,
            I => \N__3106\
        );

    \I__459\ : InMux
    port map (
            O => \N__3109\,
            I => \N__3103\
        );

    \I__458\ : LocalMux
    port map (
            O => \N__3106\,
            I => \uart.data_AuxZ0Z_0\
        );

    \I__457\ : LocalMux
    port map (
            O => \N__3103\,
            I => \uart.data_AuxZ0Z_0\
        );

    \I__456\ : InMux
    port map (
            O => \N__3098\,
            I => \N__3094\
        );

    \I__455\ : CascadeMux
    port map (
            O => \N__3097\,
            I => \N__3091\
        );

    \I__454\ : LocalMux
    port map (
            O => \N__3094\,
            I => \N__3088\
        );

    \I__453\ : InMux
    port map (
            O => \N__3091\,
            I => \N__3085\
        );

    \I__452\ : Odrv4
    port map (
            O => \N__3088\,
            I => \uart.data_AuxZ0Z_2\
        );

    \I__451\ : LocalMux
    port map (
            O => \N__3085\,
            I => \uart.data_AuxZ0Z_2\
        );

    \I__450\ : InMux
    port map (
            O => \N__3080\,
            I => \N__3076\
        );

    \I__449\ : InMux
    port map (
            O => \N__3079\,
            I => \N__3073\
        );

    \I__448\ : LocalMux
    port map (
            O => \N__3076\,
            I => \N__3070\
        );

    \I__447\ : LocalMux
    port map (
            O => \N__3073\,
            I => \uart.data_AuxZ0Z_3\
        );

    \I__446\ : Odrv4
    port map (
            O => \N__3070\,
            I => \uart.data_AuxZ0Z_3\
        );

    \I__445\ : InMux
    port map (
            O => \N__3065\,
            I => \N__3062\
        );

    \I__444\ : LocalMux
    port map (
            O => \N__3062\,
            I => \N__3058\
        );

    \I__443\ : InMux
    port map (
            O => \N__3061\,
            I => \N__3055\
        );

    \I__442\ : Odrv4
    port map (
            O => \N__3058\,
            I => \uart.data_AuxZ0Z_5\
        );

    \I__441\ : LocalMux
    port map (
            O => \N__3055\,
            I => \uart.data_AuxZ0Z_5\
        );

    \I__440\ : InMux
    port map (
            O => \N__3050\,
            I => \N__3047\
        );

    \I__439\ : LocalMux
    port map (
            O => \N__3047\,
            I => \N__3043\
        );

    \I__438\ : InMux
    port map (
            O => \N__3046\,
            I => \N__3040\
        );

    \I__437\ : Odrv4
    port map (
            O => \N__3043\,
            I => \reset_module_System.countZ0Z_16\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__3040\,
            I => \reset_module_System.countZ0Z_16\
        );

    \I__435\ : InMux
    port map (
            O => \N__3035\,
            I => \N__3031\
        );

    \I__434\ : InMux
    port map (
            O => \N__3034\,
            I => \N__3028\
        );

    \I__433\ : LocalMux
    port map (
            O => \N__3031\,
            I => \reset_module_System.countZ0Z_4\
        );

    \I__432\ : LocalMux
    port map (
            O => \N__3028\,
            I => \reset_module_System.countZ0Z_4\
        );

    \I__431\ : CascadeMux
    port map (
            O => \N__3023\,
            I => \N__3020\
        );

    \I__430\ : InMux
    port map (
            O => \N__3020\,
            I => \N__3016\
        );

    \I__429\ : InMux
    port map (
            O => \N__3019\,
            I => \N__3013\
        );

    \I__428\ : LocalMux
    port map (
            O => \N__3016\,
            I => \N__3010\
        );

    \I__427\ : LocalMux
    port map (
            O => \N__3013\,
            I => \reset_module_System.countZ0Z_18\
        );

    \I__426\ : Odrv4
    port map (
            O => \N__3010\,
            I => \reset_module_System.countZ0Z_18\
        );

    \I__425\ : CascadeMux
    port map (
            O => \N__3005\,
            I => \reset_module_System.reset6_14_cascade_\
        );

    \I__424\ : InMux
    port map (
            O => \N__3002\,
            I => \N__2998\
        );

    \I__423\ : InMux
    port map (
            O => \N__3001\,
            I => \N__2995\
        );

    \I__422\ : LocalMux
    port map (
            O => \N__2998\,
            I => \reset_module_System.countZ0Z_6\
        );

    \I__421\ : LocalMux
    port map (
            O => \N__2995\,
            I => \reset_module_System.countZ0Z_6\
        );

    \I__420\ : InMux
    port map (
            O => \N__2990\,
            I => \N__2986\
        );

    \I__419\ : InMux
    port map (
            O => \N__2989\,
            I => \N__2983\
        );

    \I__418\ : LocalMux
    port map (
            O => \N__2986\,
            I => \reset_module_System.countZ0Z_3\
        );

    \I__417\ : LocalMux
    port map (
            O => \N__2983\,
            I => \reset_module_System.countZ0Z_3\
        );

    \I__416\ : CascadeMux
    port map (
            O => \N__2978\,
            I => \N__2975\
        );

    \I__415\ : InMux
    port map (
            O => \N__2975\,
            I => \N__2971\
        );

    \I__414\ : InMux
    port map (
            O => \N__2974\,
            I => \N__2968\
        );

    \I__413\ : LocalMux
    port map (
            O => \N__2971\,
            I => \N__2965\
        );

    \I__412\ : LocalMux
    port map (
            O => \N__2968\,
            I => \reset_module_System.countZ0Z_20\
        );

    \I__411\ : Odrv4
    port map (
            O => \N__2965\,
            I => \reset_module_System.countZ0Z_20\
        );

    \I__410\ : InMux
    port map (
            O => \N__2960\,
            I => \N__2956\
        );

    \I__409\ : InMux
    port map (
            O => \N__2959\,
            I => \N__2953\
        );

    \I__408\ : LocalMux
    port map (
            O => \N__2956\,
            I => \reset_module_System.countZ0Z_8\
        );

    \I__407\ : LocalMux
    port map (
            O => \N__2953\,
            I => \reset_module_System.countZ0Z_8\
        );

    \I__406\ : InMux
    port map (
            O => \N__2948\,
            I => \N__2944\
        );

    \I__405\ : InMux
    port map (
            O => \N__2947\,
            I => \N__2941\
        );

    \I__404\ : LocalMux
    port map (
            O => \N__2944\,
            I => \reset_module_System.countZ0Z_7\
        );

    \I__403\ : LocalMux
    port map (
            O => \N__2941\,
            I => \reset_module_System.countZ0Z_7\
        );

    \I__402\ : CascadeMux
    port map (
            O => \N__2936\,
            I => \N__2932\
        );

    \I__401\ : InMux
    port map (
            O => \N__2935\,
            I => \N__2929\
        );

    \I__400\ : InMux
    port map (
            O => \N__2932\,
            I => \N__2926\
        );

    \I__399\ : LocalMux
    port map (
            O => \N__2929\,
            I => \reset_module_System.countZ0Z_9\
        );

    \I__398\ : LocalMux
    port map (
            O => \N__2926\,
            I => \reset_module_System.countZ0Z_9\
        );

    \I__397\ : InMux
    port map (
            O => \N__2921\,
            I => \N__2917\
        );

    \I__396\ : InMux
    port map (
            O => \N__2920\,
            I => \N__2914\
        );

    \I__395\ : LocalMux
    port map (
            O => \N__2917\,
            I => \reset_module_System.countZ0Z_5\
        );

    \I__394\ : LocalMux
    port map (
            O => \N__2914\,
            I => \reset_module_System.countZ0Z_5\
        );

    \I__393\ : InMux
    port map (
            O => \N__2909\,
            I => \N__2906\
        );

    \I__392\ : LocalMux
    port map (
            O => \N__2906\,
            I => \N__2903\
        );

    \I__391\ : Span4Mux_h
    port map (
            O => \N__2903\,
            I => \N__2900\
        );

    \I__390\ : Odrv4
    port map (
            O => \N__2900\,
            I => \reset_module_System.count_1_1\
        );

    \I__389\ : InMux
    port map (
            O => \N__2897\,
            I => \N__2894\
        );

    \I__388\ : LocalMux
    port map (
            O => \N__2894\,
            I => \N__2889\
        );

    \I__387\ : InMux
    port map (
            O => \N__2893\,
            I => \N__2886\
        );

    \I__386\ : InMux
    port map (
            O => \N__2892\,
            I => \N__2883\
        );

    \I__385\ : Odrv12
    port map (
            O => \N__2889\,
            I => \reset_module_System.countZ0Z_1\
        );

    \I__384\ : LocalMux
    port map (
            O => \N__2886\,
            I => \reset_module_System.countZ0Z_1\
        );

    \I__383\ : LocalMux
    port map (
            O => \N__2883\,
            I => \reset_module_System.countZ0Z_1\
        );

    \I__382\ : CascadeMux
    port map (
            O => \N__2876\,
            I => \N__2872\
        );

    \I__381\ : CascadeMux
    port map (
            O => \N__2875\,
            I => \N__2869\
        );

    \I__380\ : InMux
    port map (
            O => \N__2872\,
            I => \N__2855\
        );

    \I__379\ : InMux
    port map (
            O => \N__2869\,
            I => \N__2855\
        );

    \I__378\ : InMux
    port map (
            O => \N__2868\,
            I => \N__2855\
        );

    \I__377\ : InMux
    port map (
            O => \N__2867\,
            I => \N__2855\
        );

    \I__376\ : InMux
    port map (
            O => \N__2866\,
            I => \N__2855\
        );

    \I__375\ : LocalMux
    port map (
            O => \N__2855\,
            I => \N__2852\
        );

    \I__374\ : Span4Mux_h
    port map (
            O => \N__2852\,
            I => \N__2849\
        );

    \I__373\ : Odrv4
    port map (
            O => \N__2849\,
            I => \reset_module_System.reset6_15\
        );

    \I__372\ : CascadeMux
    port map (
            O => \N__2846\,
            I => \N__2843\
        );

    \I__371\ : InMux
    port map (
            O => \N__2843\,
            I => \N__2831\
        );

    \I__370\ : InMux
    port map (
            O => \N__2842\,
            I => \N__2831\
        );

    \I__369\ : InMux
    port map (
            O => \N__2841\,
            I => \N__2831\
        );

    \I__368\ : InMux
    port map (
            O => \N__2840\,
            I => \N__2831\
        );

    \I__367\ : LocalMux
    port map (
            O => \N__2831\,
            I => \reset_module_System.reset6_14\
        );

    \I__366\ : InMux
    port map (
            O => \N__2828\,
            I => \N__2825\
        );

    \I__365\ : LocalMux
    port map (
            O => \N__2825\,
            I => \reset_module_System.count_1_2\
        );

    \I__364\ : CascadeMux
    port map (
            O => \N__2822\,
            I => \N__2819\
        );

    \I__363\ : InMux
    port map (
            O => \N__2819\,
            I => \N__2815\
        );

    \I__362\ : InMux
    port map (
            O => \N__2818\,
            I => \N__2812\
        );

    \I__361\ : LocalMux
    port map (
            O => \N__2815\,
            I => \reset_module_System.countZ0Z_2\
        );

    \I__360\ : LocalMux
    port map (
            O => \N__2812\,
            I => \reset_module_System.countZ0Z_2\
        );

    \I__359\ : InMux
    port map (
            O => \N__2807\,
            I => \N__2803\
        );

    \I__358\ : InMux
    port map (
            O => \N__2806\,
            I => \N__2800\
        );

    \I__357\ : LocalMux
    port map (
            O => \N__2803\,
            I => \reset_module_System.countZ0Z_11\
        );

    \I__356\ : LocalMux
    port map (
            O => \N__2800\,
            I => \reset_module_System.countZ0Z_11\
        );

    \I__355\ : InMux
    port map (
            O => \N__2795\,
            I => \N__2791\
        );

    \I__354\ : InMux
    port map (
            O => \N__2794\,
            I => \N__2788\
        );

    \I__353\ : LocalMux
    port map (
            O => \N__2791\,
            I => \reset_module_System.countZ0Z_10\
        );

    \I__352\ : LocalMux
    port map (
            O => \N__2788\,
            I => \reset_module_System.countZ0Z_10\
        );

    \I__351\ : CascadeMux
    port map (
            O => \N__2783\,
            I => \N__2778\
        );

    \I__350\ : InMux
    port map (
            O => \N__2782\,
            I => \N__2771\
        );

    \I__349\ : InMux
    port map (
            O => \N__2781\,
            I => \N__2764\
        );

    \I__348\ : InMux
    port map (
            O => \N__2778\,
            I => \N__2764\
        );

    \I__347\ : InMux
    port map (
            O => \N__2777\,
            I => \N__2764\
        );

    \I__346\ : InMux
    port map (
            O => \N__2776\,
            I => \N__2757\
        );

    \I__345\ : InMux
    port map (
            O => \N__2775\,
            I => \N__2757\
        );

    \I__344\ : InMux
    port map (
            O => \N__2774\,
            I => \N__2757\
        );

    \I__343\ : LocalMux
    port map (
            O => \N__2771\,
            I => \uart.un1_state_2_0\
        );

    \I__342\ : LocalMux
    port map (
            O => \N__2764\,
            I => \uart.un1_state_2_0\
        );

    \I__341\ : LocalMux
    port map (
            O => \N__2757\,
            I => \uart.un1_state_2_0\
        );

    \I__340\ : InMux
    port map (
            O => \N__2750\,
            I => \N__2747\
        );

    \I__339\ : LocalMux
    port map (
            O => \N__2747\,
            I => \uart.data_Auxce_0_0_4\
        );

    \I__338\ : InMux
    port map (
            O => \N__2744\,
            I => \N__2741\
        );

    \I__337\ : LocalMux
    port map (
            O => \N__2741\,
            I => \uart.data_Auxce_0_0_0\
        );

    \I__336\ : InMux
    port map (
            O => \N__2738\,
            I => \N__2735\
        );

    \I__335\ : LocalMux
    port map (
            O => \N__2735\,
            I => \uart.data_Auxce_0_1\
        );

    \I__334\ : InMux
    port map (
            O => \N__2732\,
            I => \N__2729\
        );

    \I__333\ : LocalMux
    port map (
            O => \N__2729\,
            I => \N__2726\
        );

    \I__332\ : Odrv4
    port map (
            O => \N__2726\,
            I => \uart.data_Auxce_0_0_2\
        );

    \I__331\ : InMux
    port map (
            O => \N__2723\,
            I => \N__2714\
        );

    \I__330\ : InMux
    port map (
            O => \N__2722\,
            I => \N__2714\
        );

    \I__329\ : InMux
    port map (
            O => \N__2721\,
            I => \N__2714\
        );

    \I__328\ : LocalMux
    port map (
            O => \N__2714\,
            I => \uart.un1_state_5_0\
        );

    \I__327\ : CascadeMux
    port map (
            O => \N__2711\,
            I => \N__2701\
        );

    \I__326\ : CascadeMux
    port map (
            O => \N__2710\,
            I => \N__2698\
        );

    \I__325\ : InMux
    port map (
            O => \N__2709\,
            I => \N__2693\
        );

    \I__324\ : InMux
    port map (
            O => \N__2708\,
            I => \N__2682\
        );

    \I__323\ : InMux
    port map (
            O => \N__2707\,
            I => \N__2682\
        );

    \I__322\ : InMux
    port map (
            O => \N__2706\,
            I => \N__2682\
        );

    \I__321\ : InMux
    port map (
            O => \N__2705\,
            I => \N__2682\
        );

    \I__320\ : InMux
    port map (
            O => \N__2704\,
            I => \N__2682\
        );

    \I__319\ : InMux
    port map (
            O => \N__2701\,
            I => \N__2677\
        );

    \I__318\ : InMux
    port map (
            O => \N__2698\,
            I => \N__2677\
        );

    \I__317\ : InMux
    port map (
            O => \N__2697\,
            I => \N__2672\
        );

    \I__316\ : InMux
    port map (
            O => \N__2696\,
            I => \N__2672\
        );

    \I__315\ : LocalMux
    port map (
            O => \N__2693\,
            I => \uart.bit_CountZ0Z_2\
        );

    \I__314\ : LocalMux
    port map (
            O => \N__2682\,
            I => \uart.bit_CountZ0Z_2\
        );

    \I__313\ : LocalMux
    port map (
            O => \N__2677\,
            I => \uart.bit_CountZ0Z_2\
        );

    \I__312\ : LocalMux
    port map (
            O => \N__2672\,
            I => \uart.bit_CountZ0Z_2\
        );

    \I__311\ : CascadeMux
    port map (
            O => \N__2663\,
            I => \N__2658\
        );

    \I__310\ : CascadeMux
    port map (
            O => \N__2662\,
            I => \N__2653\
        );

    \I__309\ : CascadeMux
    port map (
            O => \N__2661\,
            I => \N__2645\
        );

    \I__308\ : InMux
    port map (
            O => \N__2658\,
            I => \N__2633\
        );

    \I__307\ : InMux
    port map (
            O => \N__2657\,
            I => \N__2633\
        );

    \I__306\ : InMux
    port map (
            O => \N__2656\,
            I => \N__2633\
        );

    \I__305\ : InMux
    port map (
            O => \N__2653\,
            I => \N__2633\
        );

    \I__304\ : InMux
    port map (
            O => \N__2652\,
            I => \N__2633\
        );

    \I__303\ : InMux
    port map (
            O => \N__2651\,
            I => \N__2628\
        );

    \I__302\ : InMux
    port map (
            O => \N__2650\,
            I => \N__2628\
        );

    \I__301\ : InMux
    port map (
            O => \N__2649\,
            I => \N__2623\
        );

    \I__300\ : InMux
    port map (
            O => \N__2648\,
            I => \N__2623\
        );

    \I__299\ : InMux
    port map (
            O => \N__2645\,
            I => \N__2618\
        );

    \I__298\ : InMux
    port map (
            O => \N__2644\,
            I => \N__2618\
        );

    \I__297\ : LocalMux
    port map (
            O => \N__2633\,
            I => \uart.bit_CountZ0Z_1\
        );

    \I__296\ : LocalMux
    port map (
            O => \N__2628\,
            I => \uart.bit_CountZ0Z_1\
        );

    \I__295\ : LocalMux
    port map (
            O => \N__2623\,
            I => \uart.bit_CountZ0Z_1\
        );

    \I__294\ : LocalMux
    port map (
            O => \N__2618\,
            I => \uart.bit_CountZ0Z_1\
        );

    \I__293\ : InMux
    port map (
            O => \N__2609\,
            I => \N__2587\
        );

    \I__292\ : InMux
    port map (
            O => \N__2608\,
            I => \N__2587\
        );

    \I__291\ : InMux
    port map (
            O => \N__2607\,
            I => \N__2587\
        );

    \I__290\ : InMux
    port map (
            O => \N__2606\,
            I => \N__2587\
        );

    \I__289\ : InMux
    port map (
            O => \N__2605\,
            I => \N__2587\
        );

    \I__288\ : InMux
    port map (
            O => \N__2604\,
            I => \N__2582\
        );

    \I__287\ : InMux
    port map (
            O => \N__2603\,
            I => \N__2582\
        );

    \I__286\ : InMux
    port map (
            O => \N__2602\,
            I => \N__2575\
        );

    \I__285\ : InMux
    port map (
            O => \N__2601\,
            I => \N__2575\
        );

    \I__284\ : InMux
    port map (
            O => \N__2600\,
            I => \N__2575\
        );

    \I__283\ : InMux
    port map (
            O => \N__2599\,
            I => \N__2570\
        );

    \I__282\ : InMux
    port map (
            O => \N__2598\,
            I => \N__2570\
        );

    \I__281\ : LocalMux
    port map (
            O => \N__2587\,
            I => \uart.bit_CountZ0Z_0\
        );

    \I__280\ : LocalMux
    port map (
            O => \N__2582\,
            I => \uart.bit_CountZ0Z_0\
        );

    \I__279\ : LocalMux
    port map (
            O => \N__2575\,
            I => \uart.bit_CountZ0Z_0\
        );

    \I__278\ : LocalMux
    port map (
            O => \N__2570\,
            I => \uart.bit_CountZ0Z_0\
        );

    \I__277\ : CascadeMux
    port map (
            O => \N__2561\,
            I => \N__2558\
        );

    \I__276\ : InMux
    port map (
            O => \N__2558\,
            I => \N__2555\
        );

    \I__275\ : LocalMux
    port map (
            O => \N__2555\,
            I => \uart.data_Auxce_0_3\
        );

    \I__274\ : InMux
    port map (
            O => \N__2552\,
            I => \reset_module_System.count_1_cry_18\
        );

    \I__273\ : InMux
    port map (
            O => \N__2549\,
            I => \reset_module_System.count_1_cry_19\
        );

    \I__272\ : InMux
    port map (
            O => \N__2546\,
            I => \reset_module_System.count_1_cry_20\
        );

    \I__271\ : CascadeMux
    port map (
            O => \N__2543\,
            I => \N__2539\
        );

    \I__270\ : InMux
    port map (
            O => \N__2542\,
            I => \N__2536\
        );

    \I__269\ : InMux
    port map (
            O => \N__2539\,
            I => \N__2533\
        );

    \I__268\ : LocalMux
    port map (
            O => \N__2536\,
            I => \reset_module_System.countZ0Z_21\
        );

    \I__267\ : LocalMux
    port map (
            O => \N__2533\,
            I => \reset_module_System.countZ0Z_21\
        );

    \I__266\ : InMux
    port map (
            O => \N__2528\,
            I => \N__2525\
        );

    \I__265\ : LocalMux
    port map (
            O => \N__2525\,
            I => \uart.data_Auxce_0_5\
        );

    \I__264\ : InMux
    port map (
            O => \N__2522\,
            I => \N__2519\
        );

    \I__263\ : LocalMux
    port map (
            O => \N__2519\,
            I => \N__2516\
        );

    \I__262\ : Odrv4
    port map (
            O => \N__2516\,
            I => \uart.timer_Count_RNI9M0NZ0Z_1\
        );

    \I__261\ : CascadeMux
    port map (
            O => \N__2513\,
            I => \uart.timer_Count_RNILKMA1Z0Z_0_cascade_\
        );

    \I__260\ : CascadeMux
    port map (
            O => \N__2510\,
            I => \uart.un1_state_2_0_cascade_\
        );

    \I__259\ : InMux
    port map (
            O => \N__2507\,
            I => \reset_module_System.count_1_cry_10\
        );

    \I__258\ : InMux
    port map (
            O => \N__2504\,
            I => \reset_module_System.count_1_cry_11\
        );

    \I__257\ : InMux
    port map (
            O => \N__2501\,
            I => \N__2497\
        );

    \I__256\ : InMux
    port map (
            O => \N__2500\,
            I => \N__2494\
        );

    \I__255\ : LocalMux
    port map (
            O => \N__2497\,
            I => \reset_module_System.countZ0Z_13\
        );

    \I__254\ : LocalMux
    port map (
            O => \N__2494\,
            I => \reset_module_System.countZ0Z_13\
        );

    \I__253\ : InMux
    port map (
            O => \N__2489\,
            I => \reset_module_System.count_1_cry_12\
        );

    \I__252\ : InMux
    port map (
            O => \N__2486\,
            I => \reset_module_System.count_1_cry_13\
        );

    \I__251\ : InMux
    port map (
            O => \N__2483\,
            I => \N__2479\
        );

    \I__250\ : InMux
    port map (
            O => \N__2482\,
            I => \N__2476\
        );

    \I__249\ : LocalMux
    port map (
            O => \N__2479\,
            I => \reset_module_System.countZ0Z_15\
        );

    \I__248\ : LocalMux
    port map (
            O => \N__2476\,
            I => \reset_module_System.countZ0Z_15\
        );

    \I__247\ : InMux
    port map (
            O => \N__2471\,
            I => \reset_module_System.count_1_cry_14\
        );

    \I__246\ : InMux
    port map (
            O => \N__2468\,
            I => \reset_module_System.count_1_cry_15\
        );

    \I__245\ : InMux
    port map (
            O => \N__2465\,
            I => \bfn_8_3_0_\
        );

    \I__244\ : InMux
    port map (
            O => \N__2462\,
            I => \reset_module_System.count_1_cry_17\
        );

    \I__243\ : InMux
    port map (
            O => \N__2459\,
            I => \N__2455\
        );

    \I__242\ : InMux
    port map (
            O => \N__2458\,
            I => \N__2452\
        );

    \I__241\ : LocalMux
    port map (
            O => \N__2455\,
            I => \reset_module_System.countZ0Z_19\
        );

    \I__240\ : LocalMux
    port map (
            O => \N__2452\,
            I => \reset_module_System.countZ0Z_19\
        );

    \I__239\ : InMux
    port map (
            O => \N__2447\,
            I => \reset_module_System.count_1_cry_1\
        );

    \I__238\ : InMux
    port map (
            O => \N__2444\,
            I => \reset_module_System.count_1_cry_2\
        );

    \I__237\ : InMux
    port map (
            O => \N__2441\,
            I => \reset_module_System.count_1_cry_3\
        );

    \I__236\ : InMux
    port map (
            O => \N__2438\,
            I => \reset_module_System.count_1_cry_4\
        );

    \I__235\ : InMux
    port map (
            O => \N__2435\,
            I => \reset_module_System.count_1_cry_5\
        );

    \I__234\ : InMux
    port map (
            O => \N__2432\,
            I => \reset_module_System.count_1_cry_6\
        );

    \I__233\ : InMux
    port map (
            O => \N__2429\,
            I => \reset_module_System.count_1_cry_7\
        );

    \I__232\ : InMux
    port map (
            O => \N__2426\,
            I => \bfn_8_2_0_\
        );

    \I__231\ : InMux
    port map (
            O => \N__2423\,
            I => \reset_module_System.count_1_cry_9\
        );

    \I__230\ : CascadeMux
    port map (
            O => \N__2420\,
            I => \uart.N_133_0_cascade_\
        );

    \I__229\ : InMux
    port map (
            O => \N__2417\,
            I => \N__2413\
        );

    \I__228\ : InMux
    port map (
            O => \N__2416\,
            I => \N__2410\
        );

    \I__227\ : LocalMux
    port map (
            O => \N__2413\,
            I => \uart.N_133_0\
        );

    \I__226\ : LocalMux
    port map (
            O => \N__2410\,
            I => \uart.N_133_0\
        );

    \I__225\ : CascadeMux
    port map (
            O => \N__2405\,
            I => \uart.data_Auxce_0_6_cascade_\
        );

    \I__224\ : InMux
    port map (
            O => \N__2402\,
            I => \N__2399\
        );

    \I__223\ : LocalMux
    port map (
            O => \N__2399\,
            I => \N__2396\
        );

    \I__222\ : Odrv4
    port map (
            O => \N__2396\,
            I => \uart.CO1_0\
        );

    \I__221\ : IoInMux
    port map (
            O => \N__2393\,
            I => \N__2390\
        );

    \I__220\ : LocalMux
    port map (
            O => \N__2390\,
            I => \N__2387\
        );

    \I__219\ : Span4Mux_s0_v
    port map (
            O => \N__2387\,
            I => \N__2384\
        );

    \I__218\ : Sp12to4
    port map (
            O => \N__2384\,
            I => \N__2380\
        );

    \I__217\ : CascadeMux
    port map (
            O => \N__2383\,
            I => \N__2377\
        );

    \I__216\ : Span12Mux_h
    port map (
            O => \N__2380\,
            I => \N__2374\
        );

    \I__215\ : InMux
    port map (
            O => \N__2377\,
            I => \N__2371\
        );

    \I__214\ : Odrv12
    port map (
            O => \N__2374\,
            I => frame_decoder_dv_c
        );

    \I__213\ : LocalMux
    port map (
            O => \N__2371\,
            I => frame_decoder_dv_c
        );

    \I__212\ : InMux
    port map (
            O => \N__2366\,
            I => \N__2362\
        );

    \I__211\ : IoInMux
    port map (
            O => \N__2365\,
            I => \N__2359\
        );

    \I__210\ : LocalMux
    port map (
            O => \N__2362\,
            I => \N__2356\
        );

    \I__209\ : LocalMux
    port map (
            O => \N__2359\,
            I => \N__2353\
        );

    \I__208\ : Span4Mux_h
    port map (
            O => \N__2356\,
            I => \N__2350\
        );

    \I__207\ : IoSpan4Mux
    port map (
            O => \N__2353\,
            I => \N__2347\
        );

    \I__206\ : Odrv4
    port map (
            O => \N__2350\,
            I => uart_input_c
        );

    \I__205\ : Odrv4
    port map (
            O => \N__2347\,
            I => uart_input_c
        );

    \I__204\ : InMux
    port map (
            O => \N__2342\,
            I => \N__2339\
        );

    \I__203\ : LocalMux
    port map (
            O => \N__2339\,
            I => \uart_sync.aux_0__0_Z0Z_0\
        );

    \I__202\ : InMux
    port map (
            O => \N__2336\,
            I => \N__2333\
        );

    \I__201\ : LocalMux
    port map (
            O => \N__2333\,
            I => \uart_sync.aux_1__0_Z0Z_0\
        );

    \I__200\ : InMux
    port map (
            O => \N__2330\,
            I => \N__2327\
        );

    \I__199\ : LocalMux
    port map (
            O => \N__2327\,
            I => \uart_sync.aux_2__0_Z0Z_0\
        );

    \I__198\ : InMux
    port map (
            O => \N__2324\,
            I => \N__2321\
        );

    \I__197\ : LocalMux
    port map (
            O => \N__2321\,
            I => \uart_sync.aux_3__0_Z0Z_0\
        );

    \IN_MUX_bfv_11_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_1_0_\
        );

    \IN_MUX_bfv_10_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_5_0_\
        );

    \IN_MUX_bfv_8_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_1_0_\
        );

    \IN_MUX_bfv_8_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \reset_module_System.count_1_cry_8\,
            carryinitout => \bfn_8_2_0_\
        );

    \IN_MUX_bfv_8_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \reset_module_System.count_1_cry_16\,
            carryinitout => \bfn_8_3_0_\
        );

    \IN_MUX_bfv_12_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_2_0_\
        );

    \IN_MUX_bfv_12_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \uart_frame_decoder.un1_WDT_cry_7\,
            carryinitout => \bfn_12_3_0_\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \reset_module_System.count_RNO_0_1_LC_5_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3173\,
            in2 => \_gnd_net_\,
            in3 => \N__2897\,
            lcout => \reset_module_System.count_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.source_data_valid_LC_7_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011001000"
        )
    port map (
            in0 => \N__5033\,
            in1 => \N__5501\,
            in2 => \N__2383\,
            in3 => \N__4106\,
            lcout => frame_decoder_dv_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4883\,
            ce => 'H',
            sr => \N__5551\
        );

    \uart_sync.aux_2__0__0_LC_7_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2336\,
            lcout => \uart_sync.aux_2__0_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4881\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_sync.aux_0__0__0_LC_7_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2366\,
            lcout => \uart_sync.aux_0__0_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4881\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_sync.Q_0__0_LC_7_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2324\,
            lcout => uart_input_sync,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4881\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_sync.aux_1__0__0_LC_7_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2342\,
            lcout => \uart_sync.aux_1__0_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4881\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_sync.aux_3__0__0_LC_7_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2330\,
            lcout => \uart_sync.aux_3__0_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4881\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNI34OR1_21_LC_7_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2458\,
            in1 => \N__2483\,
            in2 => \N__2543\,
            in3 => \N__2501\,
            lcout => \reset_module_System.reset6_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_5_LC_7_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101011001100"
        )
    port map (
            in0 => \N__3650\,
            in1 => \N__3061\,
            in2 => \N__2783\,
            in3 => \N__2528\,
            lcout => \uart.data_AuxZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4878\,
            ce => 'H',
            sr => \N__3455\
        );

    \uart.data_Aux_7_LC_7_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__3238\,
            in1 => \N__2781\,
            in2 => \N__3259\,
            in3 => \N__3652\,
            lcout => \uart.data_AuxZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4878\,
            ce => 'H',
            sr => \N__3455\
        );

    \uart.data_Aux_2_LC_7_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__2732\,
            in1 => \N__2777\,
            in2 => \N__3097\,
            in3 => \N__3651\,
            lcout => \uart.data_AuxZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4878\,
            ce => 'H',
            sr => \N__3455\
        );

    \uart.bit_Count_0_LC_7_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010010101010"
        )
    port map (
            in0 => \N__2601\,
            in1 => \N__2416\,
            in2 => \_gnd_net_\,
            in3 => \N__2721\,
            lcout => \uart.bit_CountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4875\,
            ce => 'H',
            sr => \N__5550\
        );

    \uart.state_RNI4ENK_3_LC_7_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110011001100"
        )
    port map (
            in0 => \N__2648\,
            in1 => \N__3371\,
            in2 => \N__2710\,
            in3 => \N__2600\,
            lcout => \uart.N_133_0\,
            ltout => \uart.N_133_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.bit_Count_1_LC_7_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110000011001100"
        )
    port map (
            in0 => \N__2602\,
            in1 => \N__2649\,
            in2 => \N__2420\,
            in3 => \N__2722\,
            lcout => \uart.bit_CountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4875\,
            ce => 'H',
            sr => \N__5550\
        );

    \uart.bit_Count_2_LC_7_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100001010000"
        )
    port map (
            in0 => \N__2723\,
            in1 => \N__2402\,
            in2 => \N__2711\,
            in3 => \N__2417\,
            lcout => \uart.bit_CountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4875\,
            ce => 'H',
            sr => \N__5550\
        );

    \uart.data_Aux_RNO_0_6_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__2651\,
            in1 => \N__2709\,
            in2 => \_gnd_net_\,
            in3 => \N__2604\,
            lcout => OPEN,
            ltout => \uart.data_Auxce_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_6_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101010001010"
        )
    port map (
            in0 => \N__4570\,
            in1 => \N__2782\,
            in2 => \N__2405\,
            in3 => \N__3672\,
            lcout => \uart.data_AuxZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4871\,
            ce => 'H',
            sr => \N__3454\
        );

    \uart.bit_Count_RNO_0_2_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__2603\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2650\,
            lcout => \uart.CO1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_1_cry_1_c_LC_8_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2892\,
            in2 => \N__3172\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_1_0_\,
            carryout => \reset_module_System.count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNO_0_2_LC_8_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2822\,
            in3 => \N__2447\,
            lcout => \reset_module_System.count_1_2\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_1\,
            carryout => \reset_module_System.count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_3_LC_8_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2990\,
            in2 => \_gnd_net_\,
            in3 => \N__2444\,
            lcout => \reset_module_System.countZ0Z_3\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_2\,
            carryout => \reset_module_System.count_1_cry_3\,
            clk => \N__4882\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_4_LC_8_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3034\,
            in2 => \_gnd_net_\,
            in3 => \N__2441\,
            lcout => \reset_module_System.countZ0Z_4\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_3\,
            carryout => \reset_module_System.count_1_cry_4\,
            clk => \N__4882\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_5_LC_8_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2921\,
            in2 => \_gnd_net_\,
            in3 => \N__2438\,
            lcout => \reset_module_System.countZ0Z_5\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_4\,
            carryout => \reset_module_System.count_1_cry_5\,
            clk => \N__4882\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_6_LC_8_1_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3002\,
            in2 => \_gnd_net_\,
            in3 => \N__2435\,
            lcout => \reset_module_System.countZ0Z_6\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_5\,
            carryout => \reset_module_System.count_1_cry_6\,
            clk => \N__4882\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_7_LC_8_1_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2948\,
            in2 => \_gnd_net_\,
            in3 => \N__2432\,
            lcout => \reset_module_System.countZ0Z_7\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_6\,
            carryout => \reset_module_System.count_1_cry_7\,
            clk => \N__4882\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_8_LC_8_1_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2960\,
            in2 => \_gnd_net_\,
            in3 => \N__2429\,
            lcout => \reset_module_System.countZ0Z_8\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_7\,
            carryout => \reset_module_System.count_1_cry_8\,
            clk => \N__4882\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_9_LC_8_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2935\,
            in2 => \_gnd_net_\,
            in3 => \N__2426\,
            lcout => \reset_module_System.countZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_8_2_0_\,
            carryout => \reset_module_System.count_1_cry_9\,
            clk => \N__4879\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_10_LC_8_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2795\,
            in2 => \_gnd_net_\,
            in3 => \N__2423\,
            lcout => \reset_module_System.countZ0Z_10\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_9\,
            carryout => \reset_module_System.count_1_cry_10\,
            clk => \N__4879\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_11_LC_8_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2807\,
            in2 => \_gnd_net_\,
            in3 => \N__2507\,
            lcout => \reset_module_System.countZ0Z_11\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_10\,
            carryout => \reset_module_System.count_1_cry_11\,
            clk => \N__4879\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_12_LC_8_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3184\,
            in2 => \_gnd_net_\,
            in3 => \N__2504\,
            lcout => \reset_module_System.countZ0Z_12\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_11\,
            carryout => \reset_module_System.count_1_cry_12\,
            clk => \N__4879\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_13_LC_8_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2500\,
            in2 => \_gnd_net_\,
            in3 => \N__2489\,
            lcout => \reset_module_System.countZ0Z_13\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_12\,
            carryout => \reset_module_System.count_1_cry_13\,
            clk => \N__4879\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_14_LC_8_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3218\,
            in2 => \_gnd_net_\,
            in3 => \N__2486\,
            lcout => \reset_module_System.countZ0Z_14\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_13\,
            carryout => \reset_module_System.count_1_cry_14\,
            clk => \N__4879\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_15_LC_8_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2482\,
            in2 => \_gnd_net_\,
            in3 => \N__2471\,
            lcout => \reset_module_System.countZ0Z_15\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_14\,
            carryout => \reset_module_System.count_1_cry_15\,
            clk => \N__4879\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_16_LC_8_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3046\,
            in2 => \_gnd_net_\,
            in3 => \N__2468\,
            lcout => \reset_module_System.countZ0Z_16\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_15\,
            carryout => \reset_module_System.count_1_cry_16\,
            clk => \N__4879\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_17_LC_8_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3206\,
            in2 => \_gnd_net_\,
            in3 => \N__2465\,
            lcout => \reset_module_System.countZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_8_3_0_\,
            carryout => \reset_module_System.count_1_cry_17\,
            clk => \N__4876\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_18_LC_8_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3019\,
            in2 => \_gnd_net_\,
            in3 => \N__2462\,
            lcout => \reset_module_System.countZ0Z_18\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_17\,
            carryout => \reset_module_System.count_1_cry_18\,
            clk => \N__4876\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_19_LC_8_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2459\,
            in2 => \_gnd_net_\,
            in3 => \N__2552\,
            lcout => \reset_module_System.countZ0Z_19\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_18\,
            carryout => \reset_module_System.count_1_cry_19\,
            clk => \N__4876\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_20_LC_8_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2974\,
            in2 => \_gnd_net_\,
            in3 => \N__2549\,
            lcout => \reset_module_System.countZ0Z_20\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_19\,
            carryout => \reset_module_System.count_1_cry_20\,
            clk => \N__4876\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_21_LC_8_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2542\,
            in2 => \_gnd_net_\,
            in3 => \N__2546\,
            lcout => \reset_module_System.countZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4876\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.bit_Count_RNIETHE_2_LC_8_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__2696\,
            in1 => \N__2644\,
            in2 => \_gnd_net_\,
            in3 => \N__2598\,
            lcout => \uart.N_177\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_RNO_0_5_LC_8_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__2599\,
            in1 => \_gnd_net_\,
            in2 => \N__2661\,
            in3 => \N__2697\,
            lcout => \uart.data_Auxce_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_RNI9M0N_1_LC_8_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100010001"
        )
    port map (
            in0 => \N__3334\,
            in1 => \N__3505\,
            in2 => \_gnd_net_\,
            in3 => \N__4156\,
            lcout => \uart.timer_Count_RNI9M0NZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_RNILKMA1_0_LC_8_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__3929\,
            in1 => \N__3971\,
            in2 => \N__4328\,
            in3 => \N__3890\,
            lcout => OPEN,
            ltout => \uart.timer_Count_RNILKMA1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNILC8T2_3_LC_8_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110111011101"
        )
    port map (
            in0 => \N__2522\,
            in1 => \N__3361\,
            in2 => \N__2513\,
            in3 => \N__4003\,
            lcout => \uart.un1_state_2_0\,
            ltout => \uart.un1_state_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_0_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111010100010"
        )
    port map (
            in0 => \N__3109\,
            in1 => \N__2744\,
            in2 => \N__2510\,
            in3 => \N__3670\,
            lcout => \uart.data_AuxZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4872\,
            ce => 'H',
            sr => \N__3453\
        );

    \uart.data_Aux_1_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__3668\,
            in1 => \N__2738\,
            in2 => \N__4240\,
            in3 => \N__2774\,
            lcout => \uart.data_AuxZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4872\,
            ce => 'H',
            sr => \N__3453\
        );

    \uart.data_Aux_3_LC_8_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101100"
        )
    port map (
            in0 => \N__3669\,
            in1 => \N__3080\,
            in2 => \N__2561\,
            in3 => \N__2775\,
            lcout => \uart.data_AuxZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4872\,
            ce => 'H',
            sr => \N__3453\
        );

    \uart.data_Aux_4_LC_8_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__2776\,
            in1 => \N__2750\,
            in2 => \N__4600\,
            in3 => \N__3671\,
            lcout => \uart.data_AuxZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4872\,
            ce => 'H',
            sr => \N__3453\
        );

    \uart.data_Aux_RNO_0_4_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__2609\,
            in1 => \_gnd_net_\,
            in2 => \N__2663\,
            in3 => \N__2708\,
            lcout => \uart.data_Auxce_0_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_RNO_0_0_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__2704\,
            in1 => \N__2652\,
            in2 => \_gnd_net_\,
            in3 => \N__2605\,
            lcout => \uart.data_Auxce_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_RNO_0_1_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001010"
        )
    port map (
            in0 => \N__2606\,
            in1 => \_gnd_net_\,
            in2 => \N__2662\,
            in3 => \N__2705\,
            lcout => \uart.data_Auxce_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_RNO_0_2_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__2706\,
            in1 => \N__2656\,
            in2 => \_gnd_net_\,
            in3 => \N__2607\,
            lcout => \uart.data_Auxce_0_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNIA73N2_4_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100010001"
        )
    port map (
            in0 => \N__3362\,
            in1 => \N__3511\,
            in2 => \_gnd_net_\,
            in3 => \N__3565\,
            lcout => \uart.un1_state_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_RNO_0_3_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__2707\,
            in1 => \N__2657\,
            in2 => \_gnd_net_\,
            in3 => \N__2608\,
            lcout => \uart.data_Auxce_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_0_LC_9_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010101010101"
        )
    port map (
            in0 => \N__3171\,
            in1 => \N__2841\,
            in2 => \N__2876\,
            in3 => \N__3133\,
            lcout => \reset_module_System.countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4880\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNI10J41_1_LC_9_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__3050\,
            in1 => \N__3035\,
            in2 => \N__3023\,
            in3 => \N__2893\,
            lcout => \reset_module_System.reset6_14\,
            ltout => \reset_module_System.reset6_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.reset_LC_9_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111111111111"
        )
    port map (
            in0 => \N__2867\,
            in1 => \_gnd_net_\,
            in2 => \N__3005\,
            in3 => \N__3131\,
            lcout => reset_system,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4880\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNI9O1P_2_LC_9_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__3001\,
            in1 => \N__2989\,
            in2 => \N__2978\,
            in3 => \N__2818\,
            lcout => \reset_module_System.reset6_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.reset_iso_LC_9_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__2868\,
            in1 => \N__2840\,
            in2 => \_gnd_net_\,
            in3 => \N__3132\,
            lcout => \reset_module_System_reset_iso\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4880\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNI97FD_5_LC_9_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2959\,
            in1 => \N__2947\,
            in2 => \N__2936\,
            in3 => \N__2920\,
            lcout => \reset_module_System.reset6_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_1_LC_9_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__2909\,
            in1 => \N__2842\,
            in2 => \N__2875\,
            in3 => \N__3134\,
            lcout => \reset_module_System.countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4880\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_2_LC_9_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3130\,
            in1 => \N__2866\,
            in2 => \N__2846\,
            in3 => \N__2828\,
            lcout => \reset_module_System.countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4880\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNIP8RT_10_LC_9_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__2806\,
            in1 => \N__2794\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \reset_module_System.reset6_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNI53692_14_LC_9_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3217\,
            in1 => \N__3205\,
            in2 => \N__3194\,
            in3 => \N__3191\,
            lcout => OPEN,
            ltout => \reset_module_System.reset6_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNIN3HK3_12_LC_9_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__3185\,
            in1 => \N__3170\,
            in2 => \N__3143\,
            in3 => \N__3140\,
            lcout => \reset_module_System.reset6_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNO_1_3_LC_9_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__3352\,
            in1 => \N__3787\,
            in2 => \N__3404\,
            in3 => \N__3818\,
            lcout => OPEN,
            ltout => \uart.N_169_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNO_0_3_LC_9_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001011"
        )
    port map (
            in0 => \N__3848\,
            in1 => \N__3305\,
            in2 => \N__3116\,
            in3 => \N__5359\,
            lcout => OPEN,
            ltout => \uart.state_srsts_i_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_3_LC_9_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000011110000"
        )
    port map (
            in0 => \N__3239\,
            in1 => \N__3403\,
            in2 => \N__3113\,
            in3 => \N__3572\,
            lcout => \uart.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4877\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_esr_0_LC_9_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3110\,
            lcout => uart_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4873\,
            ce => \N__4547\,
            sr => \N__4529\
        );

    \uart.data_esr_2_LC_9_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3098\,
            lcout => uart_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4873\,
            ce => \N__4547\,
            sr => \N__4529\
        );

    \uart.data_esr_3_LC_9_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3079\,
            lcout => uart_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4873\,
            ce => \N__4547\,
            sr => \N__4529\
        );

    \uart.data_esr_5_LC_9_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3065\,
            lcout => uart_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4873\,
            ce => \N__4547\,
            sr => \N__4529\
        );

    \uart.data_esr_7_LC_9_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3260\,
            lcout => uart_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4873\,
            ce => \N__4547\,
            sr => \N__4529\
        );

    \uart.timer_Count_RNI22NA1_6_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__3880\,
            in1 => \N__3813\,
            in2 => \N__3780\,
            in3 => \N__3842\,
            lcout => OPEN,
            ltout => \uart.timer_Count10lto5_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_RNIT4OA2_2_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000010100000"
        )
    port map (
            in0 => \N__3843\,
            in1 => \N__3920\,
            in2 => \N__3242\,
            in3 => \N__3967\,
            lcout => \uart.N_180\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_RNI1HBL_6_LC_9_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3841\,
            in2 => \_gnd_net_\,
            in3 => \N__3812\,
            lcout => \uart.N_145_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_1_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001000000"
        )
    port map (
            in0 => \N__5362\,
            in1 => \N__3422\,
            in2 => \N__3683\,
            in3 => \N__3287\,
            lcout => \uart.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4868\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNIMO1Q_4_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__3770\,
            in1 => \N__3500\,
            in2 => \_gnd_net_\,
            in3 => \N__5360\,
            lcout => \uart.state_srsts_0_a3_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNO_0_4_LC_9_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__5361\,
            in1 => \N__3237\,
            in2 => \N__3370\,
            in3 => \N__3566\,
            lcout => OPEN,
            ltout => \uart.N_168_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_4_LC_9_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__3587\,
            in1 => \_gnd_net_\,
            in2 => \N__3221\,
            in3 => \_gnd_net_\,
            lcout => \uart.stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4868\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNIB0BC_2_LC_9_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3392\,
            in2 => \_gnd_net_\,
            in3 => \N__3356\,
            lcout => \uart.N_159\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNIAFHL_4_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__3360\,
            in1 => \N__3512\,
            in2 => \_gnd_net_\,
            in3 => \N__5376\,
            lcout => \uart.state_RNIAFHLZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNO_0_2_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__3420\,
            in1 => \N__3396\,
            in2 => \_gnd_net_\,
            in3 => \N__3676\,
            lcout => OPEN,
            ltout => \uart.N_151_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_2_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010000000101"
        )
    port map (
            in0 => \N__5378\,
            in1 => \N__3421\,
            in2 => \N__3407\,
            in3 => \N__3571\,
            lcout => \uart.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4866\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNO_2_3_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__3924\,
            in1 => \N__3964\,
            in2 => \N__3369\,
            in3 => \N__3884\,
            lcout => \uart.state_srsts_i_1_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNO_1_0_LC_10_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3788\,
            in2 => \_gnd_net_\,
            in3 => \N__3520\,
            lcout => OPEN,
            ltout => \uart.N_166_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNO_0_0_LC_10_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001101"
        )
    port map (
            in0 => \N__3283\,
            in1 => \N__3681\,
            in2 => \N__3293\,
            in3 => \N__5358\,
            lcout => OPEN,
            ltout => \uart.state_srsts_0_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_0_LC_10_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111100001111"
        )
    port map (
            in0 => \N__3521\,
            in1 => \N__3539\,
            in2 => \N__3290\,
            in3 => \N__4007\,
            lcout => \uart.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4874\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_10_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.count_2_LC_10_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010100110"
        )
    port map (
            in0 => \N__4061\,
            in1 => \N__4081\,
            in2 => \N__3272\,
            in3 => \N__4094\,
            lcout => \uart_frame_decoder.countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4874\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.count_RNIV5MS_0_LC_10_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__5030\,
            in1 => \N__5455\,
            in2 => \_gnd_net_\,
            in3 => \N__4037\,
            lcout => \uart_frame_decoder.N_43\,
            ltout => \uart_frame_decoder.N_43_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.count_1_LC_10_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4080\,
            in2 => \N__3467\,
            in3 => \N__4093\,
            lcout => \uart_frame_decoder.countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4874\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNIMBMF_1_LC_10_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5026\,
            in2 => \_gnd_net_\,
            in3 => \N__5215\,
            lcout => \uart_frame_decoder.state_1_ns_i_i_a2_1_1_0\,
            ltout => \uart_frame_decoder.state_1_ns_i_i_a2_1_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNO_1_0_LC_10_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010000000"
        )
    port map (
            in0 => \N__3692\,
            in1 => \N__4269\,
            in2 => \N__3464\,
            in3 => \N__4255\,
            lcout => OPEN,
            ltout => \uart_frame_decoder.N_81_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_0_LC_10_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__4166\,
            in1 => \N__4927\,
            in2 => \N__3461\,
            in3 => \N__4334\,
            lcout => \uart_frame_decoder.state_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4869\,
            ce => 'H',
            sr => \N__5536\
        );

    \uart_frame_decoder.state_1_ns_0_i_a2_0_0_1_2_LC_10_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3721\,
            in2 => \_gnd_net_\,
            in3 => \N__3700\,
            lcout => OPEN,
            ltout => \uart_frame_decoder.state_1_ns_0_i_a2_0_0_1Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNI5BVV_1_LC_10_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__5207\,
            in1 => \N__3709\,
            in2 => \N__3458\,
            in3 => \N__3730\,
            lcout => \uart_frame_decoder.N_92\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNO_3_0_LC_10_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011101"
        )
    port map (
            in0 => \N__4182\,
            in1 => \N__5206\,
            in2 => \_gnd_net_\,
            in3 => \N__5422\,
            lcout => \uart_frame_decoder.state_1_ns_i_i_a2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_rdy_LC_10_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__3980\,
            in1 => \N__3677\,
            in2 => \_gnd_net_\,
            in3 => \N__5368\,
            lcout => uart_data_rdy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4867\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_ns_0_i_a2_1_0_2_LC_10_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5423\,
            in2 => \_gnd_net_\,
            in3 => \N__4583\,
            lcout => OPEN,
            ltout => \uart_frame_decoder.state_1_ns_0_i_a2_1_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_ns_0_i_a2_1_2_LC_10_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4559\,
            in1 => \N__3740\,
            in2 => \N__3734\,
            in3 => \N__4223\,
            lcout => \uart_frame_decoder.N_99\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_ns_0_i_a2_0_4_1_LC_10_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3731\,
            in1 => \N__3722\,
            in2 => \N__3713\,
            in3 => \N__3701\,
            lcout => \uart_frame_decoder.N_79_4\,
            ltout => \uart_frame_decoder.N_79_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNO_0_1_LC_10_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3686\,
            in3 => \N__4183\,
            lcout => \uart_frame_decoder.state_1_ns_0_i_a2_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNI78E91_4_LC_10_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001000"
        )
    port map (
            in0 => \N__3501\,
            in1 => \N__3771\,
            in2 => \N__3682\,
            in3 => \N__4000\,
            lcout => OPEN,
            ltout => \uart.data_8_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_RNIS4183_7_LC_10_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011111100"
        )
    port map (
            in0 => \N__3772\,
            in1 => \N__5363\,
            in2 => \N__3599\,
            in3 => \N__3534\,
            lcout => \uart.timer_Count_RNIS4183Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_RNIMLMA1_1_LC_10_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__4148\,
            in1 => \N__3966\,
            in2 => \N__3886\,
            in3 => \N__3919\,
            lcout => \uart.N_152_0\,
            ltout => \uart.N_152_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNIDV3Q2_4_LC_10_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3596\,
            in2 => \N__3590\,
            in3 => \N__4001\,
            lcout => \uart.N_167\,
            ltout => \uart.N_167_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNIIHDQ5_2_LC_10_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111001110"
        )
    port map (
            in0 => \N__3581\,
            in1 => \N__5364\,
            in2 => \N__3575\,
            in3 => \N__3567\,
            lcout => \uart.timer_Count_1_sqmuxa_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNIGITG2_4_LC_10_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000011000000"
        )
    port map (
            in0 => \N__3535\,
            in1 => \N__3773\,
            in2 => \N__3513\,
            in3 => \N__4002\,
            lcout => \uart.state_1_sqmuxa\,
            ltout => \uart.state_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNICNUO5_4_LC_10_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3974\,
            in3 => \N__4515\,
            lcout => \uart.state_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.un4_timer_Count_1_cry_1_c_LC_10_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4324\,
            in2 => \N__4160\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_5_0_\,
            carryout => \uart.un4_timer_Count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_2_LC_10_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3965\,
            in2 => \_gnd_net_\,
            in3 => \N__3932\,
            lcout => \uart.timer_CountZ0Z_2\,
            ltout => OPEN,
            carryin => \uart.un4_timer_Count_1_cry_1\,
            carryout => \uart.un4_timer_Count_1_cry_2\,
            clk => \N__4862\,
            ce => 'H',
            sr => \N__4294\
        );

    \uart.timer_Count_3_LC_10_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3925\,
            in2 => \_gnd_net_\,
            in3 => \N__3893\,
            lcout => \uart.timer_CountZ0Z_3\,
            ltout => OPEN,
            carryin => \uart.un4_timer_Count_1_cry_2\,
            carryout => \uart.un4_timer_Count_1_cry_3\,
            clk => \N__4862\,
            ce => 'H',
            sr => \N__4294\
        );

    \uart.timer_Count_4_LC_10_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3885\,
            in2 => \_gnd_net_\,
            in3 => \N__3851\,
            lcout => \uart.timer_CountZ0Z_4\,
            ltout => OPEN,
            carryin => \uart.un4_timer_Count_1_cry_3\,
            carryout => \uart.un4_timer_Count_1_cry_4\,
            clk => \N__4862\,
            ce => 'H',
            sr => \N__4294\
        );

    \uart.timer_Count_5_LC_10_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3847\,
            in2 => \_gnd_net_\,
            in3 => \N__3821\,
            lcout => \uart.timer_CountZ0Z_5\,
            ltout => OPEN,
            carryin => \uart.un4_timer_Count_1_cry_4\,
            carryout => \uart.un4_timer_Count_1_cry_5\,
            clk => \N__4862\,
            ce => 'H',
            sr => \N__4294\
        );

    \uart.timer_Count_6_LC_10_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3817\,
            in2 => \_gnd_net_\,
            in3 => \N__3794\,
            lcout => \uart.timer_CountZ0Z_6\,
            ltout => OPEN,
            carryin => \uart.un4_timer_Count_1_cry_5\,
            carryout => \uart.un4_timer_Count_1_cry_6\,
            clk => \N__4862\,
            ce => 'H',
            sr => \N__4294\
        );

    \uart.timer_Count_7_LC_10_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3779\,
            in2 => \_gnd_net_\,
            in3 => \N__3791\,
            lcout => \uart.timer_CountZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4862\,
            ce => 'H',
            sr => \N__4294\
        );

    \uart_frame_decoder.count8_cry_0_c_LC_11_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4019\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_1_0_\,
            carryout => \uart_frame_decoder.count8_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.count8_cry_1_c_inv_LC_11_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4127\,
            in3 => \N__4076\,
            lcout => \uart_frame_decoder.count8_axb_1\,
            ltout => OPEN,
            carryin => \uart_frame_decoder.count8_cry_0\,
            carryout => \uart_frame_decoder.count8_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.count8_cry_2_c_inv_LC_11_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4046\,
            in2 => \N__4118\,
            in3 => \N__4059\,
            lcout => \uart_frame_decoder.count_i_2\,
            ltout => OPEN,
            carryin => \uart_frame_decoder.count8_cry_1\,
            carryout => \uart_frame_decoder.count8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.count8_THRU_LUT4_0_LC_11_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4109\,
            lcout => \uart_frame_decoder.count8_THRU_CO\,
            ltout => \uart_frame_decoder.count8_THRU_CO_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.count8_cry_2_c_RNICKS21_LC_11_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001000"
        )
    port map (
            in0 => \N__5031\,
            in1 => \N__5458\,
            in2 => \N__4097\,
            in3 => \N__5372\,
            lcout => \uart_frame_decoder.N_37\,
            ltout => \uart_frame_decoder.N_37_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.count_0_LC_11_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100001000"
        )
    port map (
            in0 => \N__5459\,
            in1 => \N__5032\,
            in2 => \N__4085\,
            in3 => \N__4036\,
            lcout => \uart_frame_decoder.count8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4870\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.count_RNIHPR51_2_LC_11_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010111111111"
        )
    port map (
            in0 => \N__4035\,
            in1 => \_gnd_net_\,
            in2 => \N__4082\,
            in3 => \N__4060\,
            lcout => \uart_frame_decoder.state_1_ns_0_i_o2_0_tz_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.count8_cry_0_c_inv_LC_11_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__4045\,
            in1 => \N__4018\,
            in2 => \_gnd_net_\,
            in3 => \N__4034\,
            lcout => \uart_frame_decoder.count8_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.WDT_RNIOAVK1_5_LC_11_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011100110011"
        )
    port map (
            in0 => \N__4800\,
            in1 => \N__4727\,
            in2 => \N__4430\,
            in3 => \N__4205\,
            lcout => OPEN,
            ltout => \uart_frame_decoder.N_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.WDT_RNIGSL62_15_LC_11_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011101010101"
        )
    port map (
            in0 => \N__4953\,
            in1 => \N__4661\,
            in2 => \N__4214\,
            in3 => \N__4211\,
            lcout => \uart_frame_decoder.WDT8_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.WDT_RNIEKPB_11_LC_11_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000011111"
        )
    port map (
            in0 => \N__4704\,
            in1 => \N__4683\,
            in2 => \N__4664\,
            in3 => \N__4639\,
            lcout => \uart_frame_decoder.g0_1_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.WDT_RNIRBB11_4_LC_11_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4780\,
            in1 => \N__4446\,
            in2 => \N__4403\,
            in3 => \N__4752\,
            lcout => \uart_frame_decoder.g0_1_a3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.WDT_RNIQAB11_4_LC_11_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4447\,
            in1 => \N__4425\,
            in2 => \N__4781\,
            in3 => \N__4753\,
            lcout => \uart_frame_decoder.WDT_RNIQAB11Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.WDT_RNIVBR8_15_LC_11_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010100000"
        )
    port map (
            in0 => \N__4640\,
            in1 => \_gnd_net_\,
            in2 => \N__4955\,
            in3 => \N__4662\,
            lcout => \uart_frame_decoder.WDT8lto15\,
            ltout => \uart_frame_decoder.WDT8lto15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNILEPU1_10_LC_11_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110000000100"
        )
    port map (
            in0 => \N__5456\,
            in1 => \N__5017\,
            in2 => \N__4199\,
            in3 => \N__4196\,
            lcout => \uart_frame_decoder.state_1_ns_0_i_a2_0_0_0_10\,
            ltout => \uart_frame_decoder.state_1_ns_0_i_a2_0_0_0_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNO_2_0_LC_11_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001111"
        )
    port map (
            in0 => \N__4190\,
            in1 => \N__4184\,
            in2 => \N__4169\,
            in3 => \N__5457\,
            lcout => \uart_frame_decoder.N_35_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_1_LC_11_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4320\,
            in2 => \_gnd_net_\,
            in3 => \N__4155\,
            lcout => \uart.timer_CountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4865\,
            ce => 'H',
            sr => \N__4295\
        );

    \uart_frame_decoder.WDT_RNISS5H_11_LC_11_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100010001"
        )
    port map (
            in0 => \N__4684\,
            in1 => \N__4705\,
            in2 => \N__4733\,
            in3 => \N__4401\,
            lcout => OPEN,
            ltout => \uart_frame_decoder.WDT_RNISS5HZ0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.WDT_RNIEDQT1_7_LC_11_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010110000"
        )
    port map (
            in0 => \N__4379\,
            in1 => \N__4731\,
            in2 => \N__4373\,
            in3 => \N__4801\,
            lcout => \uart_frame_decoder.WDT8lt13\,
            ltout => \uart_frame_decoder.WDT8lt13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.WDT_RNIKVEI2_14_LC_11_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101010001"
        )
    port map (
            in0 => \N__5443\,
            in1 => \N__4345\,
            in2 => \N__4370\,
            in3 => \N__4631\,
            lcout => \uart_frame_decoder.N_85\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.WDT_RNI85RG2_14_LC_11_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__4630\,
            in1 => \N__5008\,
            in2 => \N__4361\,
            in3 => \N__5444\,
            lcout => \uart_frame_decoder.state_1_ns_0_i_a2_0_d_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNO_0_0_LC_11_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010001010"
        )
    port map (
            in0 => \N__4367\,
            in1 => \N__4357\,
            in2 => \N__4349\,
            in3 => \N__4632\,
            lcout => \uart_frame_decoder.N_80\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_0_LC_11_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4319\,
            lcout => \uart.timer_CountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4865\,
            ce => 'H',
            sr => \N__4295\
        );

    \uart_frame_decoder.state_1_1_LC_11_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__5211\,
            in1 => \N__4270\,
            in2 => \N__4283\,
            in3 => \N__4908\,
            lcout => \uart_frame_decoder.state_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4863\,
            ce => 'H',
            sr => \N__5549\
        );

    \uart_frame_decoder.state_1_2_LC_11_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__4909\,
            in1 => \N__5074\,
            in2 => \N__4274\,
            in3 => \N__4256\,
            lcout => \uart_frame_decoder.state_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4863\,
            ce => 'H',
            sr => \N__5549\
        );

    \uart.data_esr_1_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4244\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => uart_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4860\,
            ce => \N__4546\,
            sr => \N__4528\
        );

    \uart.data_esr_4_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4604\,
            lcout => uart_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4860\,
            ce => \N__4546\,
            sr => \N__4528\
        );

    \uart.data_esr_6_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4574\,
            lcout => uart_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4860\,
            ce => \N__4546\,
            sr => \N__4528\
        );

    \uart_frame_decoder.WDT_0_LC_12_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4481\,
            in2 => \N__4498\,
            in3 => \N__4499\,
            lcout => \uart_frame_decoder.WDTZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_12_2_0_\,
            carryout => \uart_frame_decoder.un1_WDT_cry_0\,
            clk => \N__4864\,
            ce => 'H',
            sr => \N__5300\
        );

    \uart_frame_decoder.WDT_1_LC_12_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4475\,
            in2 => \_gnd_net_\,
            in3 => \N__4469\,
            lcout => \uart_frame_decoder.WDTZ0Z_1\,
            ltout => OPEN,
            carryin => \uart_frame_decoder.un1_WDT_cry_0\,
            carryout => \uart_frame_decoder.un1_WDT_cry_1\,
            clk => \N__4864\,
            ce => 'H',
            sr => \N__5300\
        );

    \uart_frame_decoder.WDT_2_LC_12_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4466\,
            in2 => \_gnd_net_\,
            in3 => \N__4460\,
            lcout => \uart_frame_decoder.WDTZ0Z_2\,
            ltout => OPEN,
            carryin => \uart_frame_decoder.un1_WDT_cry_1\,
            carryout => \uart_frame_decoder.un1_WDT_cry_2\,
            clk => \N__4864\,
            ce => 'H',
            sr => \N__5300\
        );

    \uart_frame_decoder.WDT_3_LC_12_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4457\,
            in2 => \_gnd_net_\,
            in3 => \N__4451\,
            lcout => \uart_frame_decoder.WDTZ0Z_3\,
            ltout => OPEN,
            carryin => \uart_frame_decoder.un1_WDT_cry_2\,
            carryout => \uart_frame_decoder.un1_WDT_cry_3\,
            clk => \N__4864\,
            ce => 'H',
            sr => \N__5300\
        );

    \uart_frame_decoder.WDT_4_LC_12_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4448\,
            in2 => \_gnd_net_\,
            in3 => \N__4433\,
            lcout => \uart_frame_decoder.WDTZ0Z_4\,
            ltout => OPEN,
            carryin => \uart_frame_decoder.un1_WDT_cry_3\,
            carryout => \uart_frame_decoder.un1_WDT_cry_4\,
            clk => \N__4864\,
            ce => 'H',
            sr => \N__5300\
        );

    \uart_frame_decoder.WDT_5_LC_12_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4426\,
            in2 => \_gnd_net_\,
            in3 => \N__4406\,
            lcout => \uart_frame_decoder.WDTZ0Z_5\,
            ltout => OPEN,
            carryin => \uart_frame_decoder.un1_WDT_cry_4\,
            carryout => \uart_frame_decoder.un1_WDT_cry_5\,
            clk => \N__4864\,
            ce => 'H',
            sr => \N__5300\
        );

    \uart_frame_decoder.WDT_6_LC_12_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4402\,
            in2 => \_gnd_net_\,
            in3 => \N__4382\,
            lcout => \uart_frame_decoder.WDTZ0Z_6\,
            ltout => OPEN,
            carryin => \uart_frame_decoder.un1_WDT_cry_5\,
            carryout => \uart_frame_decoder.un1_WDT_cry_6\,
            clk => \N__4864\,
            ce => 'H',
            sr => \N__5300\
        );

    \uart_frame_decoder.WDT_7_LC_12_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4802\,
            in2 => \_gnd_net_\,
            in3 => \N__4784\,
            lcout => \uart_frame_decoder.WDTZ0Z_7\,
            ltout => OPEN,
            carryin => \uart_frame_decoder.un1_WDT_cry_6\,
            carryout => \uart_frame_decoder.un1_WDT_cry_7\,
            clk => \N__4864\,
            ce => 'H',
            sr => \N__5300\
        );

    \uart_frame_decoder.WDT_8_LC_12_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4779\,
            in2 => \_gnd_net_\,
            in3 => \N__4757\,
            lcout => \uart_frame_decoder.WDTZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_12_3_0_\,
            carryout => \uart_frame_decoder.un1_WDT_cry_8\,
            clk => \N__4861\,
            ce => 'H',
            sr => \N__5296\
        );

    \uart_frame_decoder.WDT_9_LC_12_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4754\,
            in2 => \_gnd_net_\,
            in3 => \N__4736\,
            lcout => \uart_frame_decoder.WDTZ0Z_9\,
            ltout => OPEN,
            carryin => \uart_frame_decoder.un1_WDT_cry_8\,
            carryout => \uart_frame_decoder.un1_WDT_cry_9\,
            clk => \N__4861\,
            ce => 'H',
            sr => \N__5296\
        );

    \uart_frame_decoder.WDT_10_LC_12_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4732\,
            in2 => \_gnd_net_\,
            in3 => \N__4709\,
            lcout => \uart_frame_decoder.WDTZ0Z_10\,
            ltout => OPEN,
            carryin => \uart_frame_decoder.un1_WDT_cry_9\,
            carryout => \uart_frame_decoder.un1_WDT_cry_10\,
            clk => \N__4861\,
            ce => 'H',
            sr => \N__5296\
        );

    \uart_frame_decoder.WDT_11_LC_12_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4706\,
            in2 => \_gnd_net_\,
            in3 => \N__4688\,
            lcout => \uart_frame_decoder.WDTZ0Z_11\,
            ltout => OPEN,
            carryin => \uart_frame_decoder.un1_WDT_cry_10\,
            carryout => \uart_frame_decoder.un1_WDT_cry_11\,
            clk => \N__4861\,
            ce => 'H',
            sr => \N__5296\
        );

    \uart_frame_decoder.WDT_12_LC_12_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4685\,
            in2 => \_gnd_net_\,
            in3 => \N__4667\,
            lcout => \uart_frame_decoder.WDTZ0Z_12\,
            ltout => OPEN,
            carryin => \uart_frame_decoder.un1_WDT_cry_11\,
            carryout => \uart_frame_decoder.un1_WDT_cry_12\,
            clk => \N__4861\,
            ce => 'H',
            sr => \N__5296\
        );

    \uart_frame_decoder.WDT_13_LC_12_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4663\,
            in2 => \_gnd_net_\,
            in3 => \N__4643\,
            lcout => \uart_frame_decoder.WDTZ0Z_13\,
            ltout => OPEN,
            carryin => \uart_frame_decoder.un1_WDT_cry_12\,
            carryout => \uart_frame_decoder.un1_WDT_cry_13\,
            clk => \N__4861\,
            ce => 'H',
            sr => \N__5296\
        );

    \uart_frame_decoder.WDT_14_LC_12_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4633\,
            in2 => \_gnd_net_\,
            in3 => \N__4607\,
            lcout => \uart_frame_decoder.WDTZ0Z_14\,
            ltout => OPEN,
            carryin => \uart_frame_decoder.un1_WDT_cry_13\,
            carryout => \uart_frame_decoder.un1_WDT_cry_14\,
            clk => \N__4861\,
            ce => 'H',
            sr => \N__5296\
        );

    \uart_frame_decoder.WDT_15_LC_12_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4954\,
            in2 => \_gnd_net_\,
            in3 => \N__4958\,
            lcout => \uart_frame_decoder.WDTZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4861\,
            ce => 'H',
            sr => \N__5296\
        );

    \uart_frame_decoder.state_1_10_LC_12_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111101010"
        )
    port map (
            in0 => \N__4937\,
            in1 => \N__5495\,
            in2 => \N__5183\,
            in3 => \N__4928\,
            lcout => \uart_frame_decoder.state_1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4859\,
            ce => 'H',
            sr => \N__5552\
        );

    \uart_frame_decoder.state_1_3_LC_12_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__5491\,
            in1 => \N__5073\,
            in2 => \N__5057\,
            in3 => \N__4910\,
            lcout => \uart_frame_decoder.state_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4859\,
            ce => 'H',
            sr => \N__5552\
        );

    \uart_frame_decoder.state_1_4_LC_12_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__4911\,
            in1 => \N__5496\,
            in2 => \N__5279\,
            in3 => \N__5051\,
            lcout => \uart_frame_decoder.state_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4859\,
            ce => 'H',
            sr => \N__5552\
        );

    \uart_frame_decoder.state_1_5_LC_12_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__5492\,
            in1 => \N__5274\,
            in2 => \N__5159\,
            in3 => \N__4912\,
            lcout => \uart_frame_decoder.state_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4859\,
            ce => 'H',
            sr => \N__5552\
        );

    \uart_frame_decoder.state_1_6_LC_12_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__4913\,
            in1 => \N__5497\,
            in2 => \N__5123\,
            in3 => \N__5153\,
            lcout => \uart_frame_decoder.state_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4859\,
            ce => 'H',
            sr => \N__5552\
        );

    \uart_frame_decoder.state_1_7_LC_12_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__5493\,
            in1 => \N__5118\,
            in2 => \N__5105\,
            in3 => \N__4914\,
            lcout => \uart_frame_decoder.state_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4859\,
            ce => 'H',
            sr => \N__5552\
        );

    \uart_frame_decoder.state_1_8_LC_12_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__4915\,
            in1 => \N__5102\,
            in2 => \N__5504\,
            in3 => \N__5244\,
            lcout => \uart_frame_decoder.state_1Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4859\,
            ce => 'H',
            sr => \N__5552\
        );

    \uart_frame_decoder.state_1_9_LC_12_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__5494\,
            in1 => \N__5180\,
            in2 => \N__5246\,
            in3 => \N__4916\,
            lcout => \uart_frame_decoder.state_1Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4859\,
            ce => 'H',
            sr => \N__5552\
        );

    \uart_frame_decoder.source_data_valid_2_sqmuxa_i_LC_13_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5460\,
            in2 => \_gnd_net_\,
            in3 => \N__5377\,
            lcout => \uart_frame_decoder.source_data_valid_2_sqmuxa_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNIUQR11_4_LC_13_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__5278\,
            in1 => \N__5084\,
            in2 => \_gnd_net_\,
            in3 => \N__5158\,
            lcout => \uart_frame_decoder_N_307_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNI8L5O_8_LC_13_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__5009\,
            in1 => \N__5245\,
            in2 => \_gnd_net_\,
            in3 => \N__5182\,
            lcout => \uart_frame_decoder_N_308_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNICQTG_7_LC_13_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5103\,
            in2 => \_gnd_net_\,
            in3 => \N__5216\,
            lcout => OPEN,
            ltout => \uart_frame_decoder.un14_i_a2_0_a2_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNI3NAA1_3_LC_13_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__5181\,
            in1 => \N__5055\,
            in2 => \N__5162\,
            in3 => \N__5157\,
            lcout => \uart_frame_decoder_N_305_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNIHVTG_6_LC_13_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__5122\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5104\,
            lcout => \uart_frame_decoder.N_306_1\,
            ltout => \uart_frame_decoder.N_306_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNID8391_2_LC_13_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__5078\,
            in1 => \N__5056\,
            in2 => \N__5036\,
            in3 => \N__5010\,
            lcout => \uart_frame_decoder_N_306_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
