------- ROM creada automaticamente por ppm2rom -----------
------- Felipe Machado -----------------------------------
------- Departamento de Tecnologia Electronica -----------
------- Universidad Rey Juan Carlos ----------------------
------- http://gtebim.es ---------------------------------
----------------------------------------------------------
--------Datos de la imagen -------------------------------
--- Fichero original    : dibujo.ppm 
--- Filas    : 60 
--- Columnas : 80 
----------------------------------------------------------
--------Codificacion de la memoria------------------------
--- Palabras de 9 bits
--- De cada palabra hay 3 bits para cada color : "RRRGGGBBB" 512 colores



------ Puertos -------------------------------------------
-- Entradas ----------------------------------------------
--    clk  :  senal de reloj
--    addr :  direccion de la memoria
-- Salidas  ----------------------------------------------
--    dout :  dato de 9 bits de la direccion addr (un ciclo despues)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;
entity ROM_RGB_9b_dibujo is
  port (
    clk  : in  std_logic;   -- reloj
    addr : in  std_logic_vector(13-1 downto 0);
    dout : out std_logic_vector(12-1 downto 0) 
  );
end ROM_RGB_9b_dibujo;


architecture BEHAVIORAL of ROM_RGB_9b_dibujo is
  signal addr_int  : natural range 0 to 2**13-1;
  type memostruct is array (natural range<>) of std_logic_vector(9-1 downto 0);
  constant filaimg : memostruct := (
     --"RRRGGGBBB"
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "000111111",
       "000111111",
       "000111111",
       "111111000",
       "111111000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "111111000",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111111000",
       "000111111",
       "000111111",
       "000111111",
       "111111000",
       "111111000",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111111111",
       "111111111",
       "111110000",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "111111111",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111110000",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111111111",
       "111111111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111111111",
       "111111111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111111111",
       "111111111",
       "111111111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "111111111",
       "111111111",
       "111111111",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111111111",
       "111111111",
       "111111111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "111111111",
       "111111111",
       "111111111",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111111111",
       "111111111",
       "111111111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "111111111",
       "111111111",
       "111111111",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111111111",
       "111111111",
       "111111111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "111111111",
       "111111111",
       "111111111",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "111111111",
       "111111111",
       "111111111",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "111111111",
       "111111111",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "111111111",
       "111111111",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "111111111",
       "111111111",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111000000",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "111111111",
       "111111111",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000111111",
       "000111111",
       "000111111",
       "111000110",
       "111000110",
       "111000110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000111111",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "000111111",
       "111000110",
       "111000110",
       "111000110",
       "000111111",
       "000111111",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "000111111",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "111111111",
       "111111111",
       "111111111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "111111111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "001000111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "001000111",
       "001000111",
       "001000111",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "111000110",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000111000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000",
       "000000000"
        );

begin

  addr_int <= TO_INTEGER(unsigned(addr));

  P_ROM: process (clk)
  begin
    if clk'event and clk='1' then
      dout <= filaimg(addr_int)(8 downto 6) & '0' & filaimg(addr_int)(5 downto 3) & '0' & filaimg(addr_int)(2 downto 0) & '0';
    end if;
  end process;

end BEHAVIORAL;

