-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     Mar 12 2019 01:42:22

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "Pc2Drone" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of Pc2Drone
entity Pc2Drone is
port (
    debug_state_output : out std_logic_vector(4 downto 0);
    uart_input : in std_logic;
    uart_data_rdy : out std_logic;
    debug_sinkdatavalid_output : out std_logic;
    uart_input_debug : out std_logic;
    frame_decoder_dv : out std_logic;
    clk_system : in std_logic);
end Pc2Drone;

-- Architecture of Pc2Drone
-- View name is \INTERFACE\
architecture \INTERFACE\ of Pc2Drone is

signal \N__5303\ : std_logic;
signal \N__5302\ : std_logic;
signal \N__5301\ : std_logic;
signal \N__5292\ : std_logic;
signal \N__5291\ : std_logic;
signal \N__5290\ : std_logic;
signal \N__5283\ : std_logic;
signal \N__5282\ : std_logic;
signal \N__5281\ : std_logic;
signal \N__5274\ : std_logic;
signal \N__5273\ : std_logic;
signal \N__5272\ : std_logic;
signal \N__5265\ : std_logic;
signal \N__5264\ : std_logic;
signal \N__5263\ : std_logic;
signal \N__5256\ : std_logic;
signal \N__5255\ : std_logic;
signal \N__5254\ : std_logic;
signal \N__5247\ : std_logic;
signal \N__5246\ : std_logic;
signal \N__5245\ : std_logic;
signal \N__5238\ : std_logic;
signal \N__5237\ : std_logic;
signal \N__5236\ : std_logic;
signal \N__5229\ : std_logic;
signal \N__5228\ : std_logic;
signal \N__5227\ : std_logic;
signal \N__5220\ : std_logic;
signal \N__5219\ : std_logic;
signal \N__5218\ : std_logic;
signal \N__5211\ : std_logic;
signal \N__5210\ : std_logic;
signal \N__5209\ : std_logic;
signal \N__5192\ : std_logic;
signal \N__5189\ : std_logic;
signal \N__5186\ : std_logic;
signal \N__5183\ : std_logic;
signal \N__5182\ : std_logic;
signal \N__5179\ : std_logic;
signal \N__5176\ : std_logic;
signal \N__5173\ : std_logic;
signal \N__5168\ : std_logic;
signal \N__5165\ : std_logic;
signal \N__5162\ : std_logic;
signal \N__5161\ : std_logic;
signal \N__5160\ : std_logic;
signal \N__5159\ : std_logic;
signal \N__5158\ : std_logic;
signal \N__5157\ : std_logic;
signal \N__5156\ : std_logic;
signal \N__5155\ : std_logic;
signal \N__5152\ : std_logic;
signal \N__5149\ : std_logic;
signal \N__5146\ : std_logic;
signal \N__5141\ : std_logic;
signal \N__5138\ : std_logic;
signal \N__5135\ : std_logic;
signal \N__5134\ : std_logic;
signal \N__5131\ : std_logic;
signal \N__5130\ : std_logic;
signal \N__5117\ : std_logic;
signal \N__5114\ : std_logic;
signal \N__5111\ : std_logic;
signal \N__5108\ : std_logic;
signal \N__5107\ : std_logic;
signal \N__5106\ : std_logic;
signal \N__5105\ : std_logic;
signal \N__5104\ : std_logic;
signal \N__5099\ : std_logic;
signal \N__5094\ : std_logic;
signal \N__5091\ : std_logic;
signal \N__5088\ : std_logic;
signal \N__5083\ : std_logic;
signal \N__5080\ : std_logic;
signal \N__5077\ : std_logic;
signal \N__5070\ : std_logic;
signal \N__5063\ : std_logic;
signal \N__5062\ : std_logic;
signal \N__5061\ : std_logic;
signal \N__5058\ : std_logic;
signal \N__5053\ : std_logic;
signal \N__5052\ : std_logic;
signal \N__5051\ : std_logic;
signal \N__5046\ : std_logic;
signal \N__5043\ : std_logic;
signal \N__5042\ : std_logic;
signal \N__5041\ : std_logic;
signal \N__5038\ : std_logic;
signal \N__5037\ : std_logic;
signal \N__5036\ : std_logic;
signal \N__5035\ : std_logic;
signal \N__5034\ : std_logic;
signal \N__5033\ : std_logic;
signal \N__5030\ : std_logic;
signal \N__5027\ : std_logic;
signal \N__5024\ : std_logic;
signal \N__5021\ : std_logic;
signal \N__5018\ : std_logic;
signal \N__5009\ : std_logic;
signal \N__5006\ : std_logic;
signal \N__4991\ : std_logic;
signal \N__4988\ : std_logic;
signal \N__4985\ : std_logic;
signal \N__4982\ : std_logic;
signal \N__4981\ : std_logic;
signal \N__4978\ : std_logic;
signal \N__4977\ : std_logic;
signal \N__4974\ : std_logic;
signal \N__4971\ : std_logic;
signal \N__4968\ : std_logic;
signal \N__4963\ : std_logic;
signal \N__4958\ : std_logic;
signal \N__4957\ : std_logic;
signal \N__4954\ : std_logic;
signal \N__4951\ : std_logic;
signal \N__4950\ : std_logic;
signal \N__4949\ : std_logic;
signal \N__4946\ : std_logic;
signal \N__4941\ : std_logic;
signal \N__4938\ : std_logic;
signal \N__4931\ : std_logic;
signal \N__4928\ : std_logic;
signal \N__4925\ : std_logic;
signal \N__4922\ : std_logic;
signal \N__4919\ : std_logic;
signal \N__4918\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4916\ : std_logic;
signal \N__4915\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4913\ : std_logic;
signal \N__4912\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4910\ : std_logic;
signal \N__4907\ : std_logic;
signal \N__4904\ : std_logic;
signal \N__4901\ : std_logic;
signal \N__4898\ : std_logic;
signal \N__4897\ : std_logic;
signal \N__4888\ : std_logic;
signal \N__4883\ : std_logic;
signal \N__4878\ : std_logic;
signal \N__4875\ : std_logic;
signal \N__4872\ : std_logic;
signal \N__4869\ : std_logic;
signal \N__4866\ : std_logic;
signal \N__4863\ : std_logic;
signal \N__4858\ : std_logic;
signal \N__4855\ : std_logic;
signal \N__4852\ : std_logic;
signal \N__4847\ : std_logic;
signal \N__4838\ : std_logic;
signal \N__4835\ : std_logic;
signal \N__4832\ : std_logic;
signal \N__4829\ : std_logic;
signal \N__4826\ : std_logic;
signal \N__4825\ : std_logic;
signal \N__4822\ : std_logic;
signal \N__4819\ : std_logic;
signal \N__4814\ : std_logic;
signal \N__4813\ : std_logic;
signal \N__4812\ : std_logic;
signal \N__4811\ : std_logic;
signal \N__4810\ : std_logic;
signal \N__4809\ : std_logic;
signal \N__4808\ : std_logic;
signal \N__4807\ : std_logic;
signal \N__4806\ : std_logic;
signal \N__4805\ : std_logic;
signal \N__4804\ : std_logic;
signal \N__4803\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4801\ : std_logic;
signal \N__4800\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4798\ : std_logic;
signal \N__4797\ : std_logic;
signal \N__4796\ : std_logic;
signal \N__4795\ : std_logic;
signal \N__4794\ : std_logic;
signal \N__4793\ : std_logic;
signal \N__4792\ : std_logic;
signal \N__4791\ : std_logic;
signal \N__4790\ : std_logic;
signal \N__4789\ : std_logic;
signal \N__4788\ : std_logic;
signal \N__4787\ : std_logic;
signal \N__4730\ : std_logic;
signal \N__4727\ : std_logic;
signal \N__4724\ : std_logic;
signal \N__4723\ : std_logic;
signal \N__4720\ : std_logic;
signal \N__4717\ : std_logic;
signal \N__4716\ : std_logic;
signal \N__4713\ : std_logic;
signal \N__4710\ : std_logic;
signal \N__4707\ : std_logic;
signal \N__4706\ : std_logic;
signal \N__4703\ : std_logic;
signal \N__4700\ : std_logic;
signal \N__4697\ : std_logic;
signal \N__4694\ : std_logic;
signal \N__4693\ : std_logic;
signal \N__4692\ : std_logic;
signal \N__4689\ : std_logic;
signal \N__4684\ : std_logic;
signal \N__4681\ : std_logic;
signal \N__4678\ : std_logic;
signal \N__4675\ : std_logic;
signal \N__4664\ : std_logic;
signal \N__4663\ : std_logic;
signal \N__4660\ : std_logic;
signal \N__4657\ : std_logic;
signal \N__4652\ : std_logic;
signal \N__4651\ : std_logic;
signal \N__4648\ : std_logic;
signal \N__4645\ : std_logic;
signal \N__4640\ : std_logic;
signal \N__4639\ : std_logic;
signal \N__4636\ : std_logic;
signal \N__4633\ : std_logic;
signal \N__4630\ : std_logic;
signal \N__4625\ : std_logic;
signal \N__4624\ : std_logic;
signal \N__4621\ : std_logic;
signal \N__4618\ : std_logic;
signal \N__4613\ : std_logic;
signal \N__4612\ : std_logic;
signal \N__4611\ : std_logic;
signal \N__4610\ : std_logic;
signal \N__4609\ : std_logic;
signal \N__4608\ : std_logic;
signal \N__4599\ : std_logic;
signal \N__4594\ : std_logic;
signal \N__4589\ : std_logic;
signal \N__4586\ : std_logic;
signal \N__4583\ : std_logic;
signal \N__4582\ : std_logic;
signal \N__4579\ : std_logic;
signal \N__4576\ : std_logic;
signal \N__4571\ : std_logic;
signal \N__4568\ : std_logic;
signal \N__4567\ : std_logic;
signal \N__4564\ : std_logic;
signal \N__4561\ : std_logic;
signal \N__4556\ : std_logic;
signal \N__4553\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4549\ : std_logic;
signal \N__4546\ : std_logic;
signal \N__4543\ : std_logic;
signal \N__4538\ : std_logic;
signal \N__4535\ : std_logic;
signal \N__4532\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4528\ : std_logic;
signal \N__4525\ : std_logic;
signal \N__4522\ : std_logic;
signal \N__4517\ : std_logic;
signal \N__4514\ : std_logic;
signal \N__4511\ : std_logic;
signal \N__4510\ : std_logic;
signal \N__4507\ : std_logic;
signal \N__4504\ : std_logic;
signal \N__4501\ : std_logic;
signal \N__4496\ : std_logic;
signal \N__4493\ : std_logic;
signal \N__4490\ : std_logic;
signal \N__4487\ : std_logic;
signal \N__4486\ : std_logic;
signal \N__4483\ : std_logic;
signal \N__4480\ : std_logic;
signal \N__4477\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4469\ : std_logic;
signal \N__4468\ : std_logic;
signal \N__4465\ : std_logic;
signal \N__4462\ : std_logic;
signal \N__4457\ : std_logic;
signal \N__4454\ : std_logic;
signal \N__4451\ : std_logic;
signal \N__4448\ : std_logic;
signal \N__4447\ : std_logic;
signal \N__4444\ : std_logic;
signal \N__4441\ : std_logic;
signal \N__4438\ : std_logic;
signal \N__4433\ : std_logic;
signal \N__4430\ : std_logic;
signal \N__4429\ : std_logic;
signal \N__4426\ : std_logic;
signal \N__4423\ : std_logic;
signal \N__4418\ : std_logic;
signal \N__4415\ : std_logic;
signal \N__4414\ : std_logic;
signal \N__4411\ : std_logic;
signal \N__4408\ : std_logic;
signal \N__4403\ : std_logic;
signal \N__4400\ : std_logic;
signal \N__4397\ : std_logic;
signal \N__4396\ : std_logic;
signal \N__4393\ : std_logic;
signal \N__4390\ : std_logic;
signal \N__4387\ : std_logic;
signal \N__4382\ : std_logic;
signal \N__4379\ : std_logic;
signal \N__4378\ : std_logic;
signal \N__4375\ : std_logic;
signal \N__4372\ : std_logic;
signal \N__4367\ : std_logic;
signal \N__4364\ : std_logic;
signal \N__4363\ : std_logic;
signal \N__4360\ : std_logic;
signal \N__4357\ : std_logic;
signal \N__4352\ : std_logic;
signal \N__4349\ : std_logic;
signal \N__4348\ : std_logic;
signal \N__4345\ : std_logic;
signal \N__4342\ : std_logic;
signal \N__4339\ : std_logic;
signal \N__4334\ : std_logic;
signal \N__4331\ : std_logic;
signal \N__4330\ : std_logic;
signal \N__4327\ : std_logic;
signal \N__4324\ : std_logic;
signal \N__4319\ : std_logic;
signal \N__4316\ : std_logic;
signal \N__4313\ : std_logic;
signal \N__4312\ : std_logic;
signal \N__4309\ : std_logic;
signal \N__4306\ : std_logic;
signal \N__4305\ : std_logic;
signal \N__4304\ : std_logic;
signal \N__4303\ : std_logic;
signal \N__4302\ : std_logic;
signal \N__4301\ : std_logic;
signal \N__4300\ : std_logic;
signal \N__4299\ : std_logic;
signal \N__4298\ : std_logic;
signal \N__4297\ : std_logic;
signal \N__4296\ : std_logic;
signal \N__4293\ : std_logic;
signal \N__4290\ : std_logic;
signal \N__4287\ : std_logic;
signal \N__4280\ : std_logic;
signal \N__4277\ : std_logic;
signal \N__4266\ : std_logic;
signal \N__4253\ : std_logic;
signal \N__4250\ : std_logic;
signal \N__4247\ : std_logic;
signal \N__4246\ : std_logic;
signal \N__4243\ : std_logic;
signal \N__4242\ : std_logic;
signal \N__4239\ : std_logic;
signal \N__4236\ : std_logic;
signal \N__4235\ : std_logic;
signal \N__4232\ : std_logic;
signal \N__4229\ : std_logic;
signal \N__4226\ : std_logic;
signal \N__4223\ : std_logic;
signal \N__4220\ : std_logic;
signal \N__4211\ : std_logic;
signal \N__4208\ : std_logic;
signal \N__4205\ : std_logic;
signal \N__4204\ : std_logic;
signal \N__4199\ : std_logic;
signal \N__4198\ : std_logic;
signal \N__4197\ : std_logic;
signal \N__4196\ : std_logic;
signal \N__4195\ : std_logic;
signal \N__4194\ : std_logic;
signal \N__4193\ : std_logic;
signal \N__4192\ : std_logic;
signal \N__4189\ : std_logic;
signal \N__4176\ : std_logic;
signal \N__4173\ : std_logic;
signal \N__4170\ : std_logic;
signal \N__4163\ : std_logic;
signal \N__4162\ : std_logic;
signal \N__4161\ : std_logic;
signal \N__4160\ : std_logic;
signal \N__4159\ : std_logic;
signal \N__4156\ : std_logic;
signal \N__4151\ : std_logic;
signal \N__4148\ : std_logic;
signal \N__4145\ : std_logic;
signal \N__4140\ : std_logic;
signal \N__4137\ : std_logic;
signal \N__4132\ : std_logic;
signal \N__4127\ : std_logic;
signal \N__4126\ : std_logic;
signal \N__4123\ : std_logic;
signal \N__4120\ : std_logic;
signal \N__4119\ : std_logic;
signal \N__4118\ : std_logic;
signal \N__4115\ : std_logic;
signal \N__4114\ : std_logic;
signal \N__4113\ : std_logic;
signal \N__4112\ : std_logic;
signal \N__4109\ : std_logic;
signal \N__4106\ : std_logic;
signal \N__4105\ : std_logic;
signal \N__4104\ : std_logic;
signal \N__4103\ : std_logic;
signal \N__4102\ : std_logic;
signal \N__4101\ : std_logic;
signal \N__4100\ : std_logic;
signal \N__4097\ : std_logic;
signal \N__4094\ : std_logic;
signal \N__4087\ : std_logic;
signal \N__4082\ : std_logic;
signal \N__4079\ : std_logic;
signal \N__4068\ : std_logic;
signal \N__4055\ : std_logic;
signal \N__4052\ : std_logic;
signal \N__4049\ : std_logic;
signal \N__4046\ : std_logic;
signal \N__4045\ : std_logic;
signal \N__4042\ : std_logic;
signal \N__4039\ : std_logic;
signal \N__4038\ : std_logic;
signal \N__4037\ : std_logic;
signal \N__4036\ : std_logic;
signal \N__4033\ : std_logic;
signal \N__4032\ : std_logic;
signal \N__4031\ : std_logic;
signal \N__4030\ : std_logic;
signal \N__4021\ : std_logic;
signal \N__4018\ : std_logic;
signal \N__4011\ : std_logic;
signal \N__4004\ : std_logic;
signal \N__4003\ : std_logic;
signal \N__4002\ : std_logic;
signal \N__3999\ : std_logic;
signal \N__3998\ : std_logic;
signal \N__3997\ : std_logic;
signal \N__3994\ : std_logic;
signal \N__3991\ : std_logic;
signal \N__3988\ : std_logic;
signal \N__3981\ : std_logic;
signal \N__3974\ : std_logic;
signal \N__3973\ : std_logic;
signal \N__3972\ : std_logic;
signal \N__3969\ : std_logic;
signal \N__3968\ : std_logic;
signal \N__3965\ : std_logic;
signal \N__3962\ : std_logic;
signal \N__3959\ : std_logic;
signal \N__3956\ : std_logic;
signal \N__3953\ : std_logic;
signal \N__3946\ : std_logic;
signal \N__3943\ : std_logic;
signal \N__3940\ : std_logic;
signal \N__3935\ : std_logic;
signal \N__3934\ : std_logic;
signal \N__3933\ : std_logic;
signal \N__3932\ : std_logic;
signal \N__3931\ : std_logic;
signal \N__3930\ : std_logic;
signal \N__3927\ : std_logic;
signal \N__3924\ : std_logic;
signal \N__3923\ : std_logic;
signal \N__3922\ : std_logic;
signal \N__3921\ : std_logic;
signal \N__3920\ : std_logic;
signal \N__3917\ : std_logic;
signal \N__3916\ : std_logic;
signal \N__3915\ : std_logic;
signal \N__3912\ : std_logic;
signal \N__3909\ : std_logic;
signal \N__3908\ : std_logic;
signal \N__3905\ : std_logic;
signal \N__3900\ : std_logic;
signal \N__3893\ : std_logic;
signal \N__3890\ : std_logic;
signal \N__3885\ : std_logic;
signal \N__3882\ : std_logic;
signal \N__3875\ : std_logic;
signal \N__3860\ : std_logic;
signal \N__3857\ : std_logic;
signal \N__3854\ : std_logic;
signal \N__3853\ : std_logic;
signal \N__3852\ : std_logic;
signal \N__3849\ : std_logic;
signal \N__3846\ : std_logic;
signal \N__3843\ : std_logic;
signal \N__3836\ : std_logic;
signal \N__3833\ : std_logic;
signal \N__3830\ : std_logic;
signal \N__3829\ : std_logic;
signal \N__3828\ : std_logic;
signal \N__3827\ : std_logic;
signal \N__3824\ : std_logic;
signal \N__3821\ : std_logic;
signal \N__3816\ : std_logic;
signal \N__3809\ : std_logic;
signal \N__3806\ : std_logic;
signal \N__3803\ : std_logic;
signal \N__3800\ : std_logic;
signal \N__3799\ : std_logic;
signal \N__3798\ : std_logic;
signal \N__3797\ : std_logic;
signal \N__3792\ : std_logic;
signal \N__3789\ : std_logic;
signal \N__3786\ : std_logic;
signal \N__3783\ : std_logic;
signal \N__3776\ : std_logic;
signal \N__3775\ : std_logic;
signal \N__3774\ : std_logic;
signal \N__3773\ : std_logic;
signal \N__3770\ : std_logic;
signal \N__3763\ : std_logic;
signal \N__3762\ : std_logic;
signal \N__3759\ : std_logic;
signal \N__3756\ : std_logic;
signal \N__3753\ : std_logic;
signal \N__3748\ : std_logic;
signal \N__3743\ : std_logic;
signal \N__3742\ : std_logic;
signal \N__3739\ : std_logic;
signal \N__3736\ : std_logic;
signal \N__3735\ : std_logic;
signal \N__3734\ : std_logic;
signal \N__3729\ : std_logic;
signal \N__3724\ : std_logic;
signal \N__3719\ : std_logic;
signal \N__3716\ : std_logic;
signal \N__3713\ : std_logic;
signal \N__3710\ : std_logic;
signal \N__3707\ : std_logic;
signal \N__3704\ : std_logic;
signal \N__3703\ : std_logic;
signal \N__3702\ : std_logic;
signal \N__3701\ : std_logic;
signal \N__3700\ : std_logic;
signal \N__3691\ : std_logic;
signal \N__3688\ : std_logic;
signal \N__3683\ : std_logic;
signal \N__3682\ : std_logic;
signal \N__3679\ : std_logic;
signal \N__3678\ : std_logic;
signal \N__3675\ : std_logic;
signal \N__3668\ : std_logic;
signal \N__3667\ : std_logic;
signal \N__3666\ : std_logic;
signal \N__3663\ : std_logic;
signal \N__3658\ : std_logic;
signal \N__3653\ : std_logic;
signal \N__3650\ : std_logic;
signal \N__3647\ : std_logic;
signal \N__3644\ : std_logic;
signal \N__3641\ : std_logic;
signal \N__3640\ : std_logic;
signal \N__3639\ : std_logic;
signal \N__3638\ : std_logic;
signal \N__3635\ : std_logic;
signal \N__3632\ : std_logic;
signal \N__3629\ : std_logic;
signal \N__3626\ : std_logic;
signal \N__3625\ : std_logic;
signal \N__3624\ : std_logic;
signal \N__3621\ : std_logic;
signal \N__3616\ : std_logic;
signal \N__3615\ : std_logic;
signal \N__3612\ : std_logic;
signal \N__3611\ : std_logic;
signal \N__3608\ : std_logic;
signal \N__3607\ : std_logic;
signal \N__3606\ : std_logic;
signal \N__3603\ : std_logic;
signal \N__3602\ : std_logic;
signal \N__3601\ : std_logic;
signal \N__3600\ : std_logic;
signal \N__3595\ : std_logic;
signal \N__3592\ : std_logic;
signal \N__3589\ : std_logic;
signal \N__3578\ : std_logic;
signal \N__3571\ : std_logic;
signal \N__3560\ : std_logic;
signal \N__3557\ : std_logic;
signal \N__3554\ : std_logic;
signal \N__3551\ : std_logic;
signal \N__3550\ : std_logic;
signal \N__3549\ : std_logic;
signal \N__3546\ : std_logic;
signal \N__3543\ : std_logic;
signal \N__3540\ : std_logic;
signal \N__3539\ : std_logic;
signal \N__3536\ : std_logic;
signal \N__3533\ : std_logic;
signal \N__3532\ : std_logic;
signal \N__3531\ : std_logic;
signal \N__3530\ : std_logic;
signal \N__3527\ : std_logic;
signal \N__3524\ : std_logic;
signal \N__3519\ : std_logic;
signal \N__3512\ : std_logic;
signal \N__3509\ : std_logic;
signal \N__3506\ : std_logic;
signal \N__3497\ : std_logic;
signal \N__3494\ : std_logic;
signal \N__3491\ : std_logic;
signal \N__3488\ : std_logic;
signal \N__3485\ : std_logic;
signal \N__3482\ : std_logic;
signal \N__3479\ : std_logic;
signal \N__3478\ : std_logic;
signal \N__3477\ : std_logic;
signal \N__3474\ : std_logic;
signal \N__3473\ : std_logic;
signal \N__3472\ : std_logic;
signal \N__3467\ : std_logic;
signal \N__3464\ : std_logic;
signal \N__3459\ : std_logic;
signal \N__3452\ : std_logic;
signal \N__3449\ : std_logic;
signal \N__3446\ : std_logic;
signal \N__3443\ : std_logic;
signal \N__3442\ : std_logic;
signal \N__3441\ : std_logic;
signal \N__3438\ : std_logic;
signal \N__3433\ : std_logic;
signal \N__3428\ : std_logic;
signal \N__3427\ : std_logic;
signal \N__3424\ : std_logic;
signal \N__3421\ : std_logic;
signal \N__3418\ : std_logic;
signal \N__3415\ : std_logic;
signal \N__3410\ : std_logic;
signal \N__3407\ : std_logic;
signal \N__3404\ : std_logic;
signal \N__3401\ : std_logic;
signal \N__3400\ : std_logic;
signal \N__3397\ : std_logic;
signal \N__3394\ : std_logic;
signal \N__3391\ : std_logic;
signal \N__3386\ : std_logic;
signal \N__3385\ : std_logic;
signal \N__3382\ : std_logic;
signal \N__3381\ : std_logic;
signal \N__3380\ : std_logic;
signal \N__3379\ : std_logic;
signal \N__3376\ : std_logic;
signal \N__3373\ : std_logic;
signal \N__3368\ : std_logic;
signal \N__3365\ : std_logic;
signal \N__3364\ : std_logic;
signal \N__3363\ : std_logic;
signal \N__3362\ : std_logic;
signal \N__3357\ : std_logic;
signal \N__3352\ : std_logic;
signal \N__3351\ : std_logic;
signal \N__3350\ : std_logic;
signal \N__3345\ : std_logic;
signal \N__3344\ : std_logic;
signal \N__3343\ : std_logic;
signal \N__3340\ : std_logic;
signal \N__3335\ : std_logic;
signal \N__3330\ : std_logic;
signal \N__3327\ : std_logic;
signal \N__3322\ : std_logic;
signal \N__3311\ : std_logic;
signal \N__3308\ : std_logic;
signal \N__3305\ : std_logic;
signal \N__3302\ : std_logic;
signal \N__3301\ : std_logic;
signal \N__3300\ : std_logic;
signal \N__3297\ : std_logic;
signal \N__3294\ : std_logic;
signal \N__3291\ : std_logic;
signal \N__3286\ : std_logic;
signal \N__3281\ : std_logic;
signal \N__3278\ : std_logic;
signal \N__3277\ : std_logic;
signal \N__3276\ : std_logic;
signal \N__3275\ : std_logic;
signal \N__3272\ : std_logic;
signal \N__3269\ : std_logic;
signal \N__3266\ : std_logic;
signal \N__3261\ : std_logic;
signal \N__3258\ : std_logic;
signal \N__3255\ : std_logic;
signal \N__3252\ : std_logic;
signal \N__3245\ : std_logic;
signal \N__3242\ : std_logic;
signal \N__3239\ : std_logic;
signal \N__3236\ : std_logic;
signal \N__3233\ : std_logic;
signal \N__3232\ : std_logic;
signal \N__3231\ : std_logic;
signal \N__3228\ : std_logic;
signal \N__3221\ : std_logic;
signal \N__3218\ : std_logic;
signal \N__3215\ : std_logic;
signal \N__3212\ : std_logic;
signal \N__3209\ : std_logic;
signal \N__3206\ : std_logic;
signal \N__3203\ : std_logic;
signal \N__3202\ : std_logic;
signal \N__3201\ : std_logic;
signal \N__3196\ : std_logic;
signal \N__3195\ : std_logic;
signal \N__3192\ : std_logic;
signal \N__3189\ : std_logic;
signal \N__3184\ : std_logic;
signal \N__3179\ : std_logic;
signal \N__3176\ : std_logic;
signal \N__3173\ : std_logic;
signal \N__3172\ : std_logic;
signal \N__3171\ : std_logic;
signal \N__3168\ : std_logic;
signal \N__3165\ : std_logic;
signal \N__3162\ : std_logic;
signal \N__3161\ : std_logic;
signal \N__3160\ : std_logic;
signal \N__3159\ : std_logic;
signal \N__3158\ : std_logic;
signal \N__3153\ : std_logic;
signal \N__3150\ : std_logic;
signal \N__3149\ : std_logic;
signal \N__3148\ : std_logic;
signal \N__3147\ : std_logic;
signal \N__3146\ : std_logic;
signal \N__3143\ : std_logic;
signal \N__3140\ : std_logic;
signal \N__3139\ : std_logic;
signal \N__3136\ : std_logic;
signal \N__3135\ : std_logic;
signal \N__3132\ : std_logic;
signal \N__3129\ : std_logic;
signal \N__3126\ : std_logic;
signal \N__3123\ : std_logic;
signal \N__3120\ : std_logic;
signal \N__3115\ : std_logic;
signal \N__3106\ : std_logic;
signal \N__3103\ : std_logic;
signal \N__3098\ : std_logic;
signal \N__3083\ : std_logic;
signal \N__3080\ : std_logic;
signal \N__3077\ : std_logic;
signal \N__3076\ : std_logic;
signal \N__3075\ : std_logic;
signal \N__3074\ : std_logic;
signal \N__3073\ : std_logic;
signal \N__3070\ : std_logic;
signal \N__3067\ : std_logic;
signal \N__3062\ : std_logic;
signal \N__3061\ : std_logic;
signal \N__3060\ : std_logic;
signal \N__3059\ : std_logic;
signal \N__3056\ : std_logic;
signal \N__3053\ : std_logic;
signal \N__3048\ : std_logic;
signal \N__3045\ : std_logic;
signal \N__3040\ : std_logic;
signal \N__3029\ : std_logic;
signal \N__3026\ : std_logic;
signal \N__3025\ : std_logic;
signal \N__3024\ : std_logic;
signal \N__3023\ : std_logic;
signal \N__3020\ : std_logic;
signal \N__3017\ : std_logic;
signal \N__3012\ : std_logic;
signal \N__3011\ : std_logic;
signal \N__3010\ : std_logic;
signal \N__3009\ : std_logic;
signal \N__3008\ : std_logic;
signal \N__3007\ : std_logic;
signal \N__3004\ : std_logic;
signal \N__2999\ : std_logic;
signal \N__2994\ : std_logic;
signal \N__2987\ : std_logic;
signal \N__2978\ : std_logic;
signal \N__2975\ : std_logic;
signal \N__2972\ : std_logic;
signal \N__2969\ : std_logic;
signal \N__2966\ : std_logic;
signal \N__2963\ : std_logic;
signal \N__2962\ : std_logic;
signal \N__2961\ : std_logic;
signal \N__2958\ : std_logic;
signal \N__2957\ : std_logic;
signal \N__2954\ : std_logic;
signal \N__2947\ : std_logic;
signal \N__2942\ : std_logic;
signal \N__2939\ : std_logic;
signal \N__2936\ : std_logic;
signal \N__2933\ : std_logic;
signal \N__2930\ : std_logic;
signal \N__2927\ : std_logic;
signal \N__2924\ : std_logic;
signal \N__2923\ : std_logic;
signal \N__2922\ : std_logic;
signal \N__2919\ : std_logic;
signal \N__2918\ : std_logic;
signal \N__2917\ : std_logic;
signal \N__2914\ : std_logic;
signal \N__2911\ : std_logic;
signal \N__2908\ : std_logic;
signal \N__2901\ : std_logic;
signal \N__2894\ : std_logic;
signal \N__2891\ : std_logic;
signal \N__2888\ : std_logic;
signal \N__2885\ : std_logic;
signal \N__2884\ : std_logic;
signal \N__2883\ : std_logic;
signal \N__2880\ : std_logic;
signal \N__2877\ : std_logic;
signal \N__2874\ : std_logic;
signal \N__2871\ : std_logic;
signal \N__2868\ : std_logic;
signal \N__2863\ : std_logic;
signal \N__2858\ : std_logic;
signal \N__2855\ : std_logic;
signal \N__2852\ : std_logic;
signal \N__2849\ : std_logic;
signal \N__2848\ : std_logic;
signal \N__2847\ : std_logic;
signal \N__2842\ : std_logic;
signal \N__2841\ : std_logic;
signal \N__2838\ : std_logic;
signal \N__2837\ : std_logic;
signal \N__2836\ : std_logic;
signal \N__2835\ : std_logic;
signal \N__2834\ : std_logic;
signal \N__2831\ : std_logic;
signal \N__2828\ : std_logic;
signal \N__2825\ : std_logic;
signal \N__2816\ : std_logic;
signal \N__2807\ : std_logic;
signal \N__2804\ : std_logic;
signal \N__2801\ : std_logic;
signal \N__2798\ : std_logic;
signal \N__2797\ : std_logic;
signal \N__2794\ : std_logic;
signal \N__2791\ : std_logic;
signal \N__2786\ : std_logic;
signal \N__2783\ : std_logic;
signal \N__2780\ : std_logic;
signal \N__2777\ : std_logic;
signal \N__2774\ : std_logic;
signal \N__2771\ : std_logic;
signal \N__2768\ : std_logic;
signal \N__2765\ : std_logic;
signal \N__2762\ : std_logic;
signal \N__2759\ : std_logic;
signal \N__2756\ : std_logic;
signal \N__2753\ : std_logic;
signal \N__2750\ : std_logic;
signal \N__2747\ : std_logic;
signal \N__2744\ : std_logic;
signal \N__2743\ : std_logic;
signal \N__2742\ : std_logic;
signal \N__2741\ : std_logic;
signal \N__2740\ : std_logic;
signal \N__2739\ : std_logic;
signal \N__2736\ : std_logic;
signal \N__2733\ : std_logic;
signal \N__2730\ : std_logic;
signal \N__2729\ : std_logic;
signal \N__2728\ : std_logic;
signal \N__2727\ : std_logic;
signal \N__2726\ : std_logic;
signal \N__2723\ : std_logic;
signal \N__2720\ : std_logic;
signal \N__2717\ : std_logic;
signal \N__2716\ : std_logic;
signal \N__2713\ : std_logic;
signal \N__2708\ : std_logic;
signal \N__2705\ : std_logic;
signal \N__2704\ : std_logic;
signal \N__2697\ : std_logic;
signal \N__2696\ : std_logic;
signal \N__2695\ : std_logic;
signal \N__2694\ : std_logic;
signal \N__2689\ : std_logic;
signal \N__2686\ : std_logic;
signal \N__2683\ : std_logic;
signal \N__2682\ : std_logic;
signal \N__2679\ : std_logic;
signal \N__2676\ : std_logic;
signal \N__2673\ : std_logic;
signal \N__2670\ : std_logic;
signal \N__2667\ : std_logic;
signal \N__2660\ : std_logic;
signal \N__2653\ : std_logic;
signal \N__2650\ : std_logic;
signal \N__2633\ : std_logic;
signal \N__2632\ : std_logic;
signal \N__2629\ : std_logic;
signal \N__2628\ : std_logic;
signal \N__2627\ : std_logic;
signal \N__2626\ : std_logic;
signal \N__2623\ : std_logic;
signal \N__2622\ : std_logic;
signal \N__2621\ : std_logic;
signal \N__2620\ : std_logic;
signal \N__2615\ : std_logic;
signal \N__2602\ : std_logic;
signal \N__2597\ : std_logic;
signal \N__2594\ : std_logic;
signal \N__2593\ : std_logic;
signal \N__2590\ : std_logic;
signal \N__2587\ : std_logic;
signal \N__2582\ : std_logic;
signal \N__2579\ : std_logic;
signal \N__2576\ : std_logic;
signal \N__2573\ : std_logic;
signal \N__2570\ : std_logic;
signal \N__2567\ : std_logic;
signal \N__2564\ : std_logic;
signal \N__2561\ : std_logic;
signal \N__2558\ : std_logic;
signal \N__2557\ : std_logic;
signal \N__2554\ : std_logic;
signal \N__2551\ : std_logic;
signal \N__2546\ : std_logic;
signal \N__2543\ : std_logic;
signal \N__2540\ : std_logic;
signal \N__2537\ : std_logic;
signal \N__2534\ : std_logic;
signal \N__2531\ : std_logic;
signal \N__2528\ : std_logic;
signal \N__2525\ : std_logic;
signal \N__2522\ : std_logic;
signal \N__2519\ : std_logic;
signal \N__2518\ : std_logic;
signal \N__2513\ : std_logic;
signal \N__2510\ : std_logic;
signal \N__2507\ : std_logic;
signal \N__2504\ : std_logic;
signal \N__2501\ : std_logic;
signal \N__2498\ : std_logic;
signal \N__2497\ : std_logic;
signal \N__2494\ : std_logic;
signal \N__2491\ : std_logic;
signal \N__2486\ : std_logic;
signal \N__2485\ : std_logic;
signal \N__2480\ : std_logic;
signal \N__2477\ : std_logic;
signal \N__2476\ : std_logic;
signal \N__2475\ : std_logic;
signal \N__2474\ : std_logic;
signal \N__2469\ : std_logic;
signal \N__2466\ : std_logic;
signal \N__2465\ : std_logic;
signal \N__2464\ : std_logic;
signal \N__2463\ : std_logic;
signal \N__2460\ : std_logic;
signal \N__2457\ : std_logic;
signal \N__2448\ : std_logic;
signal \N__2441\ : std_logic;
signal \N__2438\ : std_logic;
signal \N__2435\ : std_logic;
signal \N__2432\ : std_logic;
signal \N__2429\ : std_logic;
signal \N__2426\ : std_logic;
signal \N__2423\ : std_logic;
signal \N__2420\ : std_logic;
signal \N__2417\ : std_logic;
signal \N__2414\ : std_logic;
signal \N__2411\ : std_logic;
signal \N__2408\ : std_logic;
signal \N__2405\ : std_logic;
signal \N__2402\ : std_logic;
signal \N__2399\ : std_logic;
signal \N__2396\ : std_logic;
signal \N__2393\ : std_logic;
signal \N__2392\ : std_logic;
signal \N__2389\ : std_logic;
signal \N__2386\ : std_logic;
signal \N__2381\ : std_logic;
signal \N__2378\ : std_logic;
signal \N__2375\ : std_logic;
signal \N__2372\ : std_logic;
signal \N__2369\ : std_logic;
signal \N__2366\ : std_logic;
signal \N__2363\ : std_logic;
signal \N__2360\ : std_logic;
signal \N__2357\ : std_logic;
signal \N__2354\ : std_logic;
signal \N__2351\ : std_logic;
signal \N__2348\ : std_logic;
signal \N__2345\ : std_logic;
signal \N__2342\ : std_logic;
signal \N__2341\ : std_logic;
signal \N__2338\ : std_logic;
signal \N__2335\ : std_logic;
signal \N__2330\ : std_logic;
signal \N__2327\ : std_logic;
signal \N__2324\ : std_logic;
signal \N__2321\ : std_logic;
signal \N__2318\ : std_logic;
signal \N__2315\ : std_logic;
signal \N__2312\ : std_logic;
signal \N__2309\ : std_logic;
signal \N__2306\ : std_logic;
signal \N__2303\ : std_logic;
signal \N__2302\ : std_logic;
signal \N__2299\ : std_logic;
signal \N__2296\ : std_logic;
signal \N__2293\ : std_logic;
signal \N__2288\ : std_logic;
signal \N__2285\ : std_logic;
signal \N__2282\ : std_logic;
signal \N__2279\ : std_logic;
signal \N__2276\ : std_logic;
signal \N__2273\ : std_logic;
signal \N__2270\ : std_logic;
signal \N__2267\ : std_logic;
signal \N__2266\ : std_logic;
signal \N__2265\ : std_logic;
signal \N__2262\ : std_logic;
signal \N__2261\ : std_logic;
signal \N__2260\ : std_logic;
signal \N__2255\ : std_logic;
signal \N__2248\ : std_logic;
signal \N__2243\ : std_logic;
signal \N__2240\ : std_logic;
signal \N__2237\ : std_logic;
signal \N__2234\ : std_logic;
signal \N__2233\ : std_logic;
signal \N__2228\ : std_logic;
signal \N__2225\ : std_logic;
signal \N__2222\ : std_logic;
signal \N__2219\ : std_logic;
signal \N__2216\ : std_logic;
signal \N__2215\ : std_logic;
signal \N__2212\ : std_logic;
signal \N__2209\ : std_logic;
signal \N__2204\ : std_logic;
signal \N__2201\ : std_logic;
signal \N__2198\ : std_logic;
signal \N__2195\ : std_logic;
signal \N__2194\ : std_logic;
signal \N__2191\ : std_logic;
signal \N__2188\ : std_logic;
signal \N__2183\ : std_logic;
signal \N__2180\ : std_logic;
signal \N__2177\ : std_logic;
signal \N__2174\ : std_logic;
signal \N__2171\ : std_logic;
signal \N__2168\ : std_logic;
signal \N__2167\ : std_logic;
signal \N__2164\ : std_logic;
signal \N__2161\ : std_logic;
signal \N__2156\ : std_logic;
signal \N__2153\ : std_logic;
signal \N__2150\ : std_logic;
signal \N__2147\ : std_logic;
signal \N__2144\ : std_logic;
signal \N__2141\ : std_logic;
signal \N__2138\ : std_logic;
signal \N__2135\ : std_logic;
signal \N__2132\ : std_logic;
signal \N__2129\ : std_logic;
signal \N__2126\ : std_logic;
signal \N__2123\ : std_logic;
signal \N__2120\ : std_logic;
signal \N__2117\ : std_logic;
signal \N__2114\ : std_logic;
signal \N__2111\ : std_logic;
signal \N__2108\ : std_logic;
signal \N__2105\ : std_logic;
signal \N__2102\ : std_logic;
signal \N__2099\ : std_logic;
signal \N__2096\ : std_logic;
signal \N__2093\ : std_logic;
signal \N__2090\ : std_logic;
signal \N__2087\ : std_logic;
signal \N__2084\ : std_logic;
signal \N__2081\ : std_logic;
signal \N__2078\ : std_logic;
signal \N__2075\ : std_logic;
signal \N__2072\ : std_logic;
signal \N__2069\ : std_logic;
signal \N__2066\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \uart_frame_decoder.N_43_cascade_\ : std_logic;
signal \uart_frame_decoder.state_1_srsts_i_i_0_0_cascade_\ : std_logic;
signal \uart_frame_decoder_N_131_i\ : std_logic;
signal \uart_frame_decoder.state_1Z0Z_0\ : std_logic;
signal \uart_frame_decoder.state_1_srsts_0_i_1_1\ : std_logic;
signal \uart_frame_decoder.N_58_4\ : std_logic;
signal \uart_frame_decoder.N_58_4_cascade_\ : std_logic;
signal \uart_frame_decoder.N_32_i_1\ : std_logic;
signal \uart.state_0_sqmuxa_1_d_cascade_\ : std_logic;
signal \uart.m13_0_0_o2_2_cascade_\ : std_logic;
signal \uart.N_10_cascade_\ : std_logic;
signal \uart.data_Auxce_0_2_cascade_\ : std_logic;
signal \uart.data_Aux_esr_RNO_0Z0Z_2_cascade_\ : std_logic;
signal \uart.N_118_0\ : std_logic;
signal \uart_frame_decoder.state_1_srsts_0_i_a2_0_0_1Z0Z_2_cascade_\ : std_logic;
signal \uart_frame_decoder.N_49\ : std_logic;
signal \uart_frame_decoder.state_1Z0Z_1\ : std_logic;
signal \uart_frame_decoder_N_129_i\ : std_logic;
signal \uart_frame_decoder.state_1_srsts_i_i_a2_3_0Z0Z_0_cascade_\ : std_logic;
signal \uart_frame_decoder.N_67\ : std_logic;
signal \uart_frame_decoder.N_61\ : std_logic;
signal \uart_frame_decoder.N_67_cascade_\ : std_logic;
signal \uart_frame_decoder.state_1_srsts_0_i_a2_0_0_2\ : std_logic;
signal \uart.data_AuxZ0Z_0\ : std_logic;
signal uart_data_0 : std_logic;
signal uart_data_1 : std_logic;
signal \uart.data_AuxZ0Z_2\ : std_logic;
signal uart_data_2 : std_logic;
signal uart_data_3 : std_logic;
signal uart_data_4 : std_logic;
signal uart_data_5 : std_logic;
signal \uart.data_AuxZ0Z_6\ : std_logic;
signal uart_data_6 : std_logic;
signal \uart.data_AuxZ0Z_7\ : std_logic;
signal uart_data_7 : std_logic;
signal \uart.N_147_0_0_cascade_\ : std_logic;
signal \uart.g3_1_0_cascade_\ : std_logic;
signal \uart.g0_4_0\ : std_logic;
signal \uart.N_175_cascade_\ : std_logic;
signal \uart.data_Aux_esr_RNO_0Z0Z_0_cascade_\ : std_logic;
signal \uart.N_120_0\ : std_logic;
signal \uart.data_Auxce_0_0\ : std_logic;
signal \uart.data_Aux_esr_RNO_0Z0Z_1_cascade_\ : std_logic;
signal \uart.data_AuxZ0Z_1\ : std_logic;
signal \uart.N_119_0\ : std_logic;
signal \uart.data_Auxce_0_2\ : std_logic;
signal \uart.data_Aux_esr_RNO_0Z0Z_3_cascade_\ : std_logic;
signal \uart.data_Aux_esr_RNO_0Z0Z_4_cascade_\ : std_logic;
signal \uart.data_Auxce_0_4\ : std_logic;
signal \uart.N_113_0\ : std_logic;
signal \uart.N_133_0\ : std_logic;
signal \uart.stateZ0Z_0\ : std_logic;
signal \uart.N_175\ : std_logic;
signal \uart.data_Auxce_0_6_cascade_\ : std_logic;
signal \uart.N_114_0\ : std_logic;
signal \uart.data_Aux_esr_RNO_0Z0Z_5\ : std_logic;
signal \uart.data_AuxZ0Z_5\ : std_logic;
signal \uart.N_115_0\ : std_logic;
signal \uart.un4_timer_Count_1_c2_cascade_\ : std_logic;
signal \uart.state_srsts_0_a3_1_4_cascade_\ : std_logic;
signal \uart.timer_Count_fastZ0Z_4\ : std_logic;
signal \uart.timer_Count10lto4_0\ : std_logic;
signal \uart.timer_Count10lto4_0_cascade_\ : std_logic;
signal \uart.N_51_cascade_\ : std_logic;
signal \uart.N_146_0\ : std_logic;
signal \uart.data_14_1_cascade_\ : std_logic;
signal \uart.state_RNILS533Z0Z_4\ : std_logic;
signal \uart.state_RNILS533Z0Z_4_cascade_\ : std_logic;
signal \uart.state_1_sqmuxa_0\ : std_logic;
signal \uart.stateZ0Z_1\ : std_logic;
signal \uart.N_151\ : std_logic;
signal \uart.N_174\ : std_logic;
signal \uart.state_srsts_0_a3_2_0_4\ : std_logic;
signal \uart.state_1_sqmuxa\ : std_logic;
signal \uart.data_AuxZ0Z_3\ : std_logic;
signal \uart.N_117_0\ : std_logic;
signal \uart.data_AuxZ0Z_4\ : std_logic;
signal \uart.N_116_0\ : std_logic;
signal \uart.state_RNIAFHLZ0Z_4\ : std_logic;
signal \uart.timer_CountZ0Z_2\ : std_logic;
signal \uart.timer_Count_fastZ0Z_2\ : std_logic;
signal \reset_module_System.reset6_11_cascade_\ : std_logic;
signal \reset_module_System.reset6_19_cascade_\ : std_logic;
signal \uart.N_66\ : std_logic;
signal \uart.N_51\ : std_logic;
signal \uart.timer_Count_fastZ0Z_3\ : std_logic;
signal \uart.N_5\ : std_logic;
signal \uart.timer_Count_RNI3B101Z0Z_6\ : std_logic;
signal \uart.un4_timer_Count_1_c5\ : std_logic;
signal \uart.un1_state_2_0_a3_2\ : std_logic;
signal \uart.timer_CountZ0Z_0\ : std_logic;
signal \uart.timer_Count_RNI22NA1Z0Z_4\ : std_logic;
signal \uart.bit_CountZ0Z_0\ : std_logic;
signal \uart.bit_CountZ0Z_2\ : std_logic;
signal \uart.bit_CountZ0Z_1\ : std_logic;
signal \uart.g1_4_cascade_\ : std_logic;
signal \uart.g1_0\ : std_logic;
signal \uart.g1_3\ : std_logic;
signal \uart.stateZ0Z_2\ : std_logic;
signal \uart.un1_state_5\ : std_logic;
signal \uart.N_177\ : std_logic;
signal reset_system : std_logic;
signal \uart.N_28_mux\ : std_logic;
signal \uart.N_8_cascade_\ : std_logic;
signal \uart_frame_decoder.state_1Z0Z_4\ : std_logic;
signal \uart_frame_decoder.state_1Z0Z_5\ : std_logic;
signal \reset_module_System.reset6_3\ : std_logic;
signal \reset_module_System.reset6_14_cascade_\ : std_logic;
signal \reset_module_System.reset6_19\ : std_logic;
signal \reset_module_System.reset6_14\ : std_logic;
signal \reset_module_System.reset6_19_1\ : std_logic;
signal \reset_module_System.reset6_13\ : std_logic;
signal \uart.stateZ0Z_3\ : std_logic;
signal \uart.g3_0_0\ : std_logic;
signal \uart.timer_CountZ0Z_4\ : std_logic;
signal \uart.state_0_sqmuxa_1_d_0\ : std_logic;
signal \uart.timer_CountZ0Z_1\ : std_logic;
signal \uart.g3_cascade_\ : std_logic;
signal \uart.timer_CountZ0Z_6\ : std_logic;
signal \uart.N_167_0\ : std_logic;
signal \reset_module_System_reset_fast\ : std_logic;
signal \uart.g0_3_1\ : std_logic;
signal \uart.timer_CountZ0Z_3\ : std_logic;
signal \uart.timer_Count_4_repZ0Z1\ : std_logic;
signal \uart.timer_CountZ0Z_5\ : std_logic;
signal \uart.state_RNO_2Z0Z_3\ : std_logic;
signal \uart.un4_timer_Count_1_c2\ : std_logic;
signal \uart.timer_Count_2_repZ0Z1\ : std_logic;
signal \uart.state_RNI38F97Z0Z_2\ : std_logic;
signal \uart.timer_CountZ0Z_7\ : std_logic;
signal \uart.N_41\ : std_logic;
signal \uart.state_srsts_0_o4_0_a2_0_4\ : std_logic;
signal \uart_frame_decoder.uart_data_rdy_c_0\ : std_logic;
signal \uart_frame_decoder.state_1Z0Z_3\ : std_logic;
signal \uart_frame_decoder.state_1Z0Z_6\ : std_logic;
signal \uart_frame_decoder.state_1Z0Z_2\ : std_logic;
signal \uart_frame_decoder_N_130_i\ : std_logic;
signal \bfn_12_2_0_\ : std_logic;
signal \reset_module_System.countZ0Z_2\ : std_logic;
signal \reset_module_System.count_1_2\ : std_logic;
signal \reset_module_System.count_1_cry_1\ : std_logic;
signal \reset_module_System.countZ0Z_3\ : std_logic;
signal \reset_module_System.count_1_cry_2\ : std_logic;
signal \reset_module_System.countZ0Z_4\ : std_logic;
signal \reset_module_System.count_1_cry_3\ : std_logic;
signal \reset_module_System.countZ0Z_5\ : std_logic;
signal \reset_module_System.count_1_cry_4\ : std_logic;
signal \reset_module_System.countZ0Z_6\ : std_logic;
signal \reset_module_System.count_1_cry_5\ : std_logic;
signal \reset_module_System.countZ0Z_7\ : std_logic;
signal \reset_module_System.count_1_cry_6\ : std_logic;
signal \reset_module_System.countZ0Z_8\ : std_logic;
signal \reset_module_System.count_1_cry_7\ : std_logic;
signal \reset_module_System.count_1_cry_8\ : std_logic;
signal \reset_module_System.countZ0Z_9\ : std_logic;
signal \bfn_12_3_0_\ : std_logic;
signal \reset_module_System.countZ0Z_10\ : std_logic;
signal \reset_module_System.count_1_cry_9\ : std_logic;
signal \reset_module_System.countZ0Z_11\ : std_logic;
signal \reset_module_System.count_1_cry_10\ : std_logic;
signal \reset_module_System.countZ0Z_12\ : std_logic;
signal \reset_module_System.count_1_cry_11\ : std_logic;
signal \reset_module_System.count_1_cry_12\ : std_logic;
signal \reset_module_System.countZ0Z_14\ : std_logic;
signal \reset_module_System.count_1_cry_13\ : std_logic;
signal \reset_module_System.count_1_cry_14\ : std_logic;
signal \reset_module_System.countZ0Z_16\ : std_logic;
signal \reset_module_System.count_1_cry_15\ : std_logic;
signal \reset_module_System.count_1_cry_16\ : std_logic;
signal \reset_module_System.countZ0Z_17\ : std_logic;
signal \bfn_12_4_0_\ : std_logic;
signal \reset_module_System.countZ0Z_18\ : std_logic;
signal \reset_module_System.count_1_cry_17\ : std_logic;
signal \reset_module_System.count_1_cry_18\ : std_logic;
signal \reset_module_System.countZ0Z_20\ : std_logic;
signal \reset_module_System.count_1_cry_19\ : std_logic;
signal \reset_module_System.count_1_cry_20\ : std_logic;
signal uart_input_c : std_logic;
signal \uart.stateZ0Z_4\ : std_logic;
signal \uart.data_rdyc_0\ : std_logic;
signal \reset_module_System.countZ0Z_1\ : std_logic;
signal \reset_module_System.countZ0Z_0\ : std_logic;
signal \reset_module_System.count_1_1\ : std_logic;
signal uart_data_rdy_c : std_logic;
signal frame_decoder_dv_c : std_logic;
signal clk_system_c_g : std_logic;
signal \reset_module_System_reset_iso\ : std_logic;
signal \reset_module_System.countZ0Z_19\ : std_logic;
signal \reset_module_System.countZ0Z_15\ : std_logic;
signal \reset_module_System.countZ0Z_21\ : std_logic;
signal \reset_module_System.countZ0Z_13\ : std_logic;
signal \reset_module_System.reset6_15\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal clk_system_wire : std_logic;
signal debug_state_output_wire : std_logic_vector(4 downto 0);
signal uart_data_rdy_wire : std_logic;
signal debug_sinkdatavalid_output_wire : std_logic;
signal frame_decoder_dv_wire : std_logic;
signal uart_input_wire : std_logic;
signal uart_input_debug_wire : std_logic;

begin
    clk_system_wire <= clk_system;
    debug_state_output <= debug_state_output_wire;
    uart_data_rdy <= uart_data_rdy_wire;
    debug_sinkdatavalid_output <= debug_sinkdatavalid_output_wire;
    frame_decoder_dv <= frame_decoder_dv_wire;
    uart_input_wire <= uart_input;
    uart_input_debug <= uart_input_debug_wire;

    \clk_system_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__5301\,
            GLOBALBUFFEROUTPUT => clk_system_c_g
        );

    \clk_system_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5303\,
            DIN => \N__5302\,
            DOUT => \N__5301\,
            PACKAGEPIN => clk_system_wire
        );

    \clk_system_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5303\,
            PADOUT => \N__5302\,
            PADIN => \N__5301\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \debug_state_output_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5292\,
            DIN => \N__5291\,
            DOUT => \N__5290\,
            PACKAGEPIN => debug_state_output_wire(4)
        );

    \debug_state_output_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5292\,
            PADOUT => \N__5291\,
            PADIN => \N__5290\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \debug_state_output_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5283\,
            DIN => \N__5282\,
            DOUT => \N__5281\,
            PACKAGEPIN => debug_state_output_wire(1)
        );

    \debug_state_output_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5283\,
            PADOUT => \N__5282\,
            PADIN => \N__5281\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3719\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \uart_data_rdy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5274\,
            DIN => \N__5273\,
            DOUT => \N__5272\,
            PACKAGEPIN => uart_data_rdy_wire
        );

    \uart_data_rdy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5274\,
            PADOUT => \N__5273\,
            PADIN => \N__5272\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4922\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \debug_state_output_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5265\,
            DIN => \N__5264\,
            DOUT => \N__5263\,
            PACKAGEPIN => debug_state_output_wire(3)
        );

    \debug_state_output_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5265\,
            PADOUT => \N__5264\,
            PADIN => \N__5263\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \debug_sinkdatavalid_output_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5256\,
            DIN => \N__5255\,
            DOUT => \N__5254\,
            PACKAGEPIN => debug_sinkdatavalid_output_wire
        );

    \debug_sinkdatavalid_output_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5256\,
            PADOUT => \N__5255\,
            PADIN => \N__5254\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4918\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \frame_decoder_dv_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5247\,
            DIN => \N__5246\,
            DOUT => \N__5245\,
            PACKAGEPIN => frame_decoder_dv_wire
        );

    \frame_decoder_dv_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5247\,
            PADOUT => \N__5246\,
            PADIN => \N__5245\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4838\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \uart_input_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5238\,
            DIN => \N__5237\,
            DOUT => \N__5236\,
            PACKAGEPIN => uart_input_wire
        );

    \uart_input_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5238\,
            PADOUT => \N__5237\,
            PADIN => \N__5236\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => uart_input_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \debug_state_output_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5229\,
            DIN => \N__5228\,
            DOUT => \N__5227\,
            PACKAGEPIN => debug_state_output_wire(0)
        );

    \debug_state_output_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5229\,
            PADOUT => \N__5228\,
            PADIN => \N__5227\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2243\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \debug_state_output_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5220\,
            DIN => \N__5219\,
            DOUT => \N__5218\,
            PACKAGEPIN => debug_state_output_wire(2)
        );

    \debug_state_output_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5220\,
            PADOUT => \N__5219\,
            PADIN => \N__5218\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2096\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \uart_input_debug_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5211\,
            DIN => \N__5210\,
            DOUT => \N__5209\,
            PACKAGEPIN => uart_input_debug_wire
        );

    \uart_input_debug_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5211\,
            PADOUT => \N__5210\,
            PADIN => \N__5209\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5130\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__1217\ : InMux
    port map (
            O => \N__5192\,
            I => \reset_module_System.count_1_cry_18\
        );

    \I__1216\ : CascadeMux
    port map (
            O => \N__5189\,
            I => \N__5186\
        );

    \I__1215\ : InMux
    port map (
            O => \N__5186\,
            I => \N__5183\
        );

    \I__1214\ : LocalMux
    port map (
            O => \N__5183\,
            I => \N__5179\
        );

    \I__1213\ : InMux
    port map (
            O => \N__5182\,
            I => \N__5176\
        );

    \I__1212\ : Span4Mux_s3_v
    port map (
            O => \N__5179\,
            I => \N__5173\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__5176\,
            I => \reset_module_System.countZ0Z_20\
        );

    \I__1210\ : Odrv4
    port map (
            O => \N__5173\,
            I => \reset_module_System.countZ0Z_20\
        );

    \I__1209\ : InMux
    port map (
            O => \N__5168\,
            I => \reset_module_System.count_1_cry_19\
        );

    \I__1208\ : InMux
    port map (
            O => \N__5165\,
            I => \reset_module_System.count_1_cry_20\
        );

    \I__1207\ : InMux
    port map (
            O => \N__5162\,
            I => \N__5152\
        );

    \I__1206\ : InMux
    port map (
            O => \N__5161\,
            I => \N__5149\
        );

    \I__1205\ : InMux
    port map (
            O => \N__5160\,
            I => \N__5146\
        );

    \I__1204\ : InMux
    port map (
            O => \N__5159\,
            I => \N__5141\
        );

    \I__1203\ : InMux
    port map (
            O => \N__5158\,
            I => \N__5141\
        );

    \I__1202\ : InMux
    port map (
            O => \N__5157\,
            I => \N__5138\
        );

    \I__1201\ : InMux
    port map (
            O => \N__5156\,
            I => \N__5135\
        );

    \I__1200\ : InMux
    port map (
            O => \N__5155\,
            I => \N__5131\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__5152\,
            I => \N__5117\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__5149\,
            I => \N__5117\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__5146\,
            I => \N__5117\
        );

    \I__1196\ : LocalMux
    port map (
            O => \N__5141\,
            I => \N__5117\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__5138\,
            I => \N__5117\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__5135\,
            I => \N__5117\
        );

    \I__1193\ : InMux
    port map (
            O => \N__5134\,
            I => \N__5114\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__5131\,
            I => \N__5111\
        );

    \I__1191\ : IoInMux
    port map (
            O => \N__5130\,
            I => \N__5108\
        );

    \I__1190\ : Span4Mux_v
    port map (
            O => \N__5117\,
            I => \N__5099\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__5114\,
            I => \N__5099\
        );

    \I__1188\ : Span4Mux_v
    port map (
            O => \N__5111\,
            I => \N__5094\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__5108\,
            I => \N__5094\
        );

    \I__1186\ : InMux
    port map (
            O => \N__5107\,
            I => \N__5091\
        );

    \I__1185\ : InMux
    port map (
            O => \N__5106\,
            I => \N__5088\
        );

    \I__1184\ : InMux
    port map (
            O => \N__5105\,
            I => \N__5083\
        );

    \I__1183\ : InMux
    port map (
            O => \N__5104\,
            I => \N__5083\
        );

    \I__1182\ : IoSpan4Mux
    port map (
            O => \N__5099\,
            I => \N__5080\
        );

    \I__1181\ : IoSpan4Mux
    port map (
            O => \N__5094\,
            I => \N__5077\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__5091\,
            I => \N__5070\
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__5088\,
            I => \N__5070\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__5083\,
            I => \N__5070\
        );

    \I__1177\ : Odrv4
    port map (
            O => \N__5080\,
            I => uart_input_c
        );

    \I__1176\ : Odrv4
    port map (
            O => \N__5077\,
            I => uart_input_c
        );

    \I__1175\ : Odrv12
    port map (
            O => \N__5070\,
            I => uart_input_c
        );

    \I__1174\ : InMux
    port map (
            O => \N__5063\,
            I => \N__5058\
        );

    \I__1173\ : InMux
    port map (
            O => \N__5062\,
            I => \N__5053\
        );

    \I__1172\ : InMux
    port map (
            O => \N__5061\,
            I => \N__5053\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__5058\,
            I => \N__5046\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__5053\,
            I => \N__5046\
        );

    \I__1169\ : InMux
    port map (
            O => \N__5052\,
            I => \N__5043\
        );

    \I__1168\ : InMux
    port map (
            O => \N__5051\,
            I => \N__5038\
        );

    \I__1167\ : Span4Mux_s3_v
    port map (
            O => \N__5046\,
            I => \N__5030\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__5043\,
            I => \N__5027\
        );

    \I__1165\ : InMux
    port map (
            O => \N__5042\,
            I => \N__5024\
        );

    \I__1164\ : InMux
    port map (
            O => \N__5041\,
            I => \N__5021\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__5038\,
            I => \N__5018\
        );

    \I__1162\ : InMux
    port map (
            O => \N__5037\,
            I => \N__5009\
        );

    \I__1161\ : InMux
    port map (
            O => \N__5036\,
            I => \N__5009\
        );

    \I__1160\ : InMux
    port map (
            O => \N__5035\,
            I => \N__5009\
        );

    \I__1159\ : InMux
    port map (
            O => \N__5034\,
            I => \N__5009\
        );

    \I__1158\ : InMux
    port map (
            O => \N__5033\,
            I => \N__5006\
        );

    \I__1157\ : Odrv4
    port map (
            O => \N__5030\,
            I => \uart.stateZ0Z_4\
        );

    \I__1156\ : Odrv4
    port map (
            O => \N__5027\,
            I => \uart.stateZ0Z_4\
        );

    \I__1155\ : LocalMux
    port map (
            O => \N__5024\,
            I => \uart.stateZ0Z_4\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__5021\,
            I => \uart.stateZ0Z_4\
        );

    \I__1153\ : Odrv4
    port map (
            O => \N__5018\,
            I => \uart.stateZ0Z_4\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__5009\,
            I => \uart.stateZ0Z_4\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__5006\,
            I => \uart.stateZ0Z_4\
        );

    \I__1150\ : CascadeMux
    port map (
            O => \N__4991\,
            I => \N__4988\
        );

    \I__1149\ : InMux
    port map (
            O => \N__4988\,
            I => \N__4985\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__4985\,
            I => \uart.data_rdyc_0\
        );

    \I__1147\ : CascadeMux
    port map (
            O => \N__4982\,
            I => \N__4978\
        );

    \I__1146\ : InMux
    port map (
            O => \N__4981\,
            I => \N__4974\
        );

    \I__1145\ : InMux
    port map (
            O => \N__4978\,
            I => \N__4971\
        );

    \I__1144\ : InMux
    port map (
            O => \N__4977\,
            I => \N__4968\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__4974\,
            I => \N__4963\
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__4971\,
            I => \N__4963\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__4968\,
            I => \reset_module_System.countZ0Z_1\
        );

    \I__1140\ : Odrv4
    port map (
            O => \N__4963\,
            I => \reset_module_System.countZ0Z_1\
        );

    \I__1139\ : InMux
    port map (
            O => \N__4958\,
            I => \N__4954\
        );

    \I__1138\ : CascadeMux
    port map (
            O => \N__4957\,
            I => \N__4951\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__4954\,
            I => \N__4946\
        );

    \I__1136\ : InMux
    port map (
            O => \N__4951\,
            I => \N__4941\
        );

    \I__1135\ : InMux
    port map (
            O => \N__4950\,
            I => \N__4941\
        );

    \I__1134\ : InMux
    port map (
            O => \N__4949\,
            I => \N__4938\
        );

    \I__1133\ : Odrv4
    port map (
            O => \N__4946\,
            I => \reset_module_System.countZ0Z_0\
        );

    \I__1132\ : LocalMux
    port map (
            O => \N__4941\,
            I => \reset_module_System.countZ0Z_0\
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__4938\,
            I => \reset_module_System.countZ0Z_0\
        );

    \I__1130\ : InMux
    port map (
            O => \N__4931\,
            I => \N__4928\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__4928\,
            I => \N__4925\
        );

    \I__1128\ : Odrv4
    port map (
            O => \N__4925\,
            I => \reset_module_System.count_1_1\
        );

    \I__1127\ : IoInMux
    port map (
            O => \N__4922\,
            I => \N__4919\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__4919\,
            I => \N__4907\
        );

    \I__1125\ : IoInMux
    port map (
            O => \N__4918\,
            I => \N__4904\
        );

    \I__1124\ : CascadeMux
    port map (
            O => \N__4917\,
            I => \N__4901\
        );

    \I__1123\ : InMux
    port map (
            O => \N__4916\,
            I => \N__4898\
        );

    \I__1122\ : InMux
    port map (
            O => \N__4915\,
            I => \N__4888\
        );

    \I__1121\ : InMux
    port map (
            O => \N__4914\,
            I => \N__4888\
        );

    \I__1120\ : InMux
    port map (
            O => \N__4913\,
            I => \N__4888\
        );

    \I__1119\ : InMux
    port map (
            O => \N__4912\,
            I => \N__4888\
        );

    \I__1118\ : InMux
    port map (
            O => \N__4911\,
            I => \N__4883\
        );

    \I__1117\ : InMux
    port map (
            O => \N__4910\,
            I => \N__4883\
        );

    \I__1116\ : IoSpan4Mux
    port map (
            O => \N__4907\,
            I => \N__4878\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__4904\,
            I => \N__4878\
        );

    \I__1114\ : InMux
    port map (
            O => \N__4901\,
            I => \N__4875\
        );

    \I__1113\ : LocalMux
    port map (
            O => \N__4898\,
            I => \N__4872\
        );

    \I__1112\ : InMux
    port map (
            O => \N__4897\,
            I => \N__4869\
        );

    \I__1111\ : LocalMux
    port map (
            O => \N__4888\,
            I => \N__4866\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__4883\,
            I => \N__4863\
        );

    \I__1109\ : IoSpan4Mux
    port map (
            O => \N__4878\,
            I => \N__4858\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__4875\,
            I => \N__4858\
        );

    \I__1107\ : Span4Mux_s3_v
    port map (
            O => \N__4872\,
            I => \N__4855\
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__4869\,
            I => \N__4852\
        );

    \I__1105\ : Span4Mux_h
    port map (
            O => \N__4866\,
            I => \N__4847\
        );

    \I__1104\ : Span4Mux_h
    port map (
            O => \N__4863\,
            I => \N__4847\
        );

    \I__1103\ : Odrv4
    port map (
            O => \N__4858\,
            I => uart_data_rdy_c
        );

    \I__1102\ : Odrv4
    port map (
            O => \N__4855\,
            I => uart_data_rdy_c
        );

    \I__1101\ : Odrv4
    port map (
            O => \N__4852\,
            I => uart_data_rdy_c
        );

    \I__1100\ : Odrv4
    port map (
            O => \N__4847\,
            I => uart_data_rdy_c
        );

    \I__1099\ : IoInMux
    port map (
            O => \N__4838\,
            I => \N__4835\
        );

    \I__1098\ : LocalMux
    port map (
            O => \N__4835\,
            I => \N__4832\
        );

    \I__1097\ : IoSpan4Mux
    port map (
            O => \N__4832\,
            I => \N__4829\
        );

    \I__1096\ : Span4Mux_s2_v
    port map (
            O => \N__4829\,
            I => \N__4826\
        );

    \I__1095\ : Span4Mux_h
    port map (
            O => \N__4826\,
            I => \N__4822\
        );

    \I__1094\ : InMux
    port map (
            O => \N__4825\,
            I => \N__4819\
        );

    \I__1093\ : Odrv4
    port map (
            O => \N__4822\,
            I => frame_decoder_dv_c
        );

    \I__1092\ : LocalMux
    port map (
            O => \N__4819\,
            I => frame_decoder_dv_c
        );

    \I__1091\ : ClkMux
    port map (
            O => \N__4814\,
            I => \N__4730\
        );

    \I__1090\ : ClkMux
    port map (
            O => \N__4813\,
            I => \N__4730\
        );

    \I__1089\ : ClkMux
    port map (
            O => \N__4812\,
            I => \N__4730\
        );

    \I__1088\ : ClkMux
    port map (
            O => \N__4811\,
            I => \N__4730\
        );

    \I__1087\ : ClkMux
    port map (
            O => \N__4810\,
            I => \N__4730\
        );

    \I__1086\ : ClkMux
    port map (
            O => \N__4809\,
            I => \N__4730\
        );

    \I__1085\ : ClkMux
    port map (
            O => \N__4808\,
            I => \N__4730\
        );

    \I__1084\ : ClkMux
    port map (
            O => \N__4807\,
            I => \N__4730\
        );

    \I__1083\ : ClkMux
    port map (
            O => \N__4806\,
            I => \N__4730\
        );

    \I__1082\ : ClkMux
    port map (
            O => \N__4805\,
            I => \N__4730\
        );

    \I__1081\ : ClkMux
    port map (
            O => \N__4804\,
            I => \N__4730\
        );

    \I__1080\ : ClkMux
    port map (
            O => \N__4803\,
            I => \N__4730\
        );

    \I__1079\ : ClkMux
    port map (
            O => \N__4802\,
            I => \N__4730\
        );

    \I__1078\ : ClkMux
    port map (
            O => \N__4801\,
            I => \N__4730\
        );

    \I__1077\ : ClkMux
    port map (
            O => \N__4800\,
            I => \N__4730\
        );

    \I__1076\ : ClkMux
    port map (
            O => \N__4799\,
            I => \N__4730\
        );

    \I__1075\ : ClkMux
    port map (
            O => \N__4798\,
            I => \N__4730\
        );

    \I__1074\ : ClkMux
    port map (
            O => \N__4797\,
            I => \N__4730\
        );

    \I__1073\ : ClkMux
    port map (
            O => \N__4796\,
            I => \N__4730\
        );

    \I__1072\ : ClkMux
    port map (
            O => \N__4795\,
            I => \N__4730\
        );

    \I__1071\ : ClkMux
    port map (
            O => \N__4794\,
            I => \N__4730\
        );

    \I__1070\ : ClkMux
    port map (
            O => \N__4793\,
            I => \N__4730\
        );

    \I__1069\ : ClkMux
    port map (
            O => \N__4792\,
            I => \N__4730\
        );

    \I__1068\ : ClkMux
    port map (
            O => \N__4791\,
            I => \N__4730\
        );

    \I__1067\ : ClkMux
    port map (
            O => \N__4790\,
            I => \N__4730\
        );

    \I__1066\ : ClkMux
    port map (
            O => \N__4789\,
            I => \N__4730\
        );

    \I__1065\ : ClkMux
    port map (
            O => \N__4788\,
            I => \N__4730\
        );

    \I__1064\ : ClkMux
    port map (
            O => \N__4787\,
            I => \N__4730\
        );

    \I__1063\ : GlobalMux
    port map (
            O => \N__4730\,
            I => \N__4727\
        );

    \I__1062\ : gio2CtrlBuf
    port map (
            O => \N__4727\,
            I => clk_system_c_g
        );

    \I__1061\ : SRMux
    port map (
            O => \N__4724\,
            I => \N__4720\
        );

    \I__1060\ : SRMux
    port map (
            O => \N__4723\,
            I => \N__4717\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__4720\,
            I => \N__4713\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__4717\,
            I => \N__4710\
        );

    \I__1057\ : SRMux
    port map (
            O => \N__4716\,
            I => \N__4707\
        );

    \I__1056\ : Span4Mux_v
    port map (
            O => \N__4713\,
            I => \N__4703\
        );

    \I__1055\ : Span4Mux_v
    port map (
            O => \N__4710\,
            I => \N__4700\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__4707\,
            I => \N__4697\
        );

    \I__1053\ : SRMux
    port map (
            O => \N__4706\,
            I => \N__4694\
        );

    \I__1052\ : Span4Mux_h
    port map (
            O => \N__4703\,
            I => \N__4689\
        );

    \I__1051\ : Span4Mux_s1_v
    port map (
            O => \N__4700\,
            I => \N__4684\
        );

    \I__1050\ : Span4Mux_v
    port map (
            O => \N__4697\,
            I => \N__4684\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__4694\,
            I => \N__4681\
        );

    \I__1048\ : SRMux
    port map (
            O => \N__4693\,
            I => \N__4678\
        );

    \I__1047\ : InMux
    port map (
            O => \N__4692\,
            I => \N__4675\
        );

    \I__1046\ : Odrv4
    port map (
            O => \N__4689\,
            I => \reset_module_System_reset_iso\
        );

    \I__1045\ : Odrv4
    port map (
            O => \N__4684\,
            I => \reset_module_System_reset_iso\
        );

    \I__1044\ : Odrv12
    port map (
            O => \N__4681\,
            I => \reset_module_System_reset_iso\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__4678\,
            I => \reset_module_System_reset_iso\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__4675\,
            I => \reset_module_System_reset_iso\
        );

    \I__1041\ : InMux
    port map (
            O => \N__4664\,
            I => \N__4660\
        );

    \I__1040\ : InMux
    port map (
            O => \N__4663\,
            I => \N__4657\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__4660\,
            I => \reset_module_System.countZ0Z_19\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__4657\,
            I => \reset_module_System.countZ0Z_19\
        );

    \I__1037\ : InMux
    port map (
            O => \N__4652\,
            I => \N__4648\
        );

    \I__1036\ : InMux
    port map (
            O => \N__4651\,
            I => \N__4645\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__4648\,
            I => \reset_module_System.countZ0Z_15\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__4645\,
            I => \reset_module_System.countZ0Z_15\
        );

    \I__1033\ : CascadeMux
    port map (
            O => \N__4640\,
            I => \N__4636\
        );

    \I__1032\ : InMux
    port map (
            O => \N__4639\,
            I => \N__4633\
        );

    \I__1031\ : InMux
    port map (
            O => \N__4636\,
            I => \N__4630\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__4633\,
            I => \reset_module_System.countZ0Z_21\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__4630\,
            I => \reset_module_System.countZ0Z_21\
        );

    \I__1028\ : InMux
    port map (
            O => \N__4625\,
            I => \N__4621\
        );

    \I__1027\ : InMux
    port map (
            O => \N__4624\,
            I => \N__4618\
        );

    \I__1026\ : LocalMux
    port map (
            O => \N__4621\,
            I => \reset_module_System.countZ0Z_13\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__4618\,
            I => \reset_module_System.countZ0Z_13\
        );

    \I__1024\ : InMux
    port map (
            O => \N__4613\,
            I => \N__4599\
        );

    \I__1023\ : InMux
    port map (
            O => \N__4612\,
            I => \N__4599\
        );

    \I__1022\ : InMux
    port map (
            O => \N__4611\,
            I => \N__4599\
        );

    \I__1021\ : InMux
    port map (
            O => \N__4610\,
            I => \N__4599\
        );

    \I__1020\ : InMux
    port map (
            O => \N__4609\,
            I => \N__4594\
        );

    \I__1019\ : InMux
    port map (
            O => \N__4608\,
            I => \N__4594\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__4599\,
            I => \N__4589\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__4594\,
            I => \N__4589\
        );

    \I__1016\ : Span4Mux_h
    port map (
            O => \N__4589\,
            I => \N__4586\
        );

    \I__1015\ : Odrv4
    port map (
            O => \N__4586\,
            I => \reset_module_System.reset6_15\
        );

    \I__1014\ : InMux
    port map (
            O => \N__4583\,
            I => \N__4579\
        );

    \I__1013\ : InMux
    port map (
            O => \N__4582\,
            I => \N__4576\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__4579\,
            I => \reset_module_System.countZ0Z_11\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__4576\,
            I => \reset_module_System.countZ0Z_11\
        );

    \I__1010\ : InMux
    port map (
            O => \N__4571\,
            I => \reset_module_System.count_1_cry_10\
        );

    \I__1009\ : InMux
    port map (
            O => \N__4568\,
            I => \N__4564\
        );

    \I__1008\ : InMux
    port map (
            O => \N__4567\,
            I => \N__4561\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__4564\,
            I => \reset_module_System.countZ0Z_12\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__4561\,
            I => \reset_module_System.countZ0Z_12\
        );

    \I__1005\ : InMux
    port map (
            O => \N__4556\,
            I => \reset_module_System.count_1_cry_11\
        );

    \I__1004\ : InMux
    port map (
            O => \N__4553\,
            I => \reset_module_System.count_1_cry_12\
        );

    \I__1003\ : InMux
    port map (
            O => \N__4550\,
            I => \N__4546\
        );

    \I__1002\ : InMux
    port map (
            O => \N__4549\,
            I => \N__4543\
        );

    \I__1001\ : LocalMux
    port map (
            O => \N__4546\,
            I => \reset_module_System.countZ0Z_14\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__4543\,
            I => \reset_module_System.countZ0Z_14\
        );

    \I__999\ : InMux
    port map (
            O => \N__4538\,
            I => \reset_module_System.count_1_cry_13\
        );

    \I__998\ : InMux
    port map (
            O => \N__4535\,
            I => \reset_module_System.count_1_cry_14\
        );

    \I__997\ : InMux
    port map (
            O => \N__4532\,
            I => \N__4529\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__4529\,
            I => \N__4525\
        );

    \I__995\ : InMux
    port map (
            O => \N__4528\,
            I => \N__4522\
        );

    \I__994\ : Odrv4
    port map (
            O => \N__4525\,
            I => \reset_module_System.countZ0Z_16\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__4522\,
            I => \reset_module_System.countZ0Z_16\
        );

    \I__992\ : InMux
    port map (
            O => \N__4517\,
            I => \reset_module_System.count_1_cry_15\
        );

    \I__991\ : CascadeMux
    port map (
            O => \N__4514\,
            I => \N__4511\
        );

    \I__990\ : InMux
    port map (
            O => \N__4511\,
            I => \N__4507\
        );

    \I__989\ : InMux
    port map (
            O => \N__4510\,
            I => \N__4504\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__4507\,
            I => \N__4501\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__4504\,
            I => \reset_module_System.countZ0Z_17\
        );

    \I__986\ : Odrv4
    port map (
            O => \N__4501\,
            I => \reset_module_System.countZ0Z_17\
        );

    \I__985\ : InMux
    port map (
            O => \N__4496\,
            I => \bfn_12_4_0_\
        );

    \I__984\ : CascadeMux
    port map (
            O => \N__4493\,
            I => \N__4490\
        );

    \I__983\ : InMux
    port map (
            O => \N__4490\,
            I => \N__4487\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__4487\,
            I => \N__4483\
        );

    \I__981\ : InMux
    port map (
            O => \N__4486\,
            I => \N__4480\
        );

    \I__980\ : Span4Mux_s1_v
    port map (
            O => \N__4483\,
            I => \N__4477\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__4480\,
            I => \reset_module_System.countZ0Z_18\
        );

    \I__978\ : Odrv4
    port map (
            O => \N__4477\,
            I => \reset_module_System.countZ0Z_18\
        );

    \I__977\ : InMux
    port map (
            O => \N__4472\,
            I => \reset_module_System.count_1_cry_17\
        );

    \I__976\ : InMux
    port map (
            O => \N__4469\,
            I => \N__4465\
        );

    \I__975\ : InMux
    port map (
            O => \N__4468\,
            I => \N__4462\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__4465\,
            I => \reset_module_System.countZ0Z_2\
        );

    \I__973\ : LocalMux
    port map (
            O => \N__4462\,
            I => \reset_module_System.countZ0Z_2\
        );

    \I__972\ : InMux
    port map (
            O => \N__4457\,
            I => \N__4454\
        );

    \I__971\ : LocalMux
    port map (
            O => \N__4454\,
            I => \reset_module_System.count_1_2\
        );

    \I__970\ : InMux
    port map (
            O => \N__4451\,
            I => \reset_module_System.count_1_cry_1\
        );

    \I__969\ : InMux
    port map (
            O => \N__4448\,
            I => \N__4444\
        );

    \I__968\ : InMux
    port map (
            O => \N__4447\,
            I => \N__4441\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__4444\,
            I => \N__4438\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__4441\,
            I => \reset_module_System.countZ0Z_3\
        );

    \I__965\ : Odrv4
    port map (
            O => \N__4438\,
            I => \reset_module_System.countZ0Z_3\
        );

    \I__964\ : InMux
    port map (
            O => \N__4433\,
            I => \reset_module_System.count_1_cry_2\
        );

    \I__963\ : InMux
    port map (
            O => \N__4430\,
            I => \N__4426\
        );

    \I__962\ : InMux
    port map (
            O => \N__4429\,
            I => \N__4423\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__4426\,
            I => \reset_module_System.countZ0Z_4\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__4423\,
            I => \reset_module_System.countZ0Z_4\
        );

    \I__959\ : InMux
    port map (
            O => \N__4418\,
            I => \reset_module_System.count_1_cry_3\
        );

    \I__958\ : InMux
    port map (
            O => \N__4415\,
            I => \N__4411\
        );

    \I__957\ : InMux
    port map (
            O => \N__4414\,
            I => \N__4408\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__4411\,
            I => \reset_module_System.countZ0Z_5\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__4408\,
            I => \reset_module_System.countZ0Z_5\
        );

    \I__954\ : InMux
    port map (
            O => \N__4403\,
            I => \reset_module_System.count_1_cry_4\
        );

    \I__953\ : InMux
    port map (
            O => \N__4400\,
            I => \N__4397\
        );

    \I__952\ : LocalMux
    port map (
            O => \N__4397\,
            I => \N__4393\
        );

    \I__951\ : InMux
    port map (
            O => \N__4396\,
            I => \N__4390\
        );

    \I__950\ : Span4Mux_s1_v
    port map (
            O => \N__4393\,
            I => \N__4387\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__4390\,
            I => \reset_module_System.countZ0Z_6\
        );

    \I__948\ : Odrv4
    port map (
            O => \N__4387\,
            I => \reset_module_System.countZ0Z_6\
        );

    \I__947\ : InMux
    port map (
            O => \N__4382\,
            I => \reset_module_System.count_1_cry_5\
        );

    \I__946\ : InMux
    port map (
            O => \N__4379\,
            I => \N__4375\
        );

    \I__945\ : InMux
    port map (
            O => \N__4378\,
            I => \N__4372\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__4375\,
            I => \reset_module_System.countZ0Z_7\
        );

    \I__943\ : LocalMux
    port map (
            O => \N__4372\,
            I => \reset_module_System.countZ0Z_7\
        );

    \I__942\ : InMux
    port map (
            O => \N__4367\,
            I => \reset_module_System.count_1_cry_6\
        );

    \I__941\ : InMux
    port map (
            O => \N__4364\,
            I => \N__4360\
        );

    \I__940\ : InMux
    port map (
            O => \N__4363\,
            I => \N__4357\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__4360\,
            I => \reset_module_System.countZ0Z_8\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__4357\,
            I => \reset_module_System.countZ0Z_8\
        );

    \I__937\ : InMux
    port map (
            O => \N__4352\,
            I => \reset_module_System.count_1_cry_7\
        );

    \I__936\ : CascadeMux
    port map (
            O => \N__4349\,
            I => \N__4345\
        );

    \I__935\ : InMux
    port map (
            O => \N__4348\,
            I => \N__4342\
        );

    \I__934\ : InMux
    port map (
            O => \N__4345\,
            I => \N__4339\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__4342\,
            I => \reset_module_System.countZ0Z_9\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__4339\,
            I => \reset_module_System.countZ0Z_9\
        );

    \I__931\ : InMux
    port map (
            O => \N__4334\,
            I => \bfn_12_3_0_\
        );

    \I__930\ : InMux
    port map (
            O => \N__4331\,
            I => \N__4327\
        );

    \I__929\ : InMux
    port map (
            O => \N__4330\,
            I => \N__4324\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__4327\,
            I => \reset_module_System.countZ0Z_10\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__4324\,
            I => \reset_module_System.countZ0Z_10\
        );

    \I__926\ : InMux
    port map (
            O => \N__4319\,
            I => \reset_module_System.count_1_cry_9\
        );

    \I__925\ : CascadeMux
    port map (
            O => \N__4316\,
            I => \uart.g3_cascade_\
        );

    \I__924\ : InMux
    port map (
            O => \N__4313\,
            I => \N__4309\
        );

    \I__923\ : InMux
    port map (
            O => \N__4312\,
            I => \N__4306\
        );

    \I__922\ : LocalMux
    port map (
            O => \N__4309\,
            I => \N__4293\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__4306\,
            I => \N__4290\
        );

    \I__920\ : InMux
    port map (
            O => \N__4305\,
            I => \N__4287\
        );

    \I__919\ : InMux
    port map (
            O => \N__4304\,
            I => \N__4280\
        );

    \I__918\ : InMux
    port map (
            O => \N__4303\,
            I => \N__4280\
        );

    \I__917\ : InMux
    port map (
            O => \N__4302\,
            I => \N__4280\
        );

    \I__916\ : InMux
    port map (
            O => \N__4301\,
            I => \N__4277\
        );

    \I__915\ : InMux
    port map (
            O => \N__4300\,
            I => \N__4266\
        );

    \I__914\ : InMux
    port map (
            O => \N__4299\,
            I => \N__4266\
        );

    \I__913\ : InMux
    port map (
            O => \N__4298\,
            I => \N__4266\
        );

    \I__912\ : InMux
    port map (
            O => \N__4297\,
            I => \N__4266\
        );

    \I__911\ : InMux
    port map (
            O => \N__4296\,
            I => \N__4266\
        );

    \I__910\ : Odrv4
    port map (
            O => \N__4293\,
            I => \uart.timer_CountZ0Z_6\
        );

    \I__909\ : Odrv4
    port map (
            O => \N__4290\,
            I => \uart.timer_CountZ0Z_6\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__4287\,
            I => \uart.timer_CountZ0Z_6\
        );

    \I__907\ : LocalMux
    port map (
            O => \N__4280\,
            I => \uart.timer_CountZ0Z_6\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__4277\,
            I => \uart.timer_CountZ0Z_6\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__4266\,
            I => \uart.timer_CountZ0Z_6\
        );

    \I__904\ : InMux
    port map (
            O => \N__4253\,
            I => \N__4250\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__4250\,
            I => \uart.N_167_0\
        );

    \I__902\ : InMux
    port map (
            O => \N__4247\,
            I => \N__4243\
        );

    \I__901\ : InMux
    port map (
            O => \N__4246\,
            I => \N__4239\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__4243\,
            I => \N__4236\
        );

    \I__899\ : CascadeMux
    port map (
            O => \N__4242\,
            I => \N__4232\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__4239\,
            I => \N__4229\
        );

    \I__897\ : Span4Mux_s1_v
    port map (
            O => \N__4236\,
            I => \N__4226\
        );

    \I__896\ : InMux
    port map (
            O => \N__4235\,
            I => \N__4223\
        );

    \I__895\ : InMux
    port map (
            O => \N__4232\,
            I => \N__4220\
        );

    \I__894\ : Odrv4
    port map (
            O => \N__4229\,
            I => \reset_module_System_reset_fast\
        );

    \I__893\ : Odrv4
    port map (
            O => \N__4226\,
            I => \reset_module_System_reset_fast\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__4223\,
            I => \reset_module_System_reset_fast\
        );

    \I__891\ : LocalMux
    port map (
            O => \N__4220\,
            I => \reset_module_System_reset_fast\
        );

    \I__890\ : InMux
    port map (
            O => \N__4211\,
            I => \N__4208\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__4208\,
            I => \uart.g0_3_1\
        );

    \I__888\ : InMux
    port map (
            O => \N__4205\,
            I => \N__4199\
        );

    \I__887\ : InMux
    port map (
            O => \N__4204\,
            I => \N__4199\
        );

    \I__886\ : LocalMux
    port map (
            O => \N__4199\,
            I => \N__4189\
        );

    \I__885\ : InMux
    port map (
            O => \N__4198\,
            I => \N__4176\
        );

    \I__884\ : InMux
    port map (
            O => \N__4197\,
            I => \N__4176\
        );

    \I__883\ : InMux
    port map (
            O => \N__4196\,
            I => \N__4176\
        );

    \I__882\ : InMux
    port map (
            O => \N__4195\,
            I => \N__4176\
        );

    \I__881\ : InMux
    port map (
            O => \N__4194\,
            I => \N__4176\
        );

    \I__880\ : InMux
    port map (
            O => \N__4193\,
            I => \N__4176\
        );

    \I__879\ : InMux
    port map (
            O => \N__4192\,
            I => \N__4173\
        );

    \I__878\ : Span4Mux_h
    port map (
            O => \N__4189\,
            I => \N__4170\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__4176\,
            I => \uart.timer_CountZ0Z_3\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__4173\,
            I => \uart.timer_CountZ0Z_3\
        );

    \I__875\ : Odrv4
    port map (
            O => \N__4170\,
            I => \uart.timer_CountZ0Z_3\
        );

    \I__874\ : InMux
    port map (
            O => \N__4163\,
            I => \N__4156\
        );

    \I__873\ : InMux
    port map (
            O => \N__4162\,
            I => \N__4151\
        );

    \I__872\ : InMux
    port map (
            O => \N__4161\,
            I => \N__4151\
        );

    \I__871\ : CascadeMux
    port map (
            O => \N__4160\,
            I => \N__4148\
        );

    \I__870\ : InMux
    port map (
            O => \N__4159\,
            I => \N__4145\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__4156\,
            I => \N__4140\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__4151\,
            I => \N__4140\
        );

    \I__867\ : InMux
    port map (
            O => \N__4148\,
            I => \N__4137\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__4145\,
            I => \N__4132\
        );

    \I__865\ : Span4Mux_h
    port map (
            O => \N__4140\,
            I => \N__4132\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__4137\,
            I => \uart.timer_Count_4_repZ0Z1\
        );

    \I__863\ : Odrv4
    port map (
            O => \N__4132\,
            I => \uart.timer_Count_4_repZ0Z1\
        );

    \I__862\ : CascadeMux
    port map (
            O => \N__4127\,
            I => \N__4123\
        );

    \I__861\ : InMux
    port map (
            O => \N__4126\,
            I => \N__4120\
        );

    \I__860\ : InMux
    port map (
            O => \N__4123\,
            I => \N__4115\
        );

    \I__859\ : LocalMux
    port map (
            O => \N__4120\,
            I => \N__4109\
        );

    \I__858\ : InMux
    port map (
            O => \N__4119\,
            I => \N__4106\
        );

    \I__857\ : InMux
    port map (
            O => \N__4118\,
            I => \N__4097\
        );

    \I__856\ : LocalMux
    port map (
            O => \N__4115\,
            I => \N__4094\
        );

    \I__855\ : InMux
    port map (
            O => \N__4114\,
            I => \N__4087\
        );

    \I__854\ : InMux
    port map (
            O => \N__4113\,
            I => \N__4087\
        );

    \I__853\ : InMux
    port map (
            O => \N__4112\,
            I => \N__4087\
        );

    \I__852\ : Span4Mux_h
    port map (
            O => \N__4109\,
            I => \N__4082\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__4106\,
            I => \N__4082\
        );

    \I__850\ : InMux
    port map (
            O => \N__4105\,
            I => \N__4079\
        );

    \I__849\ : InMux
    port map (
            O => \N__4104\,
            I => \N__4068\
        );

    \I__848\ : InMux
    port map (
            O => \N__4103\,
            I => \N__4068\
        );

    \I__847\ : InMux
    port map (
            O => \N__4102\,
            I => \N__4068\
        );

    \I__846\ : InMux
    port map (
            O => \N__4101\,
            I => \N__4068\
        );

    \I__845\ : InMux
    port map (
            O => \N__4100\,
            I => \N__4068\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__4097\,
            I => \uart.timer_CountZ0Z_5\
        );

    \I__843\ : Odrv4
    port map (
            O => \N__4094\,
            I => \uart.timer_CountZ0Z_5\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__4087\,
            I => \uart.timer_CountZ0Z_5\
        );

    \I__841\ : Odrv4
    port map (
            O => \N__4082\,
            I => \uart.timer_CountZ0Z_5\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__4079\,
            I => \uart.timer_CountZ0Z_5\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__4068\,
            I => \uart.timer_CountZ0Z_5\
        );

    \I__838\ : CascadeMux
    port map (
            O => \N__4055\,
            I => \N__4052\
        );

    \I__837\ : InMux
    port map (
            O => \N__4052\,
            I => \N__4049\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__4049\,
            I => \uart.state_RNO_2Z0Z_3\
        );

    \I__835\ : InMux
    port map (
            O => \N__4046\,
            I => \N__4042\
        );

    \I__834\ : CascadeMux
    port map (
            O => \N__4045\,
            I => \N__4039\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__4042\,
            I => \N__4033\
        );

    \I__832\ : InMux
    port map (
            O => \N__4039\,
            I => \N__4021\
        );

    \I__831\ : InMux
    port map (
            O => \N__4038\,
            I => \N__4021\
        );

    \I__830\ : InMux
    port map (
            O => \N__4037\,
            I => \N__4021\
        );

    \I__829\ : InMux
    port map (
            O => \N__4036\,
            I => \N__4021\
        );

    \I__828\ : Span4Mux_h
    port map (
            O => \N__4033\,
            I => \N__4018\
        );

    \I__827\ : InMux
    port map (
            O => \N__4032\,
            I => \N__4011\
        );

    \I__826\ : InMux
    port map (
            O => \N__4031\,
            I => \N__4011\
        );

    \I__825\ : InMux
    port map (
            O => \N__4030\,
            I => \N__4011\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__4021\,
            I => \uart.un4_timer_Count_1_c2\
        );

    \I__823\ : Odrv4
    port map (
            O => \N__4018\,
            I => \uart.un4_timer_Count_1_c2\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__4011\,
            I => \uart.un4_timer_Count_1_c2\
        );

    \I__821\ : CascadeMux
    port map (
            O => \N__4004\,
            I => \N__3999\
        );

    \I__820\ : CascadeMux
    port map (
            O => \N__4003\,
            I => \N__3994\
        );

    \I__819\ : InMux
    port map (
            O => \N__4002\,
            I => \N__3991\
        );

    \I__818\ : InMux
    port map (
            O => \N__3999\,
            I => \N__3988\
        );

    \I__817\ : InMux
    port map (
            O => \N__3998\,
            I => \N__3981\
        );

    \I__816\ : InMux
    port map (
            O => \N__3997\,
            I => \N__3981\
        );

    \I__815\ : InMux
    port map (
            O => \N__3994\,
            I => \N__3981\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__3991\,
            I => \uart.timer_Count_2_repZ0Z1\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__3988\,
            I => \uart.timer_Count_2_repZ0Z1\
        );

    \I__812\ : LocalMux
    port map (
            O => \N__3981\,
            I => \uart.timer_Count_2_repZ0Z1\
        );

    \I__811\ : SRMux
    port map (
            O => \N__3974\,
            I => \N__3969\
        );

    \I__810\ : SRMux
    port map (
            O => \N__3973\,
            I => \N__3965\
        );

    \I__809\ : SRMux
    port map (
            O => \N__3972\,
            I => \N__3962\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__3969\,
            I => \N__3959\
        );

    \I__807\ : SRMux
    port map (
            O => \N__3968\,
            I => \N__3956\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__3965\,
            I => \N__3953\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__3962\,
            I => \N__3946\
        );

    \I__804\ : Span4Mux_v
    port map (
            O => \N__3959\,
            I => \N__3946\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__3956\,
            I => \N__3946\
        );

    \I__802\ : Span4Mux_v
    port map (
            O => \N__3953\,
            I => \N__3943\
        );

    \I__801\ : Span4Mux_s0_v
    port map (
            O => \N__3946\,
            I => \N__3940\
        );

    \I__800\ : Odrv4
    port map (
            O => \N__3943\,
            I => \uart.state_RNI38F97Z0Z_2\
        );

    \I__799\ : Odrv4
    port map (
            O => \N__3940\,
            I => \uart.state_RNI38F97Z0Z_2\
        );

    \I__798\ : InMux
    port map (
            O => \N__3935\,
            I => \N__3927\
        );

    \I__797\ : InMux
    port map (
            O => \N__3934\,
            I => \N__3924\
        );

    \I__796\ : CascadeMux
    port map (
            O => \N__3933\,
            I => \N__3917\
        );

    \I__795\ : CascadeMux
    port map (
            O => \N__3932\,
            I => \N__3912\
        );

    \I__794\ : CascadeMux
    port map (
            O => \N__3931\,
            I => \N__3909\
        );

    \I__793\ : InMux
    port map (
            O => \N__3930\,
            I => \N__3905\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__3927\,
            I => \N__3900\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__3924\,
            I => \N__3900\
        );

    \I__790\ : InMux
    port map (
            O => \N__3923\,
            I => \N__3893\
        );

    \I__789\ : InMux
    port map (
            O => \N__3922\,
            I => \N__3893\
        );

    \I__788\ : InMux
    port map (
            O => \N__3921\,
            I => \N__3893\
        );

    \I__787\ : InMux
    port map (
            O => \N__3920\,
            I => \N__3890\
        );

    \I__786\ : InMux
    port map (
            O => \N__3917\,
            I => \N__3885\
        );

    \I__785\ : InMux
    port map (
            O => \N__3916\,
            I => \N__3885\
        );

    \I__784\ : InMux
    port map (
            O => \N__3915\,
            I => \N__3882\
        );

    \I__783\ : InMux
    port map (
            O => \N__3912\,
            I => \N__3875\
        );

    \I__782\ : InMux
    port map (
            O => \N__3909\,
            I => \N__3875\
        );

    \I__781\ : InMux
    port map (
            O => \N__3908\,
            I => \N__3875\
        );

    \I__780\ : LocalMux
    port map (
            O => \N__3905\,
            I => \uart.timer_CountZ0Z_7\
        );

    \I__779\ : Odrv4
    port map (
            O => \N__3900\,
            I => \uart.timer_CountZ0Z_7\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__3893\,
            I => \uart.timer_CountZ0Z_7\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__3890\,
            I => \uart.timer_CountZ0Z_7\
        );

    \I__776\ : LocalMux
    port map (
            O => \N__3885\,
            I => \uart.timer_CountZ0Z_7\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__3882\,
            I => \uart.timer_CountZ0Z_7\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__3875\,
            I => \uart.timer_CountZ0Z_7\
        );

    \I__773\ : InMux
    port map (
            O => \N__3860\,
            I => \N__3857\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__3857\,
            I => \N__3854\
        );

    \I__771\ : Span4Mux_h
    port map (
            O => \N__3854\,
            I => \N__3849\
        );

    \I__770\ : InMux
    port map (
            O => \N__3853\,
            I => \N__3846\
        );

    \I__769\ : InMux
    port map (
            O => \N__3852\,
            I => \N__3843\
        );

    \I__768\ : Odrv4
    port map (
            O => \N__3849\,
            I => \uart.N_41\
        );

    \I__767\ : LocalMux
    port map (
            O => \N__3846\,
            I => \uart.N_41\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__3843\,
            I => \uart.N_41\
        );

    \I__765\ : InMux
    port map (
            O => \N__3836\,
            I => \N__3833\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__3833\,
            I => \N__3830\
        );

    \I__763\ : Span4Mux_h
    port map (
            O => \N__3830\,
            I => \N__3824\
        );

    \I__762\ : InMux
    port map (
            O => \N__3829\,
            I => \N__3821\
        );

    \I__761\ : InMux
    port map (
            O => \N__3828\,
            I => \N__3816\
        );

    \I__760\ : InMux
    port map (
            O => \N__3827\,
            I => \N__3816\
        );

    \I__759\ : Odrv4
    port map (
            O => \N__3824\,
            I => \uart.state_srsts_0_o4_0_a2_0_4\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__3821\,
            I => \uart.state_srsts_0_o4_0_a2_0_4\
        );

    \I__757\ : LocalMux
    port map (
            O => \N__3816\,
            I => \uart.state_srsts_0_o4_0_a2_0_4\
        );

    \I__756\ : CEMux
    port map (
            O => \N__3809\,
            I => \N__3806\
        );

    \I__755\ : LocalMux
    port map (
            O => \N__3806\,
            I => \N__3803\
        );

    \I__754\ : Odrv4
    port map (
            O => \N__3803\,
            I => \uart_frame_decoder.uart_data_rdy_c_0\
        );

    \I__753\ : InMux
    port map (
            O => \N__3800\,
            I => \N__3792\
        );

    \I__752\ : InMux
    port map (
            O => \N__3799\,
            I => \N__3792\
        );

    \I__751\ : InMux
    port map (
            O => \N__3798\,
            I => \N__3789\
        );

    \I__750\ : InMux
    port map (
            O => \N__3797\,
            I => \N__3786\
        );

    \I__749\ : LocalMux
    port map (
            O => \N__3792\,
            I => \N__3783\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__3789\,
            I => \uart_frame_decoder.state_1Z0Z_3\
        );

    \I__747\ : LocalMux
    port map (
            O => \N__3786\,
            I => \uart_frame_decoder.state_1Z0Z_3\
        );

    \I__746\ : Odrv12
    port map (
            O => \N__3783\,
            I => \uart_frame_decoder.state_1Z0Z_3\
        );

    \I__745\ : InMux
    port map (
            O => \N__3776\,
            I => \N__3770\
        );

    \I__744\ : InMux
    port map (
            O => \N__3775\,
            I => \N__3763\
        );

    \I__743\ : InMux
    port map (
            O => \N__3774\,
            I => \N__3763\
        );

    \I__742\ : InMux
    port map (
            O => \N__3773\,
            I => \N__3763\
        );

    \I__741\ : LocalMux
    port map (
            O => \N__3770\,
            I => \N__3759\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__3763\,
            I => \N__3756\
        );

    \I__739\ : InMux
    port map (
            O => \N__3762\,
            I => \N__3753\
        );

    \I__738\ : Span4Mux_s1_v
    port map (
            O => \N__3759\,
            I => \N__3748\
        );

    \I__737\ : Span4Mux_s1_v
    port map (
            O => \N__3756\,
            I => \N__3748\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__3753\,
            I => \uart_frame_decoder.state_1Z0Z_6\
        );

    \I__735\ : Odrv4
    port map (
            O => \N__3748\,
            I => \uart_frame_decoder.state_1Z0Z_6\
        );

    \I__734\ : InMux
    port map (
            O => \N__3743\,
            I => \N__3739\
        );

    \I__733\ : InMux
    port map (
            O => \N__3742\,
            I => \N__3736\
        );

    \I__732\ : LocalMux
    port map (
            O => \N__3739\,
            I => \N__3729\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__3736\,
            I => \N__3729\
        );

    \I__730\ : InMux
    port map (
            O => \N__3735\,
            I => \N__3724\
        );

    \I__729\ : InMux
    port map (
            O => \N__3734\,
            I => \N__3724\
        );

    \I__728\ : Odrv12
    port map (
            O => \N__3729\,
            I => \uart_frame_decoder.state_1Z0Z_2\
        );

    \I__727\ : LocalMux
    port map (
            O => \N__3724\,
            I => \uart_frame_decoder.state_1Z0Z_2\
        );

    \I__726\ : IoInMux
    port map (
            O => \N__3719\,
            I => \N__3716\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__3716\,
            I => \N__3713\
        );

    \I__724\ : IoSpan4Mux
    port map (
            O => \N__3713\,
            I => \N__3710\
        );

    \I__723\ : Odrv4
    port map (
            O => \N__3710\,
            I => \uart_frame_decoder_N_130_i\
        );

    \I__722\ : CascadeMux
    port map (
            O => \N__3707\,
            I => \reset_module_System.reset6_14_cascade_\
        );

    \I__721\ : InMux
    port map (
            O => \N__3704\,
            I => \N__3691\
        );

    \I__720\ : InMux
    port map (
            O => \N__3703\,
            I => \N__3691\
        );

    \I__719\ : InMux
    port map (
            O => \N__3702\,
            I => \N__3691\
        );

    \I__718\ : InMux
    port map (
            O => \N__3701\,
            I => \N__3691\
        );

    \I__717\ : InMux
    port map (
            O => \N__3700\,
            I => \N__3688\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__3691\,
            I => \reset_module_System.reset6_19\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__3688\,
            I => \reset_module_System.reset6_19\
        );

    \I__714\ : CascadeMux
    port map (
            O => \N__3683\,
            I => \N__3679\
        );

    \I__713\ : CascadeMux
    port map (
            O => \N__3682\,
            I => \N__3675\
        );

    \I__712\ : InMux
    port map (
            O => \N__3679\,
            I => \N__3668\
        );

    \I__711\ : InMux
    port map (
            O => \N__3678\,
            I => \N__3668\
        );

    \I__710\ : InMux
    port map (
            O => \N__3675\,
            I => \N__3668\
        );

    \I__709\ : LocalMux
    port map (
            O => \N__3668\,
            I => \N__3663\
        );

    \I__708\ : InMux
    port map (
            O => \N__3667\,
            I => \N__3658\
        );

    \I__707\ : InMux
    port map (
            O => \N__3666\,
            I => \N__3658\
        );

    \I__706\ : Odrv4
    port map (
            O => \N__3663\,
            I => \reset_module_System.reset6_14\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__3658\,
            I => \reset_module_System.reset6_14\
        );

    \I__704\ : InMux
    port map (
            O => \N__3653\,
            I => \N__3650\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__3650\,
            I => \reset_module_System.reset6_19_1\
        );

    \I__702\ : InMux
    port map (
            O => \N__3647\,
            I => \N__3644\
        );

    \I__701\ : LocalMux
    port map (
            O => \N__3644\,
            I => \reset_module_System.reset6_13\
        );

    \I__700\ : InMux
    port map (
            O => \N__3641\,
            I => \N__3635\
        );

    \I__699\ : InMux
    port map (
            O => \N__3640\,
            I => \N__3632\
        );

    \I__698\ : InMux
    port map (
            O => \N__3639\,
            I => \N__3629\
        );

    \I__697\ : InMux
    port map (
            O => \N__3638\,
            I => \N__3626\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__3635\,
            I => \N__3621\
        );

    \I__695\ : LocalMux
    port map (
            O => \N__3632\,
            I => \N__3616\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__3629\,
            I => \N__3616\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__3626\,
            I => \N__3612\
        );

    \I__692\ : CascadeMux
    port map (
            O => \N__3625\,
            I => \N__3608\
        );

    \I__691\ : CascadeMux
    port map (
            O => \N__3624\,
            I => \N__3603\
        );

    \I__690\ : Span4Mux_h
    port map (
            O => \N__3621\,
            I => \N__3595\
        );

    \I__689\ : Span4Mux_h
    port map (
            O => \N__3616\,
            I => \N__3595\
        );

    \I__688\ : InMux
    port map (
            O => \N__3615\,
            I => \N__3592\
        );

    \I__687\ : Span4Mux_h
    port map (
            O => \N__3612\,
            I => \N__3589\
        );

    \I__686\ : InMux
    port map (
            O => \N__3611\,
            I => \N__3578\
        );

    \I__685\ : InMux
    port map (
            O => \N__3608\,
            I => \N__3578\
        );

    \I__684\ : InMux
    port map (
            O => \N__3607\,
            I => \N__3578\
        );

    \I__683\ : InMux
    port map (
            O => \N__3606\,
            I => \N__3578\
        );

    \I__682\ : InMux
    port map (
            O => \N__3603\,
            I => \N__3578\
        );

    \I__681\ : InMux
    port map (
            O => \N__3602\,
            I => \N__3571\
        );

    \I__680\ : InMux
    port map (
            O => \N__3601\,
            I => \N__3571\
        );

    \I__679\ : InMux
    port map (
            O => \N__3600\,
            I => \N__3571\
        );

    \I__678\ : Odrv4
    port map (
            O => \N__3595\,
            I => \uart.stateZ0Z_3\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__3592\,
            I => \uart.stateZ0Z_3\
        );

    \I__676\ : Odrv4
    port map (
            O => \N__3589\,
            I => \uart.stateZ0Z_3\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__3578\,
            I => \uart.stateZ0Z_3\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__3571\,
            I => \uart.stateZ0Z_3\
        );

    \I__673\ : CascadeMux
    port map (
            O => \N__3560\,
            I => \N__3557\
        );

    \I__672\ : InMux
    port map (
            O => \N__3557\,
            I => \N__3554\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__3554\,
            I => \uart.g3_0_0\
        );

    \I__670\ : InMux
    port map (
            O => \N__3551\,
            I => \N__3546\
        );

    \I__669\ : InMux
    port map (
            O => \N__3550\,
            I => \N__3543\
        );

    \I__668\ : CascadeMux
    port map (
            O => \N__3549\,
            I => \N__3540\
        );

    \I__667\ : LocalMux
    port map (
            O => \N__3546\,
            I => \N__3536\
        );

    \I__666\ : LocalMux
    port map (
            O => \N__3543\,
            I => \N__3533\
        );

    \I__665\ : InMux
    port map (
            O => \N__3540\,
            I => \N__3527\
        );

    \I__664\ : InMux
    port map (
            O => \N__3539\,
            I => \N__3524\
        );

    \I__663\ : Span4Mux_v
    port map (
            O => \N__3536\,
            I => \N__3519\
        );

    \I__662\ : Span4Mux_v
    port map (
            O => \N__3533\,
            I => \N__3519\
        );

    \I__661\ : InMux
    port map (
            O => \N__3532\,
            I => \N__3512\
        );

    \I__660\ : InMux
    port map (
            O => \N__3531\,
            I => \N__3512\
        );

    \I__659\ : InMux
    port map (
            O => \N__3530\,
            I => \N__3512\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__3527\,
            I => \N__3509\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__3524\,
            I => \N__3506\
        );

    \I__656\ : Odrv4
    port map (
            O => \N__3519\,
            I => \uart.timer_CountZ0Z_4\
        );

    \I__655\ : LocalMux
    port map (
            O => \N__3512\,
            I => \uart.timer_CountZ0Z_4\
        );

    \I__654\ : Odrv4
    port map (
            O => \N__3509\,
            I => \uart.timer_CountZ0Z_4\
        );

    \I__653\ : Odrv4
    port map (
            O => \N__3506\,
            I => \uart.timer_CountZ0Z_4\
        );

    \I__652\ : InMux
    port map (
            O => \N__3497\,
            I => \N__3494\
        );

    \I__651\ : LocalMux
    port map (
            O => \N__3494\,
            I => \N__3491\
        );

    \I__650\ : Span4Mux_h
    port map (
            O => \N__3491\,
            I => \N__3488\
        );

    \I__649\ : Odrv4
    port map (
            O => \N__3488\,
            I => \uart.state_0_sqmuxa_1_d_0\
        );

    \I__648\ : CascadeMux
    port map (
            O => \N__3485\,
            I => \N__3482\
        );

    \I__647\ : InMux
    port map (
            O => \N__3482\,
            I => \N__3479\
        );

    \I__646\ : LocalMux
    port map (
            O => \N__3479\,
            I => \N__3474\
        );

    \I__645\ : InMux
    port map (
            O => \N__3478\,
            I => \N__3467\
        );

    \I__644\ : InMux
    port map (
            O => \N__3477\,
            I => \N__3467\
        );

    \I__643\ : Span4Mux_h
    port map (
            O => \N__3474\,
            I => \N__3464\
        );

    \I__642\ : InMux
    port map (
            O => \N__3473\,
            I => \N__3459\
        );

    \I__641\ : InMux
    port map (
            O => \N__3472\,
            I => \N__3459\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__3467\,
            I => \uart.timer_CountZ0Z_1\
        );

    \I__639\ : Odrv4
    port map (
            O => \N__3464\,
            I => \uart.timer_CountZ0Z_1\
        );

    \I__638\ : LocalMux
    port map (
            O => \N__3459\,
            I => \uart.timer_CountZ0Z_1\
        );

    \I__637\ : InMux
    port map (
            O => \N__3452\,
            I => \N__3449\
        );

    \I__636\ : LocalMux
    port map (
            O => \N__3449\,
            I => \uart.g1_3\
        );

    \I__635\ : InMux
    port map (
            O => \N__3446\,
            I => \N__3443\
        );

    \I__634\ : LocalMux
    port map (
            O => \N__3443\,
            I => \N__3438\
        );

    \I__633\ : InMux
    port map (
            O => \N__3442\,
            I => \N__3433\
        );

    \I__632\ : InMux
    port map (
            O => \N__3441\,
            I => \N__3433\
        );

    \I__631\ : Odrv4
    port map (
            O => \N__3438\,
            I => \uart.stateZ0Z_2\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__3433\,
            I => \uart.stateZ0Z_2\
        );

    \I__629\ : InMux
    port map (
            O => \N__3428\,
            I => \N__3424\
        );

    \I__628\ : InMux
    port map (
            O => \N__3427\,
            I => \N__3421\
        );

    \I__627\ : LocalMux
    port map (
            O => \N__3424\,
            I => \N__3418\
        );

    \I__626\ : LocalMux
    port map (
            O => \N__3421\,
            I => \N__3415\
        );

    \I__625\ : Span4Mux_s3_v
    port map (
            O => \N__3418\,
            I => \N__3410\
        );

    \I__624\ : Span4Mux_v
    port map (
            O => \N__3415\,
            I => \N__3410\
        );

    \I__623\ : Odrv4
    port map (
            O => \N__3410\,
            I => \uart.un1_state_5\
        );

    \I__622\ : InMux
    port map (
            O => \N__3407\,
            I => \N__3404\
        );

    \I__621\ : LocalMux
    port map (
            O => \N__3404\,
            I => \N__3401\
        );

    \I__620\ : Span4Mux_v
    port map (
            O => \N__3401\,
            I => \N__3397\
        );

    \I__619\ : InMux
    port map (
            O => \N__3400\,
            I => \N__3394\
        );

    \I__618\ : Span4Mux_h
    port map (
            O => \N__3397\,
            I => \N__3391\
        );

    \I__617\ : LocalMux
    port map (
            O => \N__3394\,
            I => \uart.N_177\
        );

    \I__616\ : Odrv4
    port map (
            O => \N__3391\,
            I => \uart.N_177\
        );

    \I__615\ : CascadeMux
    port map (
            O => \N__3386\,
            I => \N__3382\
        );

    \I__614\ : InMux
    port map (
            O => \N__3385\,
            I => \N__3376\
        );

    \I__613\ : InMux
    port map (
            O => \N__3382\,
            I => \N__3373\
        );

    \I__612\ : InMux
    port map (
            O => \N__3381\,
            I => \N__3368\
        );

    \I__611\ : InMux
    port map (
            O => \N__3380\,
            I => \N__3368\
        );

    \I__610\ : InMux
    port map (
            O => \N__3379\,
            I => \N__3365\
        );

    \I__609\ : LocalMux
    port map (
            O => \N__3376\,
            I => \N__3357\
        );

    \I__608\ : LocalMux
    port map (
            O => \N__3373\,
            I => \N__3357\
        );

    \I__607\ : LocalMux
    port map (
            O => \N__3368\,
            I => \N__3352\
        );

    \I__606\ : LocalMux
    port map (
            O => \N__3365\,
            I => \N__3352\
        );

    \I__605\ : InMux
    port map (
            O => \N__3364\,
            I => \N__3345\
        );

    \I__604\ : InMux
    port map (
            O => \N__3363\,
            I => \N__3345\
        );

    \I__603\ : InMux
    port map (
            O => \N__3362\,
            I => \N__3340\
        );

    \I__602\ : Span4Mux_v
    port map (
            O => \N__3357\,
            I => \N__3335\
        );

    \I__601\ : Span4Mux_s1_v
    port map (
            O => \N__3352\,
            I => \N__3335\
        );

    \I__600\ : InMux
    port map (
            O => \N__3351\,
            I => \N__3330\
        );

    \I__599\ : InMux
    port map (
            O => \N__3350\,
            I => \N__3330\
        );

    \I__598\ : LocalMux
    port map (
            O => \N__3345\,
            I => \N__3327\
        );

    \I__597\ : InMux
    port map (
            O => \N__3344\,
            I => \N__3322\
        );

    \I__596\ : InMux
    port map (
            O => \N__3343\,
            I => \N__3322\
        );

    \I__595\ : LocalMux
    port map (
            O => \N__3340\,
            I => reset_system
        );

    \I__594\ : Odrv4
    port map (
            O => \N__3335\,
            I => reset_system
        );

    \I__593\ : LocalMux
    port map (
            O => \N__3330\,
            I => reset_system
        );

    \I__592\ : Odrv12
    port map (
            O => \N__3327\,
            I => reset_system
        );

    \I__591\ : LocalMux
    port map (
            O => \N__3322\,
            I => reset_system
        );

    \I__590\ : InMux
    port map (
            O => \N__3311\,
            I => \N__3308\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__3308\,
            I => \uart.N_28_mux\
        );

    \I__588\ : CascadeMux
    port map (
            O => \N__3305\,
            I => \uart.N_8_cascade_\
        );

    \I__587\ : InMux
    port map (
            O => \N__3302\,
            I => \N__3297\
        );

    \I__586\ : InMux
    port map (
            O => \N__3301\,
            I => \N__3294\
        );

    \I__585\ : InMux
    port map (
            O => \N__3300\,
            I => \N__3291\
        );

    \I__584\ : LocalMux
    port map (
            O => \N__3297\,
            I => \N__3286\
        );

    \I__583\ : LocalMux
    port map (
            O => \N__3294\,
            I => \N__3286\
        );

    \I__582\ : LocalMux
    port map (
            O => \N__3291\,
            I => \N__3281\
        );

    \I__581\ : Span4Mux_h
    port map (
            O => \N__3286\,
            I => \N__3281\
        );

    \I__580\ : Odrv4
    port map (
            O => \N__3281\,
            I => \uart_frame_decoder.state_1Z0Z_4\
        );

    \I__579\ : CascadeMux
    port map (
            O => \N__3278\,
            I => \N__3272\
        );

    \I__578\ : InMux
    port map (
            O => \N__3277\,
            I => \N__3269\
        );

    \I__577\ : InMux
    port map (
            O => \N__3276\,
            I => \N__3266\
        );

    \I__576\ : InMux
    port map (
            O => \N__3275\,
            I => \N__3261\
        );

    \I__575\ : InMux
    port map (
            O => \N__3272\,
            I => \N__3261\
        );

    \I__574\ : LocalMux
    port map (
            O => \N__3269\,
            I => \N__3258\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__3266\,
            I => \N__3255\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__3261\,
            I => \N__3252\
        );

    \I__571\ : Odrv12
    port map (
            O => \N__3258\,
            I => \uart_frame_decoder.state_1Z0Z_5\
        );

    \I__570\ : Odrv4
    port map (
            O => \N__3255\,
            I => \uart_frame_decoder.state_1Z0Z_5\
        );

    \I__569\ : Odrv4
    port map (
            O => \N__3252\,
            I => \uart_frame_decoder.state_1Z0Z_5\
        );

    \I__568\ : InMux
    port map (
            O => \N__3245\,
            I => \N__3242\
        );

    \I__567\ : LocalMux
    port map (
            O => \N__3242\,
            I => \reset_module_System.reset6_3\
        );

    \I__566\ : InMux
    port map (
            O => \N__3239\,
            I => \N__3236\
        );

    \I__565\ : LocalMux
    port map (
            O => \N__3236\,
            I => \uart.timer_Count_RNI3B101Z0Z_6\
        );

    \I__564\ : CascadeMux
    port map (
            O => \N__3233\,
            I => \N__3228\
        );

    \I__563\ : InMux
    port map (
            O => \N__3232\,
            I => \N__3221\
        );

    \I__562\ : InMux
    port map (
            O => \N__3231\,
            I => \N__3221\
        );

    \I__561\ : InMux
    port map (
            O => \N__3228\,
            I => \N__3221\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__3221\,
            I => \N__3218\
        );

    \I__559\ : Odrv4
    port map (
            O => \N__3218\,
            I => \uart.un4_timer_Count_1_c5\
        );

    \I__558\ : InMux
    port map (
            O => \N__3215\,
            I => \N__3212\
        );

    \I__557\ : LocalMux
    port map (
            O => \N__3212\,
            I => \N__3209\
        );

    \I__556\ : Odrv4
    port map (
            O => \N__3209\,
            I => \uart.un1_state_2_0_a3_2\
        );

    \I__555\ : CascadeMux
    port map (
            O => \N__3206\,
            I => \N__3203\
        );

    \I__554\ : InMux
    port map (
            O => \N__3203\,
            I => \N__3196\
        );

    \I__553\ : InMux
    port map (
            O => \N__3202\,
            I => \N__3196\
        );

    \I__552\ : CascadeMux
    port map (
            O => \N__3201\,
            I => \N__3192\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__3196\,
            I => \N__3189\
        );

    \I__550\ : InMux
    port map (
            O => \N__3195\,
            I => \N__3184\
        );

    \I__549\ : InMux
    port map (
            O => \N__3192\,
            I => \N__3184\
        );

    \I__548\ : Odrv4
    port map (
            O => \N__3189\,
            I => \uart.timer_CountZ0Z_0\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__3184\,
            I => \uart.timer_CountZ0Z_0\
        );

    \I__546\ : InMux
    port map (
            O => \N__3179\,
            I => \N__3176\
        );

    \I__545\ : LocalMux
    port map (
            O => \N__3176\,
            I => \uart.timer_Count_RNI22NA1Z0Z_4\
        );

    \I__544\ : CascadeMux
    port map (
            O => \N__3173\,
            I => \N__3168\
        );

    \I__543\ : CascadeMux
    port map (
            O => \N__3172\,
            I => \N__3165\
        );

    \I__542\ : InMux
    port map (
            O => \N__3171\,
            I => \N__3162\
        );

    \I__541\ : InMux
    port map (
            O => \N__3168\,
            I => \N__3153\
        );

    \I__540\ : InMux
    port map (
            O => \N__3165\,
            I => \N__3153\
        );

    \I__539\ : LocalMux
    port map (
            O => \N__3162\,
            I => \N__3150\
        );

    \I__538\ : CascadeMux
    port map (
            O => \N__3161\,
            I => \N__3143\
        );

    \I__537\ : CascadeMux
    port map (
            O => \N__3160\,
            I => \N__3140\
        );

    \I__536\ : CascadeMux
    port map (
            O => \N__3159\,
            I => \N__3136\
        );

    \I__535\ : InMux
    port map (
            O => \N__3158\,
            I => \N__3132\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__3153\,
            I => \N__3129\
        );

    \I__533\ : Span4Mux_h
    port map (
            O => \N__3150\,
            I => \N__3126\
        );

    \I__532\ : InMux
    port map (
            O => \N__3149\,
            I => \N__3123\
        );

    \I__531\ : InMux
    port map (
            O => \N__3148\,
            I => \N__3120\
        );

    \I__530\ : InMux
    port map (
            O => \N__3147\,
            I => \N__3115\
        );

    \I__529\ : InMux
    port map (
            O => \N__3146\,
            I => \N__3115\
        );

    \I__528\ : InMux
    port map (
            O => \N__3143\,
            I => \N__3106\
        );

    \I__527\ : InMux
    port map (
            O => \N__3140\,
            I => \N__3106\
        );

    \I__526\ : InMux
    port map (
            O => \N__3139\,
            I => \N__3106\
        );

    \I__525\ : InMux
    port map (
            O => \N__3136\,
            I => \N__3106\
        );

    \I__524\ : InMux
    port map (
            O => \N__3135\,
            I => \N__3103\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__3132\,
            I => \N__3098\
        );

    \I__522\ : Span4Mux_h
    port map (
            O => \N__3129\,
            I => \N__3098\
        );

    \I__521\ : Odrv4
    port map (
            O => \N__3126\,
            I => \uart.bit_CountZ0Z_0\
        );

    \I__520\ : LocalMux
    port map (
            O => \N__3123\,
            I => \uart.bit_CountZ0Z_0\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__3120\,
            I => \uart.bit_CountZ0Z_0\
        );

    \I__518\ : LocalMux
    port map (
            O => \N__3115\,
            I => \uart.bit_CountZ0Z_0\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__3106\,
            I => \uart.bit_CountZ0Z_0\
        );

    \I__516\ : LocalMux
    port map (
            O => \N__3103\,
            I => \uart.bit_CountZ0Z_0\
        );

    \I__515\ : Odrv4
    port map (
            O => \N__3098\,
            I => \uart.bit_CountZ0Z_0\
        );

    \I__514\ : CascadeMux
    port map (
            O => \N__3083\,
            I => \N__3080\
        );

    \I__513\ : InMux
    port map (
            O => \N__3080\,
            I => \N__3077\
        );

    \I__512\ : LocalMux
    port map (
            O => \N__3077\,
            I => \N__3070\
        );

    \I__511\ : InMux
    port map (
            O => \N__3076\,
            I => \N__3067\
        );

    \I__510\ : InMux
    port map (
            O => \N__3075\,
            I => \N__3062\
        );

    \I__509\ : InMux
    port map (
            O => \N__3074\,
            I => \N__3062\
        );

    \I__508\ : InMux
    port map (
            O => \N__3073\,
            I => \N__3056\
        );

    \I__507\ : Span4Mux_v
    port map (
            O => \N__3070\,
            I => \N__3053\
        );

    \I__506\ : LocalMux
    port map (
            O => \N__3067\,
            I => \N__3048\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__3062\,
            I => \N__3048\
        );

    \I__504\ : InMux
    port map (
            O => \N__3061\,
            I => \N__3045\
        );

    \I__503\ : InMux
    port map (
            O => \N__3060\,
            I => \N__3040\
        );

    \I__502\ : InMux
    port map (
            O => \N__3059\,
            I => \N__3040\
        );

    \I__501\ : LocalMux
    port map (
            O => \N__3056\,
            I => \uart.bit_CountZ0Z_2\
        );

    \I__500\ : Odrv4
    port map (
            O => \N__3053\,
            I => \uart.bit_CountZ0Z_2\
        );

    \I__499\ : Odrv4
    port map (
            O => \N__3048\,
            I => \uart.bit_CountZ0Z_2\
        );

    \I__498\ : LocalMux
    port map (
            O => \N__3045\,
            I => \uart.bit_CountZ0Z_2\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__3040\,
            I => \uart.bit_CountZ0Z_2\
        );

    \I__496\ : InMux
    port map (
            O => \N__3029\,
            I => \N__3026\
        );

    \I__495\ : LocalMux
    port map (
            O => \N__3026\,
            I => \N__3020\
        );

    \I__494\ : InMux
    port map (
            O => \N__3025\,
            I => \N__3017\
        );

    \I__493\ : InMux
    port map (
            O => \N__3024\,
            I => \N__3012\
        );

    \I__492\ : InMux
    port map (
            O => \N__3023\,
            I => \N__3012\
        );

    \I__491\ : Span4Mux_h
    port map (
            O => \N__3020\,
            I => \N__3004\
        );

    \I__490\ : LocalMux
    port map (
            O => \N__3017\,
            I => \N__2999\
        );

    \I__489\ : LocalMux
    port map (
            O => \N__3012\,
            I => \N__2999\
        );

    \I__488\ : InMux
    port map (
            O => \N__3011\,
            I => \N__2994\
        );

    \I__487\ : InMux
    port map (
            O => \N__3010\,
            I => \N__2994\
        );

    \I__486\ : InMux
    port map (
            O => \N__3009\,
            I => \N__2987\
        );

    \I__485\ : InMux
    port map (
            O => \N__3008\,
            I => \N__2987\
        );

    \I__484\ : InMux
    port map (
            O => \N__3007\,
            I => \N__2987\
        );

    \I__483\ : Odrv4
    port map (
            O => \N__3004\,
            I => \uart.bit_CountZ0Z_1\
        );

    \I__482\ : Odrv4
    port map (
            O => \N__2999\,
            I => \uart.bit_CountZ0Z_1\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__2994\,
            I => \uart.bit_CountZ0Z_1\
        );

    \I__480\ : LocalMux
    port map (
            O => \N__2987\,
            I => \uart.bit_CountZ0Z_1\
        );

    \I__479\ : CascadeMux
    port map (
            O => \N__2978\,
            I => \uart.g1_4_cascade_\
        );

    \I__478\ : InMux
    port map (
            O => \N__2975\,
            I => \N__2972\
        );

    \I__477\ : LocalMux
    port map (
            O => \N__2972\,
            I => \N__2969\
        );

    \I__476\ : Span4Mux_v
    port map (
            O => \N__2969\,
            I => \N__2966\
        );

    \I__475\ : Odrv4
    port map (
            O => \N__2966\,
            I => \uart.g1_0\
        );

    \I__474\ : CascadeMux
    port map (
            O => \N__2963\,
            I => \N__2958\
        );

    \I__473\ : InMux
    port map (
            O => \N__2962\,
            I => \N__2954\
        );

    \I__472\ : InMux
    port map (
            O => \N__2961\,
            I => \N__2947\
        );

    \I__471\ : InMux
    port map (
            O => \N__2958\,
            I => \N__2947\
        );

    \I__470\ : InMux
    port map (
            O => \N__2957\,
            I => \N__2947\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__2954\,
            I => \uart.timer_Count_fastZ0Z_2\
        );

    \I__468\ : LocalMux
    port map (
            O => \N__2947\,
            I => \uart.timer_Count_fastZ0Z_2\
        );

    \I__467\ : CascadeMux
    port map (
            O => \N__2942\,
            I => \reset_module_System.reset6_11_cascade_\
        );

    \I__466\ : CascadeMux
    port map (
            O => \N__2939\,
            I => \reset_module_System.reset6_19_cascade_\
        );

    \I__465\ : InMux
    port map (
            O => \N__2936\,
            I => \N__2933\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__2933\,
            I => \uart.N_66\
        );

    \I__463\ : InMux
    port map (
            O => \N__2930\,
            I => \N__2927\
        );

    \I__462\ : LocalMux
    port map (
            O => \N__2927\,
            I => \uart.N_51\
        );

    \I__461\ : InMux
    port map (
            O => \N__2924\,
            I => \N__2919\
        );

    \I__460\ : CascadeMux
    port map (
            O => \N__2923\,
            I => \N__2914\
        );

    \I__459\ : InMux
    port map (
            O => \N__2922\,
            I => \N__2911\
        );

    \I__458\ : LocalMux
    port map (
            O => \N__2919\,
            I => \N__2908\
        );

    \I__457\ : InMux
    port map (
            O => \N__2918\,
            I => \N__2901\
        );

    \I__456\ : InMux
    port map (
            O => \N__2917\,
            I => \N__2901\
        );

    \I__455\ : InMux
    port map (
            O => \N__2914\,
            I => \N__2901\
        );

    \I__454\ : LocalMux
    port map (
            O => \N__2911\,
            I => \uart.timer_Count_fastZ0Z_3\
        );

    \I__453\ : Odrv4
    port map (
            O => \N__2908\,
            I => \uart.timer_Count_fastZ0Z_3\
        );

    \I__452\ : LocalMux
    port map (
            O => \N__2901\,
            I => \uart.timer_Count_fastZ0Z_3\
        );

    \I__451\ : InMux
    port map (
            O => \N__2894\,
            I => \N__2891\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__2891\,
            I => \N__2888\
        );

    \I__449\ : Odrv12
    port map (
            O => \N__2888\,
            I => \uart.N_5\
        );

    \I__448\ : CascadeMux
    port map (
            O => \N__2885\,
            I => \N__2880\
        );

    \I__447\ : CascadeMux
    port map (
            O => \N__2884\,
            I => \N__2877\
        );

    \I__446\ : InMux
    port map (
            O => \N__2883\,
            I => \N__2874\
        );

    \I__445\ : InMux
    port map (
            O => \N__2880\,
            I => \N__2871\
        );

    \I__444\ : InMux
    port map (
            O => \N__2877\,
            I => \N__2868\
        );

    \I__443\ : LocalMux
    port map (
            O => \N__2874\,
            I => \N__2863\
        );

    \I__442\ : LocalMux
    port map (
            O => \N__2871\,
            I => \N__2863\
        );

    \I__441\ : LocalMux
    port map (
            O => \N__2868\,
            I => \uart.stateZ0Z_1\
        );

    \I__440\ : Odrv4
    port map (
            O => \N__2863\,
            I => \uart.stateZ0Z_1\
        );

    \I__439\ : InMux
    port map (
            O => \N__2858\,
            I => \N__2855\
        );

    \I__438\ : LocalMux
    port map (
            O => \N__2855\,
            I => \uart.N_151\
        );

    \I__437\ : CascadeMux
    port map (
            O => \N__2852\,
            I => \N__2849\
        );

    \I__436\ : InMux
    port map (
            O => \N__2849\,
            I => \N__2842\
        );

    \I__435\ : InMux
    port map (
            O => \N__2848\,
            I => \N__2842\
        );

    \I__434\ : InMux
    port map (
            O => \N__2847\,
            I => \N__2838\
        );

    \I__433\ : LocalMux
    port map (
            O => \N__2842\,
            I => \N__2831\
        );

    \I__432\ : InMux
    port map (
            O => \N__2841\,
            I => \N__2828\
        );

    \I__431\ : LocalMux
    port map (
            O => \N__2838\,
            I => \N__2825\
        );

    \I__430\ : InMux
    port map (
            O => \N__2837\,
            I => \N__2816\
        );

    \I__429\ : InMux
    port map (
            O => \N__2836\,
            I => \N__2816\
        );

    \I__428\ : InMux
    port map (
            O => \N__2835\,
            I => \N__2816\
        );

    \I__427\ : InMux
    port map (
            O => \N__2834\,
            I => \N__2816\
        );

    \I__426\ : Odrv4
    port map (
            O => \N__2831\,
            I => \uart.N_174\
        );

    \I__425\ : LocalMux
    port map (
            O => \N__2828\,
            I => \uart.N_174\
        );

    \I__424\ : Odrv4
    port map (
            O => \N__2825\,
            I => \uart.N_174\
        );

    \I__423\ : LocalMux
    port map (
            O => \N__2816\,
            I => \uart.N_174\
        );

    \I__422\ : InMux
    port map (
            O => \N__2807\,
            I => \N__2804\
        );

    \I__421\ : LocalMux
    port map (
            O => \N__2804\,
            I => \uart.state_srsts_0_a3_2_0_4\
        );

    \I__420\ : InMux
    port map (
            O => \N__2801\,
            I => \N__2798\
        );

    \I__419\ : LocalMux
    port map (
            O => \N__2798\,
            I => \N__2794\
        );

    \I__418\ : InMux
    port map (
            O => \N__2797\,
            I => \N__2791\
        );

    \I__417\ : Odrv4
    port map (
            O => \N__2794\,
            I => \uart.state_1_sqmuxa\
        );

    \I__416\ : LocalMux
    port map (
            O => \N__2791\,
            I => \uart.state_1_sqmuxa\
        );

    \I__415\ : InMux
    port map (
            O => \N__2786\,
            I => \N__2783\
        );

    \I__414\ : LocalMux
    port map (
            O => \N__2783\,
            I => \N__2780\
        );

    \I__413\ : Odrv4
    port map (
            O => \N__2780\,
            I => \uart.data_AuxZ0Z_3\
        );

    \I__412\ : CEMux
    port map (
            O => \N__2777\,
            I => \N__2774\
        );

    \I__411\ : LocalMux
    port map (
            O => \N__2774\,
            I => \N__2771\
        );

    \I__410\ : Odrv12
    port map (
            O => \N__2771\,
            I => \uart.N_117_0\
        );

    \I__409\ : InMux
    port map (
            O => \N__2768\,
            I => \N__2765\
        );

    \I__408\ : LocalMux
    port map (
            O => \N__2765\,
            I => \N__2762\
        );

    \I__407\ : Span4Mux_h
    port map (
            O => \N__2762\,
            I => \N__2759\
        );

    \I__406\ : Odrv4
    port map (
            O => \N__2759\,
            I => \uart.data_AuxZ0Z_4\
        );

    \I__405\ : CEMux
    port map (
            O => \N__2756\,
            I => \N__2753\
        );

    \I__404\ : LocalMux
    port map (
            O => \N__2753\,
            I => \N__2750\
        );

    \I__403\ : Span4Mux_h
    port map (
            O => \N__2750\,
            I => \N__2747\
        );

    \I__402\ : Odrv4
    port map (
            O => \N__2747\,
            I => \uart.N_116_0\
        );

    \I__401\ : SRMux
    port map (
            O => \N__2744\,
            I => \N__2736\
        );

    \I__400\ : SRMux
    port map (
            O => \N__2743\,
            I => \N__2733\
        );

    \I__399\ : SRMux
    port map (
            O => \N__2742\,
            I => \N__2730\
        );

    \I__398\ : SRMux
    port map (
            O => \N__2741\,
            I => \N__2723\
        );

    \I__397\ : SRMux
    port map (
            O => \N__2740\,
            I => \N__2720\
        );

    \I__396\ : SRMux
    port map (
            O => \N__2739\,
            I => \N__2717\
        );

    \I__395\ : LocalMux
    port map (
            O => \N__2736\,
            I => \N__2713\
        );

    \I__394\ : LocalMux
    port map (
            O => \N__2733\,
            I => \N__2708\
        );

    \I__393\ : LocalMux
    port map (
            O => \N__2730\,
            I => \N__2708\
        );

    \I__392\ : SRMux
    port map (
            O => \N__2729\,
            I => \N__2705\
        );

    \I__391\ : InMux
    port map (
            O => \N__2728\,
            I => \N__2697\
        );

    \I__390\ : InMux
    port map (
            O => \N__2727\,
            I => \N__2697\
        );

    \I__389\ : InMux
    port map (
            O => \N__2726\,
            I => \N__2697\
        );

    \I__388\ : LocalMux
    port map (
            O => \N__2723\,
            I => \N__2689\
        );

    \I__387\ : LocalMux
    port map (
            O => \N__2720\,
            I => \N__2689\
        );

    \I__386\ : LocalMux
    port map (
            O => \N__2717\,
            I => \N__2686\
        );

    \I__385\ : InMux
    port map (
            O => \N__2716\,
            I => \N__2683\
        );

    \I__384\ : Span4Mux_h
    port map (
            O => \N__2713\,
            I => \N__2679\
        );

    \I__383\ : Span4Mux_v
    port map (
            O => \N__2708\,
            I => \N__2676\
        );

    \I__382\ : LocalMux
    port map (
            O => \N__2705\,
            I => \N__2673\
        );

    \I__381\ : SRMux
    port map (
            O => \N__2704\,
            I => \N__2670\
        );

    \I__380\ : LocalMux
    port map (
            O => \N__2697\,
            I => \N__2667\
        );

    \I__379\ : InMux
    port map (
            O => \N__2696\,
            I => \N__2660\
        );

    \I__378\ : InMux
    port map (
            O => \N__2695\,
            I => \N__2660\
        );

    \I__377\ : InMux
    port map (
            O => \N__2694\,
            I => \N__2660\
        );

    \I__376\ : Span4Mux_v
    port map (
            O => \N__2689\,
            I => \N__2653\
        );

    \I__375\ : Span4Mux_s2_v
    port map (
            O => \N__2686\,
            I => \N__2653\
        );

    \I__374\ : LocalMux
    port map (
            O => \N__2683\,
            I => \N__2653\
        );

    \I__373\ : InMux
    port map (
            O => \N__2682\,
            I => \N__2650\
        );

    \I__372\ : Odrv4
    port map (
            O => \N__2679\,
            I => \uart.state_RNIAFHLZ0Z_4\
        );

    \I__371\ : Odrv4
    port map (
            O => \N__2676\,
            I => \uart.state_RNIAFHLZ0Z_4\
        );

    \I__370\ : Odrv12
    port map (
            O => \N__2673\,
            I => \uart.state_RNIAFHLZ0Z_4\
        );

    \I__369\ : LocalMux
    port map (
            O => \N__2670\,
            I => \uart.state_RNIAFHLZ0Z_4\
        );

    \I__368\ : Odrv4
    port map (
            O => \N__2667\,
            I => \uart.state_RNIAFHLZ0Z_4\
        );

    \I__367\ : LocalMux
    port map (
            O => \N__2660\,
            I => \uart.state_RNIAFHLZ0Z_4\
        );

    \I__366\ : Odrv4
    port map (
            O => \N__2653\,
            I => \uart.state_RNIAFHLZ0Z_4\
        );

    \I__365\ : LocalMux
    port map (
            O => \N__2650\,
            I => \uart.state_RNIAFHLZ0Z_4\
        );

    \I__364\ : CascadeMux
    port map (
            O => \N__2633\,
            I => \N__2629\
        );

    \I__363\ : CascadeMux
    port map (
            O => \N__2632\,
            I => \N__2623\
        );

    \I__362\ : InMux
    port map (
            O => \N__2629\,
            I => \N__2615\
        );

    \I__361\ : InMux
    port map (
            O => \N__2628\,
            I => \N__2615\
        );

    \I__360\ : InMux
    port map (
            O => \N__2627\,
            I => \N__2602\
        );

    \I__359\ : InMux
    port map (
            O => \N__2626\,
            I => \N__2602\
        );

    \I__358\ : InMux
    port map (
            O => \N__2623\,
            I => \N__2602\
        );

    \I__357\ : InMux
    port map (
            O => \N__2622\,
            I => \N__2602\
        );

    \I__356\ : InMux
    port map (
            O => \N__2621\,
            I => \N__2602\
        );

    \I__355\ : InMux
    port map (
            O => \N__2620\,
            I => \N__2602\
        );

    \I__354\ : LocalMux
    port map (
            O => \N__2615\,
            I => \uart.timer_CountZ0Z_2\
        );

    \I__353\ : LocalMux
    port map (
            O => \N__2602\,
            I => \uart.timer_CountZ0Z_2\
        );

    \I__352\ : CascadeMux
    port map (
            O => \N__2597\,
            I => \uart.state_srsts_0_a3_1_4_cascade_\
        );

    \I__351\ : InMux
    port map (
            O => \N__2594\,
            I => \N__2590\
        );

    \I__350\ : InMux
    port map (
            O => \N__2593\,
            I => \N__2587\
        );

    \I__349\ : LocalMux
    port map (
            O => \N__2590\,
            I => \uart.timer_Count_fastZ0Z_4\
        );

    \I__348\ : LocalMux
    port map (
            O => \N__2587\,
            I => \uart.timer_Count_fastZ0Z_4\
        );

    \I__347\ : CascadeMux
    port map (
            O => \N__2582\,
            I => \N__2579\
        );

    \I__346\ : InMux
    port map (
            O => \N__2579\,
            I => \N__2576\
        );

    \I__345\ : LocalMux
    port map (
            O => \N__2576\,
            I => \N__2573\
        );

    \I__344\ : Span4Mux_v
    port map (
            O => \N__2573\,
            I => \N__2570\
        );

    \I__343\ : Odrv4
    port map (
            O => \N__2570\,
            I => \uart.timer_Count10lto4_0\
        );

    \I__342\ : CascadeMux
    port map (
            O => \N__2567\,
            I => \uart.timer_Count10lto4_0_cascade_\
        );

    \I__341\ : CascadeMux
    port map (
            O => \N__2564\,
            I => \uart.N_51_cascade_\
        );

    \I__340\ : CascadeMux
    port map (
            O => \N__2561\,
            I => \N__2558\
        );

    \I__339\ : InMux
    port map (
            O => \N__2558\,
            I => \N__2554\
        );

    \I__338\ : InMux
    port map (
            O => \N__2557\,
            I => \N__2551\
        );

    \I__337\ : LocalMux
    port map (
            O => \N__2554\,
            I => \uart.N_146_0\
        );

    \I__336\ : LocalMux
    port map (
            O => \N__2551\,
            I => \uart.N_146_0\
        );

    \I__335\ : CascadeMux
    port map (
            O => \N__2546\,
            I => \uart.data_14_1_cascade_\
        );

    \I__334\ : SRMux
    port map (
            O => \N__2543\,
            I => \N__2540\
        );

    \I__333\ : LocalMux
    port map (
            O => \N__2540\,
            I => \N__2537\
        );

    \I__332\ : Span4Mux_s2_v
    port map (
            O => \N__2537\,
            I => \N__2534\
        );

    \I__331\ : Odrv4
    port map (
            O => \N__2534\,
            I => \uart.state_RNILS533Z0Z_4\
        );

    \I__330\ : CascadeMux
    port map (
            O => \N__2531\,
            I => \uart.state_RNILS533Z0Z_4_cascade_\
        );

    \I__329\ : CEMux
    port map (
            O => \N__2528\,
            I => \N__2525\
        );

    \I__328\ : LocalMux
    port map (
            O => \N__2525\,
            I => \uart.state_1_sqmuxa_0\
        );

    \I__327\ : CascadeMux
    port map (
            O => \N__2522\,
            I => \uart.un4_timer_Count_1_c2_cascade_\
        );

    \I__326\ : InMux
    port map (
            O => \N__2519\,
            I => \N__2513\
        );

    \I__325\ : InMux
    port map (
            O => \N__2518\,
            I => \N__2513\
        );

    \I__324\ : LocalMux
    port map (
            O => \N__2513\,
            I => \uart.data_Auxce_0_4\
        );

    \I__323\ : CEMux
    port map (
            O => \N__2510\,
            I => \N__2507\
        );

    \I__322\ : LocalMux
    port map (
            O => \N__2507\,
            I => \N__2504\
        );

    \I__321\ : Odrv4
    port map (
            O => \N__2504\,
            I => \uart.N_113_0\
        );

    \I__320\ : InMux
    port map (
            O => \N__2501\,
            I => \N__2498\
        );

    \I__319\ : LocalMux
    port map (
            O => \N__2498\,
            I => \N__2494\
        );

    \I__318\ : InMux
    port map (
            O => \N__2497\,
            I => \N__2491\
        );

    \I__317\ : Odrv4
    port map (
            O => \N__2494\,
            I => \uart.N_133_0\
        );

    \I__316\ : LocalMux
    port map (
            O => \N__2491\,
            I => \uart.N_133_0\
        );

    \I__315\ : InMux
    port map (
            O => \N__2486\,
            I => \N__2480\
        );

    \I__314\ : InMux
    port map (
            O => \N__2485\,
            I => \N__2480\
        );

    \I__313\ : LocalMux
    port map (
            O => \N__2480\,
            I => \uart.stateZ0Z_0\
        );

    \I__312\ : InMux
    port map (
            O => \N__2477\,
            I => \N__2469\
        );

    \I__311\ : InMux
    port map (
            O => \N__2476\,
            I => \N__2469\
        );

    \I__310\ : CascadeMux
    port map (
            O => \N__2475\,
            I => \N__2466\
        );

    \I__309\ : InMux
    port map (
            O => \N__2474\,
            I => \N__2460\
        );

    \I__308\ : LocalMux
    port map (
            O => \N__2469\,
            I => \N__2457\
        );

    \I__307\ : InMux
    port map (
            O => \N__2466\,
            I => \N__2448\
        );

    \I__306\ : InMux
    port map (
            O => \N__2465\,
            I => \N__2448\
        );

    \I__305\ : InMux
    port map (
            O => \N__2464\,
            I => \N__2448\
        );

    \I__304\ : InMux
    port map (
            O => \N__2463\,
            I => \N__2448\
        );

    \I__303\ : LocalMux
    port map (
            O => \N__2460\,
            I => \uart.N_175\
        );

    \I__302\ : Odrv4
    port map (
            O => \N__2457\,
            I => \uart.N_175\
        );

    \I__301\ : LocalMux
    port map (
            O => \N__2448\,
            I => \uart.N_175\
        );

    \I__300\ : CascadeMux
    port map (
            O => \N__2441\,
            I => \uart.data_Auxce_0_6_cascade_\
        );

    \I__299\ : CEMux
    port map (
            O => \N__2438\,
            I => \N__2435\
        );

    \I__298\ : LocalMux
    port map (
            O => \N__2435\,
            I => \N__2432\
        );

    \I__297\ : Odrv4
    port map (
            O => \N__2432\,
            I => \uart.N_114_0\
        );

    \I__296\ : InMux
    port map (
            O => \N__2429\,
            I => \N__2426\
        );

    \I__295\ : LocalMux
    port map (
            O => \N__2426\,
            I => \uart.data_Aux_esr_RNO_0Z0Z_5\
        );

    \I__294\ : InMux
    port map (
            O => \N__2423\,
            I => \N__2420\
        );

    \I__293\ : LocalMux
    port map (
            O => \N__2420\,
            I => \N__2417\
        );

    \I__292\ : Odrv12
    port map (
            O => \N__2417\,
            I => \uart.data_AuxZ0Z_5\
        );

    \I__291\ : CEMux
    port map (
            O => \N__2414\,
            I => \N__2411\
        );

    \I__290\ : LocalMux
    port map (
            O => \N__2411\,
            I => \N__2408\
        );

    \I__289\ : Odrv4
    port map (
            O => \N__2408\,
            I => \uart.N_115_0\
        );

    \I__288\ : CascadeMux
    port map (
            O => \N__2405\,
            I => \uart.data_Aux_esr_RNO_0Z0Z_0_cascade_\
        );

    \I__287\ : CEMux
    port map (
            O => \N__2402\,
            I => \N__2399\
        );

    \I__286\ : LocalMux
    port map (
            O => \N__2399\,
            I => \N__2396\
        );

    \I__285\ : Odrv4
    port map (
            O => \N__2396\,
            I => \uart.N_120_0\
        );

    \I__284\ : InMux
    port map (
            O => \N__2393\,
            I => \N__2389\
        );

    \I__283\ : InMux
    port map (
            O => \N__2392\,
            I => \N__2386\
        );

    \I__282\ : LocalMux
    port map (
            O => \N__2389\,
            I => \uart.data_Auxce_0_0\
        );

    \I__281\ : LocalMux
    port map (
            O => \N__2386\,
            I => \uart.data_Auxce_0_0\
        );

    \I__280\ : CascadeMux
    port map (
            O => \N__2381\,
            I => \uart.data_Aux_esr_RNO_0Z0Z_1_cascade_\
        );

    \I__279\ : InMux
    port map (
            O => \N__2378\,
            I => \N__2375\
        );

    \I__278\ : LocalMux
    port map (
            O => \N__2375\,
            I => \N__2372\
        );

    \I__277\ : Odrv4
    port map (
            O => \N__2372\,
            I => \uart.data_AuxZ0Z_1\
        );

    \I__276\ : CEMux
    port map (
            O => \N__2369\,
            I => \N__2366\
        );

    \I__275\ : LocalMux
    port map (
            O => \N__2366\,
            I => \N__2363\
        );

    \I__274\ : Odrv4
    port map (
            O => \N__2363\,
            I => \uart.N_119_0\
        );

    \I__273\ : InMux
    port map (
            O => \N__2360\,
            I => \N__2357\
        );

    \I__272\ : LocalMux
    port map (
            O => \N__2357\,
            I => \uart.data_Auxce_0_2\
        );

    \I__271\ : CascadeMux
    port map (
            O => \N__2354\,
            I => \uart.data_Aux_esr_RNO_0Z0Z_3_cascade_\
        );

    \I__270\ : CascadeMux
    port map (
            O => \N__2351\,
            I => \uart.data_Aux_esr_RNO_0Z0Z_4_cascade_\
        );

    \I__269\ : InMux
    port map (
            O => \N__2348\,
            I => \N__2345\
        );

    \I__268\ : LocalMux
    port map (
            O => \N__2345\,
            I => uart_data_4
        );

    \I__267\ : InMux
    port map (
            O => \N__2342\,
            I => \N__2338\
        );

    \I__266\ : InMux
    port map (
            O => \N__2341\,
            I => \N__2335\
        );

    \I__265\ : LocalMux
    port map (
            O => \N__2338\,
            I => uart_data_5
        );

    \I__264\ : LocalMux
    port map (
            O => \N__2335\,
            I => uart_data_5
        );

    \I__263\ : InMux
    port map (
            O => \N__2330\,
            I => \N__2327\
        );

    \I__262\ : LocalMux
    port map (
            O => \N__2327\,
            I => \N__2324\
        );

    \I__261\ : Span4Mux_s2_v
    port map (
            O => \N__2324\,
            I => \N__2321\
        );

    \I__260\ : Odrv4
    port map (
            O => \N__2321\,
            I => \uart.data_AuxZ0Z_6\
        );

    \I__259\ : InMux
    port map (
            O => \N__2318\,
            I => \N__2315\
        );

    \I__258\ : LocalMux
    port map (
            O => \N__2315\,
            I => uart_data_6
        );

    \I__257\ : InMux
    port map (
            O => \N__2312\,
            I => \N__2309\
        );

    \I__256\ : LocalMux
    port map (
            O => \N__2309\,
            I => \N__2306\
        );

    \I__255\ : Odrv4
    port map (
            O => \N__2306\,
            I => \uart.data_AuxZ0Z_7\
        );

    \I__254\ : CascadeMux
    port map (
            O => \N__2303\,
            I => \N__2299\
        );

    \I__253\ : InMux
    port map (
            O => \N__2302\,
            I => \N__2296\
        );

    \I__252\ : InMux
    port map (
            O => \N__2299\,
            I => \N__2293\
        );

    \I__251\ : LocalMux
    port map (
            O => \N__2296\,
            I => uart_data_7
        );

    \I__250\ : LocalMux
    port map (
            O => \N__2293\,
            I => uart_data_7
        );

    \I__249\ : CascadeMux
    port map (
            O => \N__2288\,
            I => \uart.N_147_0_0_cascade_\
        );

    \I__248\ : CascadeMux
    port map (
            O => \N__2285\,
            I => \uart.g3_1_0_cascade_\
        );

    \I__247\ : InMux
    port map (
            O => \N__2282\,
            I => \N__2279\
        );

    \I__246\ : LocalMux
    port map (
            O => \N__2279\,
            I => \N__2276\
        );

    \I__245\ : Span4Mux_s2_v
    port map (
            O => \N__2276\,
            I => \N__2273\
        );

    \I__244\ : Odrv4
    port map (
            O => \N__2273\,
            I => \uart.g0_4_0\
        );

    \I__243\ : CascadeMux
    port map (
            O => \N__2270\,
            I => \uart.N_175_cascade_\
        );

    \I__242\ : CascadeMux
    port map (
            O => \N__2267\,
            I => \N__2262\
        );

    \I__241\ : InMux
    port map (
            O => \N__2266\,
            I => \N__2255\
        );

    \I__240\ : InMux
    port map (
            O => \N__2265\,
            I => \N__2255\
        );

    \I__239\ : InMux
    port map (
            O => \N__2262\,
            I => \N__2248\
        );

    \I__238\ : InMux
    port map (
            O => \N__2261\,
            I => \N__2248\
        );

    \I__237\ : InMux
    port map (
            O => \N__2260\,
            I => \N__2248\
        );

    \I__236\ : LocalMux
    port map (
            O => \N__2255\,
            I => \uart_frame_decoder.state_1Z0Z_1\
        );

    \I__235\ : LocalMux
    port map (
            O => \N__2248\,
            I => \uart_frame_decoder.state_1Z0Z_1\
        );

    \I__234\ : IoInMux
    port map (
            O => \N__2243\,
            I => \N__2240\
        );

    \I__233\ : LocalMux
    port map (
            O => \N__2240\,
            I => \uart_frame_decoder_N_129_i\
        );

    \I__232\ : CascadeMux
    port map (
            O => \N__2237\,
            I => \uart_frame_decoder.state_1_srsts_i_i_a2_3_0Z0Z_0_cascade_\
        );

    \I__231\ : InMux
    port map (
            O => \N__2234\,
            I => \N__2228\
        );

    \I__230\ : InMux
    port map (
            O => \N__2233\,
            I => \N__2228\
        );

    \I__229\ : LocalMux
    port map (
            O => \N__2228\,
            I => \uart_frame_decoder.N_67\
        );

    \I__228\ : InMux
    port map (
            O => \N__2225\,
            I => \N__2222\
        );

    \I__227\ : LocalMux
    port map (
            O => \N__2222\,
            I => \uart_frame_decoder.N_61\
        );

    \I__226\ : CascadeMux
    port map (
            O => \N__2219\,
            I => \uart_frame_decoder.N_67_cascade_\
        );

    \I__225\ : InMux
    port map (
            O => \N__2216\,
            I => \N__2212\
        );

    \I__224\ : InMux
    port map (
            O => \N__2215\,
            I => \N__2209\
        );

    \I__223\ : LocalMux
    port map (
            O => \N__2212\,
            I => \uart_frame_decoder.state_1_srsts_0_i_a2_0_0_2\
        );

    \I__222\ : LocalMux
    port map (
            O => \N__2209\,
            I => \uart_frame_decoder.state_1_srsts_0_i_a2_0_0_2\
        );

    \I__221\ : InMux
    port map (
            O => \N__2204\,
            I => \N__2201\
        );

    \I__220\ : LocalMux
    port map (
            O => \N__2201\,
            I => \N__2198\
        );

    \I__219\ : Odrv4
    port map (
            O => \N__2198\,
            I => \uart.data_AuxZ0Z_0\
        );

    \I__218\ : InMux
    port map (
            O => \N__2195\,
            I => \N__2191\
        );

    \I__217\ : InMux
    port map (
            O => \N__2194\,
            I => \N__2188\
        );

    \I__216\ : LocalMux
    port map (
            O => \N__2191\,
            I => uart_data_0
        );

    \I__215\ : LocalMux
    port map (
            O => \N__2188\,
            I => uart_data_0
        );

    \I__214\ : InMux
    port map (
            O => \N__2183\,
            I => \N__2180\
        );

    \I__213\ : LocalMux
    port map (
            O => \N__2180\,
            I => \N__2177\
        );

    \I__212\ : Odrv4
    port map (
            O => \N__2177\,
            I => uart_data_1
        );

    \I__211\ : InMux
    port map (
            O => \N__2174\,
            I => \N__2171\
        );

    \I__210\ : LocalMux
    port map (
            O => \N__2171\,
            I => \uart.data_AuxZ0Z_2\
        );

    \I__209\ : InMux
    port map (
            O => \N__2168\,
            I => \N__2164\
        );

    \I__208\ : InMux
    port map (
            O => \N__2167\,
            I => \N__2161\
        );

    \I__207\ : LocalMux
    port map (
            O => \N__2164\,
            I => uart_data_2
        );

    \I__206\ : LocalMux
    port map (
            O => \N__2161\,
            I => uart_data_2
        );

    \I__205\ : InMux
    port map (
            O => \N__2156\,
            I => \N__2153\
        );

    \I__204\ : LocalMux
    port map (
            O => \N__2153\,
            I => \N__2150\
        );

    \I__203\ : Odrv4
    port map (
            O => \N__2150\,
            I => uart_data_3
        );

    \I__202\ : CascadeMux
    port map (
            O => \N__2147\,
            I => \uart.data_Aux_esr_RNO_0Z0Z_2_cascade_\
        );

    \I__201\ : CEMux
    port map (
            O => \N__2144\,
            I => \N__2141\
        );

    \I__200\ : LocalMux
    port map (
            O => \N__2141\,
            I => \N__2138\
        );

    \I__199\ : Odrv4
    port map (
            O => \N__2138\,
            I => \uart.N_118_0\
        );

    \I__198\ : CascadeMux
    port map (
            O => \N__2135\,
            I => \uart_frame_decoder.state_1_srsts_0_i_a2_0_0_1Z0Z_2_cascade_\
        );

    \I__197\ : InMux
    port map (
            O => \N__2132\,
            I => \N__2129\
        );

    \I__196\ : LocalMux
    port map (
            O => \N__2129\,
            I => \uart_frame_decoder.N_49\
        );

    \I__195\ : CascadeMux
    port map (
            O => \N__2126\,
            I => \uart_frame_decoder.N_58_4_cascade_\
        );

    \I__194\ : InMux
    port map (
            O => \N__2123\,
            I => \N__2120\
        );

    \I__193\ : LocalMux
    port map (
            O => \N__2120\,
            I => \N__2117\
        );

    \I__192\ : Odrv4
    port map (
            O => \N__2117\,
            I => \uart_frame_decoder.N_32_i_1\
        );

    \I__191\ : CascadeMux
    port map (
            O => \N__2114\,
            I => \uart.state_0_sqmuxa_1_d_cascade_\
        );

    \I__190\ : CascadeMux
    port map (
            O => \N__2111\,
            I => \uart.m13_0_0_o2_2_cascade_\
        );

    \I__189\ : CascadeMux
    port map (
            O => \N__2108\,
            I => \uart.N_10_cascade_\
        );

    \I__188\ : CascadeMux
    port map (
            O => \N__2105\,
            I => \uart.data_Auxce_0_2_cascade_\
        );

    \I__187\ : CascadeMux
    port map (
            O => \N__2102\,
            I => \uart_frame_decoder.N_43_cascade_\
        );

    \I__186\ : CascadeMux
    port map (
            O => \N__2099\,
            I => \uart_frame_decoder.state_1_srsts_i_i_0_0_cascade_\
        );

    \I__185\ : IoInMux
    port map (
            O => \N__2096\,
            I => \N__2093\
        );

    \I__184\ : LocalMux
    port map (
            O => \N__2093\,
            I => \N__2090\
        );

    \I__183\ : Span4Mux_s0_v
    port map (
            O => \N__2090\,
            I => \N__2087\
        );

    \I__182\ : Odrv4
    port map (
            O => \N__2087\,
            I => \uart_frame_decoder_N_131_i\
        );

    \I__181\ : CascadeMux
    port map (
            O => \N__2084\,
            I => \N__2081\
        );

    \I__180\ : InMux
    port map (
            O => \N__2081\,
            I => \N__2078\
        );

    \I__179\ : LocalMux
    port map (
            O => \N__2078\,
            I => \uart_frame_decoder.state_1Z0Z_0\
        );

    \I__178\ : InMux
    port map (
            O => \N__2075\,
            I => \N__2072\
        );

    \I__177\ : LocalMux
    port map (
            O => \N__2072\,
            I => \uart_frame_decoder.state_1_srsts_0_i_1_1\
        );

    \I__176\ : InMux
    port map (
            O => \N__2069\,
            I => \N__2066\
        );

    \I__175\ : LocalMux
    port map (
            O => \N__2066\,
            I => \uart_frame_decoder.N_58_4\
        );

    \IN_MUX_bfv_12_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_2_0_\
        );

    \IN_MUX_bfv_12_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \reset_module_System.count_1_cry_8\,
            carryinitout => \bfn_12_3_0_\
        );

    \IN_MUX_bfv_12_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \reset_module_System.count_1_cry_16\,
            carryinitout => \bfn_12_4_0_\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNO_2_0_LC_7_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__3773\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2260\,
            lcout => OPEN,
            ltout => \uart_frame_decoder.N_43_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNO_1_0_LC_7_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100010000"
        )
    port map (
            in0 => \N__3381\,
            in1 => \N__4914\,
            in2 => \N__2102\,
            in3 => \N__2132\,
            lcout => OPEN,
            ltout => \uart_frame_decoder.state_1_srsts_i_i_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_0_LC_7_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100000111"
        )
    port map (
            in0 => \N__2215\,
            in1 => \N__2233\,
            in2 => \N__2099\,
            in3 => \N__2123\,
            lcout => \uart_frame_decoder.state_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4814\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_1_LC_7_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010001000"
        )
    port map (
            in0 => \N__2234\,
            in1 => \N__4915\,
            in2 => \N__2267\,
            in3 => \N__2075\,
            lcout => \uart_frame_decoder.state_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4814\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_esr_RNI7FFE_4_LC_7_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__3775\,
            in1 => \N__3302\,
            in2 => \_gnd_net_\,
            in3 => \N__3277\,
            lcout => \uart_frame_decoder_N_131_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNO_0_1_LC_7_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110111011101"
        )
    port map (
            in0 => \N__3380\,
            in1 => \N__4913\,
            in2 => \N__2084\,
            in3 => \N__2069\,
            lcout => \uart_frame_decoder.state_1_srsts_0_i_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_srsts_0_i_a2_0_4_1_LC_7_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2341\,
            in1 => \N__2167\,
            in2 => \N__2303\,
            in3 => \N__2194\,
            lcout => \uart_frame_decoder.N_58_4\,
            ltout => \uart_frame_decoder.N_58_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNO_0_0_LC_7_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__2261\,
            in1 => \N__4912\,
            in2 => \N__2126\,
            in3 => \N__3774\,
            lcout => \uart_frame_decoder.N_32_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_esr_2_LC_7_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5134\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uart.data_AuxZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4812\,
            ce => \N__2144\,
            sr => \N__2739\
        );

    \uart.bit_Count_RNO_0_0_LC_7_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111010101"
        )
    port map (
            in0 => \N__3639\,
            in1 => \N__3551\,
            in2 => \N__2582\,
            in3 => \N__4126\,
            lcout => OPEN,
            ltout => \uart.state_0_sqmuxa_1_d_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.bit_Count_0_LC_7_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110001001100"
        )
    port map (
            in0 => \N__3428\,
            in1 => \N__3147\,
            in2 => \N__2114\,
            in3 => \N__2501\,
            lcout => \uart.bit_CountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4809\,
            ce => 'H',
            sr => \N__4724\
        );

    \uart.bit_Count_RNO_2_2_LC_7_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__3011\,
            in1 => \N__3135\,
            in2 => \_gnd_net_\,
            in3 => \N__4313\,
            lcout => OPEN,
            ltout => \uart.m13_0_0_o2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.bit_Count_RNO_0_2_LC_7_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__2894\,
            in1 => \N__3935\,
            in2 => \N__2111\,
            in3 => \N__5061\,
            lcout => OPEN,
            ltout => \uart.N_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.bit_Count_2_LC_7_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110000000001110"
        )
    port map (
            in0 => \N__5062\,
            in1 => \N__3641\,
            in2 => \N__2108\,
            in3 => \N__3073\,
            lcout => \uart.bit_CountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4809\,
            ce => 'H',
            sr => \N__4724\
        );

    \uart.bit_Count_RNILKM9_0_2_LC_7_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3061\,
            in2 => \_gnd_net_\,
            in3 => \N__3010\,
            lcout => \uart.data_Auxce_0_2\,
            ltout => \uart.data_Auxce_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_esr_RNO_0_2_LC_7_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001000000"
        )
    port map (
            in0 => \N__3146\,
            in1 => \N__2847\,
            in2 => \N__2105\,
            in3 => \N__2474\,
            lcout => OPEN,
            ltout => \uart.data_Aux_esr_RNO_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_esr_RNO_2_LC_7_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__2716\,
            in1 => \_gnd_net_\,
            in2 => \N__2147\,
            in3 => \_gnd_net_\,
            lcout => \uart.N_118_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_esr_0_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5157\,
            lcout => \uart.data_AuxZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4806\,
            ce => \N__2402\,
            sr => \N__2740\
        );

    \uart.bit_Count_RNIETHE_2_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__3158\,
            in1 => \N__3076\,
            in2 => \_gnd_net_\,
            in3 => \N__3025\,
            lcout => \uart.N_177\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_esr_7_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5161\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uart.data_AuxZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4803\,
            ce => \N__2510\,
            sr => \N__2744\
        );

    \uart.bit_Count_RNO_0_1_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3427\,
            in2 => \_gnd_net_\,
            in3 => \N__2497\,
            lcout => \uart.g0_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_esr_6_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5162\,
            lcout => \uart.data_AuxZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4798\,
            ce => \N__2438\,
            sr => \N__2741\
        );

    \uart_frame_decoder.state_1_srsts_0_i_a2_0_0_1_2_LC_8_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2342\,
            in2 => \_gnd_net_\,
            in3 => \N__2168\,
            lcout => OPEN,
            ltout => \uart_frame_decoder.state_1_srsts_0_i_a2_0_0_1Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNI5BVV_1_LC_8_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__2265\,
            in1 => \N__2195\,
            in2 => \N__2135\,
            in3 => \N__2302\,
            lcout => \uart_frame_decoder.state_1_srsts_0_i_a2_0_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNO_0_2_LC_8_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__3735\,
            in1 => \N__4910\,
            in2 => \_gnd_net_\,
            in3 => \N__3379\,
            lcout => \uart_frame_decoder.N_61\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNO_3_0_LC_8_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3301\,
            in1 => \N__3799\,
            in2 => \N__3278\,
            in3 => \N__3734\,
            lcout => \uart_frame_decoder.N_49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_esr_RNI19FE_3_LC_8_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__3800\,
            in1 => \N__3275\,
            in2 => \_gnd_net_\,
            in3 => \N__2266\,
            lcout => \uart_frame_decoder_N_129_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_srsts_i_i_a2_3_0_0_LC_8_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2348\,
            in2 => \_gnd_net_\,
            in3 => \N__4247\,
            lcout => OPEN,
            ltout => \uart_frame_decoder.state_1_srsts_i_i_a2_3_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_srsts_i_i_a2_3_0_LC_8_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2156\,
            in1 => \N__2318\,
            in2 => \N__2237\,
            in3 => \N__2183\,
            lcout => \uart_frame_decoder.N_67\,
            ltout => \uart_frame_decoder.N_67_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_2_LC_8_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__4911\,
            in1 => \N__2225\,
            in2 => \N__2219\,
            in3 => \N__2216\,
            lcout => \uart_frame_decoder.state_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4813\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_esr_0_LC_8_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2204\,
            lcout => uart_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4810\,
            ce => \N__2528\,
            sr => \N__2543\
        );

    \uart.data_esr_1_LC_8_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2378\,
            lcout => uart_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4810\,
            ce => \N__2528\,
            sr => \N__2543\
        );

    \uart.data_esr_2_LC_8_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2174\,
            lcout => uart_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4810\,
            ce => \N__2528\,
            sr => \N__2543\
        );

    \uart.data_esr_3_LC_8_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__2786\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => uart_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4810\,
            ce => \N__2528\,
            sr => \N__2543\
        );

    \uart.data_esr_4_LC_8_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2768\,
            lcout => uart_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4810\,
            ce => \N__2528\,
            sr => \N__2543\
        );

    \uart.data_esr_5_LC_8_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2423\,
            lcout => uart_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4810\,
            ce => \N__2528\,
            sr => \N__2543\
        );

    \uart.data_esr_6_LC_8_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2330\,
            lcout => uart_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4810\,
            ce => \N__2528\,
            sr => \N__2543\
        );

    \uart.data_esr_7_LC_8_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__2312\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => uart_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4810\,
            ce => \N__2528\,
            sr => \N__2543\
        );

    \uart.bit_Count_RNO_3_1_LC_8_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3934\,
            in2 => \_gnd_net_\,
            in3 => \N__4312\,
            lcout => OPEN,
            ltout => \uart.N_147_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.bit_Count_RNO_1_1_LC_8_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100010"
        )
    port map (
            in0 => \N__3149\,
            in1 => \N__3640\,
            in2 => \N__2288\,
            in3 => \N__5063\,
            lcout => OPEN,
            ltout => \uart.g3_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.bit_Count_1_LC_8_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001001101010"
        )
    port map (
            in0 => \N__3009\,
            in1 => \N__3497\,
            in2 => \N__2285\,
            in3 => \N__2282\,
            lcout => \uart.bit_CountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4807\,
            ce => 'H',
            sr => \N__4723\
        );

    \uart.bit_Count_RNILKM9_2_LC_8_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3059\,
            in2 => \_gnd_net_\,
            in3 => \N__3007\,
            lcout => \uart.data_Auxce_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_RNI3UCP2_4_LC_8_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__4119\,
            in1 => \N__2557\,
            in2 => \N__3549\,
            in3 => \N__3215\,
            lcout => \uart.N_175\,
            ltout => \uart.N_175_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_esr_RNO_0_0_LC_8_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000000000"
        )
    port map (
            in0 => \N__2841\,
            in1 => \N__3148\,
            in2 => \N__2270\,
            in3 => \N__2392\,
            lcout => OPEN,
            ltout => \uart.data_Aux_esr_RNO_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_esr_RNO_0_LC_8_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2405\,
            in3 => \N__2682\,
            lcout => \uart.N_120_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.bit_Count_RNILKM9_1_2_LC_8_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3060\,
            in2 => \_gnd_net_\,
            in3 => \N__3008\,
            lcout => \uart.data_Auxce_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_esr_RNO_0_1_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__2837\,
            in1 => \N__3139\,
            in2 => \N__2475\,
            in3 => \N__2393\,
            lcout => OPEN,
            ltout => \uart.data_Aux_esr_RNO_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_esr_RNO_1_LC_8_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__2694\,
            in1 => \_gnd_net_\,
            in2 => \N__2381\,
            in3 => \_gnd_net_\,
            lcout => \uart.N_119_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_esr_1_LC_8_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5156\,
            lcout => \uart.data_AuxZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4804\,
            ce => \N__2369\,
            sr => \N__2742\
        );

    \uart.data_Aux_esr_RNO_0_3_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__2360\,
            in1 => \N__2836\,
            in2 => \N__3160\,
            in3 => \N__2465\,
            lcout => OPEN,
            ltout => \uart.data_Aux_esr_RNO_0Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_esr_RNO_3_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2354\,
            in3 => \N__2695\,
            lcout => \uart.N_117_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_esr_RNO_0_4_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001000"
        )
    port map (
            in0 => \N__2519\,
            in1 => \N__2835\,
            in2 => \N__3161\,
            in3 => \N__2464\,
            lcout => OPEN,
            ltout => \uart.data_Aux_esr_RNO_0Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_esr_RNO_4_LC_8_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2351\,
            in3 => \N__2696\,
            lcout => \uart.N_116_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_esr_RNO_0_5_LC_8_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__2518\,
            in1 => \N__2834\,
            in2 => \N__3159\,
            in3 => \N__2463\,
            lcout => \uart.data_Aux_esr_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_0_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111110010"
        )
    port map (
            in0 => \N__2485\,
            in1 => \N__5158\,
            in2 => \N__3386\,
            in3 => \N__2801\,
            lcout => \uart.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4799\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_esr_RNO_7_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111010101010"
        )
    port map (
            in0 => \N__2728\,
            in1 => \N__2476\,
            in2 => \N__2852\,
            in3 => \N__3400\,
            lcout => \uart.N_113_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.bit_Count_RNI4ENK_2_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3074\,
            in1 => \N__3023\,
            in2 => \N__3172\,
            in3 => \N__3638\,
            lcout => \uart.N_133_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_1_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001000"
        )
    port map (
            in0 => \N__2486\,
            in1 => \N__5159\,
            in2 => \N__2884\,
            in3 => \N__3385\,
            lcout => \uart.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4799\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_esr_RNO_0_6_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__3075\,
            in1 => \_gnd_net_\,
            in2 => \N__3173\,
            in3 => \N__3024\,
            lcout => OPEN,
            ltout => \uart.data_Auxce_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_esr_RNO_6_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011101100"
        )
    port map (
            in0 => \N__2477\,
            in1 => \N__2727\,
            in2 => \N__2441\,
            in3 => \N__2848\,
            lcout => \uart.N_114_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_esr_RNO_5_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__2726\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2429\,
            lcout => \uart.N_115_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_esr_5_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5160\,
            lcout => \uart.data_AuxZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4794\,
            ce => \N__2414\,
            sr => \N__2743\
        );

    \uart.state_RNO_1_4_LC_9_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__4193\,
            in1 => \N__3530\,
            in2 => \N__4127\,
            in3 => \N__2620\,
            lcout => \uart.g1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_RNIN6BL_0_LC_9_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3202\,
            in2 => \_gnd_net_\,
            in3 => \N__3477\,
            lcout => \uart.un4_timer_Count_1_c2\,
            ltout => \uart.un4_timer_Count_1_c2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_RNIH8CL1_4_LC_9_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4194\,
            in1 => \N__2621\,
            in2 => \N__2522\,
            in3 => \N__3531\,
            lcout => \uart.un4_timer_Count_1_c5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_4_LC_9_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__3532\,
            in1 => \N__4037\,
            in2 => \N__2632\,
            in3 => \N__4196\,
            lcout => \uart.timer_CountZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4811\,
            ce => 'H',
            sr => \N__3972\
        );

    \uart.timer_Count_1_LC_9_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__3478\,
            in1 => \_gnd_net_\,
            in2 => \N__3206\,
            in3 => \_gnd_net_\,
            lcout => \uart.timer_CountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4811\,
            ce => 'H',
            sr => \N__3972\
        );

    \uart.timer_Count_3_LC_9_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__2622\,
            in1 => \N__4036\,
            in2 => \_gnd_net_\,
            in3 => \N__4195\,
            lcout => \uart.timer_CountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4811\,
            ce => 'H',
            sr => \N__3972\
        );

    \uart.timer_Count_fast_4_LC_9_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__4198\,
            in1 => \N__2627\,
            in2 => \N__4045\,
            in3 => \N__2594\,
            lcout => \uart.timer_Count_fastZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4811\,
            ce => 'H',
            sr => \N__3972\
        );

    \uart.timer_Count_4_rep1_LC_9_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__2626\,
            in1 => \N__4197\,
            in2 => \N__4160\,
            in3 => \N__4038\,
            lcout => \uart.timer_Count_4_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4811\,
            ce => 'H',
            sr => \N__3972\
        );

    \uart.timer_Count_RNI1HBL_6_LC_9_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4301\,
            in2 => \_gnd_net_\,
            in3 => \N__4105\,
            lcout => \uart.state_srsts_0_o4_0_a2_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNI3TGU_4_LC_9_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001010"
        )
    port map (
            in0 => \N__5051\,
            in1 => \_gnd_net_\,
            in2 => \N__4242\,
            in3 => \N__3915\,
            lcout => OPEN,
            ltout => \uart.state_srsts_0_a3_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNICGLN3_2_LC_9_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101000001010"
        )
    port map (
            in0 => \N__2807\,
            in1 => \N__3852\,
            in2 => \N__2597\,
            in3 => \N__3829\,
            lcout => \uart.N_66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_fast_RNIHHG81_2_LC_9_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2957\,
            in2 => \N__2923\,
            in3 => \N__3472\,
            lcout => \uart.N_146_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_fast_RNIT1EN1_4_LC_9_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__3473\,
            in1 => \N__2593\,
            in2 => \N__2963\,
            in3 => \N__2917\,
            lcout => \uart.N_41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_fast_RNILTQT_2_LC_9_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__2918\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2961\,
            lcout => \uart.timer_Count10lto4_0\,
            ltout => \uart.timer_Count10lto4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_RNIQAJ83_4_LC_9_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__3239\,
            in1 => \_gnd_net_\,
            in2 => \N__2567\,
            in3 => \N__3179\,
            lcout => \uart.N_51\,
            ltout => \uart.N_51_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_2_LC_9_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000101"
        )
    port map (
            in0 => \N__2858\,
            in1 => \N__2883\,
            in2 => \N__2564\,
            in3 => \N__3362\,
            lcout => \uart.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4808\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_4_rep1_RNIHBMA2_LC_9_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100110011"
        )
    port map (
            in0 => \N__4159\,
            in1 => \N__3916\,
            in2 => \N__2561\,
            in3 => \N__3827\,
            lcout => OPEN,
            ltout => \uart.data_14_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNILS533_4_LC_9_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101110101010"
        )
    port map (
            in0 => \N__3344\,
            in1 => \N__5104\,
            in2 => \N__2546\,
            in3 => \N__5037\,
            lcout => \uart.state_RNILS533Z0Z_4\,
            ltout => \uart.state_RNILS533Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNICRQ06_4_LC_9_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__2797\,
            in1 => \_gnd_net_\,
            in2 => \N__2531\,
            in3 => \_gnd_net_\,
            lcout => \uart.state_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNO_0_2_LC_9_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010100000101"
        )
    port map (
            in0 => \N__3442\,
            in1 => \_gnd_net_\,
            in2 => \N__2885\,
            in3 => \N__5105\,
            lcout => \uart.N_151\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNIAFHL_4_LC_9_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011101"
        )
    port map (
            in0 => \N__5035\,
            in1 => \N__3343\,
            in2 => \_gnd_net_\,
            in3 => \N__3602\,
            lcout => \uart.state_RNIAFHLZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNID2BC_4_LC_9_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__3601\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5034\,
            lcout => \uart.N_174\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNIB0BC_2_LC_9_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3600\,
            in2 => \_gnd_net_\,
            in3 => \N__3441\,
            lcout => \uart.state_srsts_0_a3_2_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNINUKT2_4_LC_9_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000000000"
        )
    port map (
            in0 => \N__3828\,
            in1 => \N__3853\,
            in2 => \N__3933\,
            in3 => \N__5036\,
            lcout => \uart.state_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_esr_3_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5106\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uart.data_AuxZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4800\,
            ce => \N__2777\,
            sr => \N__2704\
        );

    \uart.data_Aux_esr_4_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5107\,
            lcout => \uart.data_AuxZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4795\,
            ce => \N__2756\,
            sr => \N__2729\
        );

    \uart.timer_Count_fast_3_LC_10_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__4032\,
            in1 => \_gnd_net_\,
            in2 => \N__2633\,
            in3 => \N__2922\,
            lcout => \uart.timer_Count_fastZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4805\,
            ce => 'H',
            sr => \N__3968\
        );

    \uart.timer_Count_2_LC_10_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2628\,
            in2 => \_gnd_net_\,
            in3 => \N__4030\,
            lcout => \uart.timer_CountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4805\,
            ce => 'H',
            sr => \N__3968\
        );

    \uart.timer_Count_fast_2_LC_10_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__4031\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2962\,
            lcout => \uart.timer_Count_fastZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4805\,
            ce => 'H',
            sr => \N__3968\
        );

    \uart_frame_decoder.state_1_6_LC_10_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__3351\,
            in1 => \N__3276\,
            in2 => \N__4917\,
            in3 => \N__3762\,
            lcout => \uart_frame_decoder.state_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4801\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNI9O1P_2_LC_10_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__4400\,
            in1 => \N__4448\,
            in2 => \N__5189\,
            in3 => \N__4468\,
            lcout => OPEN,
            ltout => \reset_module_System.reset6_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNIN3HK3_2_LC_10_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3653\,
            in1 => \N__3647\,
            in2 => \N__2942\,
            in3 => \N__3245\,
            lcout => \reset_module_System.reset6_19\,
            ltout => \reset_module_System.reset6_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.reset_fast_LC_10_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111111111111"
        )
    port map (
            in0 => \N__4609\,
            in1 => \_gnd_net_\,
            in2 => \N__2939\,
            in3 => \N__3667\,
            lcout => \reset_module_System_reset_fast\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4801\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.reset_LC_10_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__4608\,
            in1 => \N__3666\,
            in2 => \_gnd_net_\,
            in3 => \N__3700\,
            lcout => reset_system,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4801\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNI38F97_2_LC_10_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__3350\,
            in1 => \N__2936\,
            in2 => \_gnd_net_\,
            in3 => \N__2930\,
            lcout => \uart.state_RNI38F97Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.bit_Count_RNO_4_1_LC_10_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4002\,
            in2 => \_gnd_net_\,
            in3 => \N__4192\,
            lcout => \uart.g3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.bit_Count_RNO_1_2_LC_10_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__4163\,
            in1 => \N__4102\,
            in2 => \N__4004\,
            in3 => \N__2924\,
            lcout => \uart.N_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_5_LC_10_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__4103\,
            in1 => \_gnd_net_\,
            in2 => \N__3233\,
            in3 => \_gnd_net_\,
            lcout => \uart.timer_CountZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4796\,
            ce => 'H',
            sr => \N__3974\
        );

    \uart.timer_Count_RNI3B101_6_LC_10_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__4297\,
            in1 => \N__3908\,
            in2 => \_gnd_net_\,
            in3 => \N__4100\,
            lcout => \uart.timer_Count_RNI3B101Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_7_LC_10_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__3232\,
            in1 => \N__4118\,
            in2 => \N__3932\,
            in3 => \N__4300\,
            lcout => \uart.timer_CountZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4796\,
            ce => 'H',
            sr => \N__3974\
        );

    \uart.timer_Count_6_LC_10_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__4299\,
            in1 => \N__3231\,
            in2 => \_gnd_net_\,
            in3 => \N__4104\,
            lcout => \uart.timer_CountZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4796\,
            ce => 'H',
            sr => \N__3974\
        );

    \uart.timer_Count_RNIJTGR_0_LC_10_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4296\,
            in2 => \N__3201\,
            in3 => \N__5033\,
            lcout => \uart.un1_state_2_0_a3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_0_LC_10_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3195\,
            lcout => \uart.timer_CountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4796\,
            ce => 'H',
            sr => \N__3974\
        );

    \uart.timer_Count_RNI22NA1_4_LC_10_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__4101\,
            in1 => \N__3539\,
            in2 => \N__3931\,
            in3 => \N__4298\,
            lcout => \uart.timer_Count_RNI22NA1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNO_3_4_LC_10_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3607\,
            in1 => \N__3171\,
            in2 => \N__3083\,
            in3 => \N__3029\,
            lcout => OPEN,
            ltout => \uart.g1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_4_LC_10_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__4253\,
            in1 => \N__3452\,
            in2 => \N__2978\,
            in3 => \N__2975\,
            lcout => \uart.stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4791\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNO_2_4_LC_10_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__3922\,
            in1 => \N__3363\,
            in2 => \_gnd_net_\,
            in3 => \N__4304\,
            lcout => \uart.g1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNO_1_3_LC_10_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001110110011"
        )
    port map (
            in0 => \N__4303\,
            in1 => \N__3606\,
            in2 => \N__4055\,
            in3 => \N__3446\,
            lcout => \uart.N_28_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNIGLM11_4_LC_10_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001111"
        )
    port map (
            in0 => \N__3921\,
            in1 => \N__4302\,
            in2 => \N__3624\,
            in3 => \N__5041\,
            lcout => \uart.un1_state_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNO_0_3_LC_10_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110101"
        )
    port map (
            in0 => \N__3923\,
            in1 => \N__3407\,
            in2 => \N__3625\,
            in3 => \N__4246\,
            lcout => OPEN,
            ltout => \uart.N_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_3_LC_10_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101001100000011"
        )
    port map (
            in0 => \N__3364\,
            in1 => \N__3311\,
            in2 => \N__3305\,
            in3 => \N__3611\,
            lcout => \uart.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4791\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_esr_3_LC_11_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3742\,
            lcout => \uart_frame_decoder.state_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4802\,
            ce => \N__3809\,
            sr => \N__4693\
        );

    \uart_frame_decoder.state_1_esr_4_LC_11_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3797\,
            lcout => \uart_frame_decoder.state_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4802\,
            ce => \N__3809\,
            sr => \N__4693\
        );

    \uart_frame_decoder.state_1_esr_5_LC_11_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3300\,
            lcout => \uart_frame_decoder.state_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4802\,
            ce => \N__3809\,
            sr => \N__4693\
        );

    \reset_module_System.count_RNIP8RT_10_LC_11_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4582\,
            in2 => \_gnd_net_\,
            in3 => \N__4330\,
            lcout => \reset_module_System.reset6_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_2_LC_11_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3704\,
            in1 => \N__4613\,
            in2 => \N__3682\,
            in3 => \N__4457\,
            lcout => \reset_module_System.countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4797\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_0_LC_11_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111100001111"
        )
    port map (
            in0 => \N__4611\,
            in1 => \N__3678\,
            in2 => \N__4957\,
            in3 => \N__3702\,
            lcout => \reset_module_System.countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4797\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNI10J41_1_LC_11_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__4532\,
            in1 => \N__4430\,
            in2 => \N__4493\,
            in3 => \N__4977\,
            lcout => \reset_module_System.reset6_14\,
            ltout => \reset_module_System.reset6_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.reset_iso_LC_11_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111111111111"
        )
    port map (
            in0 => \N__4610\,
            in1 => \_gnd_net_\,
            in2 => \N__3707\,
            in3 => \N__3701\,
            lcout => \reset_module_System_reset_iso\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4797\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_1_LC_11_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__3703\,
            in1 => \N__4931\,
            in2 => \N__3683\,
            in3 => \N__4612\,
            lcout => \reset_module_System.countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4797\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNICR4G1_12_LC_11_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__4950\,
            in1 => \N__4549\,
            in2 => \N__4514\,
            in3 => \N__4567\,
            lcout => \reset_module_System.reset6_19_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNI97FD_5_LC_11_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4363\,
            in1 => \N__4378\,
            in2 => \N__4349\,
            in3 => \N__4414\,
            lcout => \reset_module_System.reset6_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.bit_Count_RNO_2_1_LC_11_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101110111011"
        )
    port map (
            in0 => \N__4113\,
            in1 => \N__3615\,
            in2 => \N__3560\,
            in3 => \N__3550\,
            lcout => \uart.state_0_sqmuxa_1_d_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNO_5_4_LC_11_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__4162\,
            in1 => \N__4205\,
            in2 => \N__3485\,
            in3 => \N__3997\,
            lcout => OPEN,
            ltout => \uart.g3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNO_0_4_LC_11_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001010101010"
        )
    port map (
            in0 => \N__4211\,
            in1 => \N__4114\,
            in2 => \N__4316\,
            in3 => \N__4305\,
            lcout => \uart.N_167_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNO_4_4_LC_11_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__4235\,
            in1 => \N__3920\,
            in2 => \_gnd_net_\,
            in3 => \N__5042\,
            lcout => \uart.g0_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNO_2_3_LC_11_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__4204\,
            in1 => \N__4161\,
            in2 => \N__4003\,
            in3 => \N__4112\,
            lcout => \uart.state_RNO_2Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_2_rep1_LC_11_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__3998\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4046\,
            lcout => \uart.timer_Count_2_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4792\,
            ce => 'H',
            sr => \N__3973\
        );

    \uart.data_rdy_LC_11_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110000010100000"
        )
    port map (
            in0 => \N__3930\,
            in1 => \N__3860\,
            in2 => \N__4991\,
            in3 => \N__3836\,
            lcout => uart_data_rdy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4789\,
            ce => 'H',
            sr => \N__4706\
        );

    \uart_frame_decoder.state_1_esr_ctle_5_LC_12_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__4692\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4897\,
            lcout => \uart_frame_decoder.uart_data_rdy_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_esr_RNIQ0UJ_3_LC_12_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__3798\,
            in1 => \N__3776\,
            in2 => \_gnd_net_\,
            in3 => \N__3743\,
            lcout => \uart_frame_decoder_N_130_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_1_cry_1_c_LC_12_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4949\,
            in2 => \N__4982\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_2_0_\,
            carryout => \reset_module_System.count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNO_0_2_LC_12_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4469\,
            in2 => \_gnd_net_\,
            in3 => \N__4451\,
            lcout => \reset_module_System.count_1_2\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_1\,
            carryout => \reset_module_System.count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_3_LC_12_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4447\,
            in2 => \_gnd_net_\,
            in3 => \N__4433\,
            lcout => \reset_module_System.countZ0Z_3\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_2\,
            carryout => \reset_module_System.count_1_cry_3\,
            clk => \N__4790\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_4_LC_12_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4429\,
            in2 => \_gnd_net_\,
            in3 => \N__4418\,
            lcout => \reset_module_System.countZ0Z_4\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_3\,
            carryout => \reset_module_System.count_1_cry_4\,
            clk => \N__4790\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_5_LC_12_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4415\,
            in2 => \_gnd_net_\,
            in3 => \N__4403\,
            lcout => \reset_module_System.countZ0Z_5\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_4\,
            carryout => \reset_module_System.count_1_cry_5\,
            clk => \N__4790\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_6_LC_12_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4396\,
            in2 => \_gnd_net_\,
            in3 => \N__4382\,
            lcout => \reset_module_System.countZ0Z_6\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_5\,
            carryout => \reset_module_System.count_1_cry_6\,
            clk => \N__4790\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_7_LC_12_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4379\,
            in2 => \_gnd_net_\,
            in3 => \N__4367\,
            lcout => \reset_module_System.countZ0Z_7\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_6\,
            carryout => \reset_module_System.count_1_cry_7\,
            clk => \N__4790\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_8_LC_12_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4364\,
            in2 => \_gnd_net_\,
            in3 => \N__4352\,
            lcout => \reset_module_System.countZ0Z_8\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_7\,
            carryout => \reset_module_System.count_1_cry_8\,
            clk => \N__4790\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_9_LC_12_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4348\,
            in2 => \_gnd_net_\,
            in3 => \N__4334\,
            lcout => \reset_module_System.countZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_12_3_0_\,
            carryout => \reset_module_System.count_1_cry_9\,
            clk => \N__4788\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_10_LC_12_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4331\,
            in2 => \_gnd_net_\,
            in3 => \N__4319\,
            lcout => \reset_module_System.countZ0Z_10\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_9\,
            carryout => \reset_module_System.count_1_cry_10\,
            clk => \N__4788\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_11_LC_12_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4583\,
            in2 => \_gnd_net_\,
            in3 => \N__4571\,
            lcout => \reset_module_System.countZ0Z_11\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_10\,
            carryout => \reset_module_System.count_1_cry_11\,
            clk => \N__4788\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_12_LC_12_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4568\,
            in2 => \_gnd_net_\,
            in3 => \N__4556\,
            lcout => \reset_module_System.countZ0Z_12\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_11\,
            carryout => \reset_module_System.count_1_cry_12\,
            clk => \N__4788\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_13_LC_12_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4624\,
            in2 => \_gnd_net_\,
            in3 => \N__4553\,
            lcout => \reset_module_System.countZ0Z_13\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_12\,
            carryout => \reset_module_System.count_1_cry_13\,
            clk => \N__4788\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_14_LC_12_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4550\,
            in2 => \_gnd_net_\,
            in3 => \N__4538\,
            lcout => \reset_module_System.countZ0Z_14\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_13\,
            carryout => \reset_module_System.count_1_cry_14\,
            clk => \N__4788\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_15_LC_12_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4651\,
            in2 => \_gnd_net_\,
            in3 => \N__4535\,
            lcout => \reset_module_System.countZ0Z_15\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_14\,
            carryout => \reset_module_System.count_1_cry_15\,
            clk => \N__4788\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_16_LC_12_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4528\,
            in2 => \_gnd_net_\,
            in3 => \N__4517\,
            lcout => \reset_module_System.countZ0Z_16\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_15\,
            carryout => \reset_module_System.count_1_cry_16\,
            clk => \N__4788\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_17_LC_12_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4510\,
            in2 => \_gnd_net_\,
            in3 => \N__4496\,
            lcout => \reset_module_System.countZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_12_4_0_\,
            carryout => \reset_module_System.count_1_cry_17\,
            clk => \N__4787\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_18_LC_12_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4486\,
            in2 => \_gnd_net_\,
            in3 => \N__4472\,
            lcout => \reset_module_System.countZ0Z_18\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_17\,
            carryout => \reset_module_System.count_1_cry_18\,
            clk => \N__4787\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_19_LC_12_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4664\,
            in2 => \_gnd_net_\,
            in3 => \N__5192\,
            lcout => \reset_module_System.countZ0Z_19\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_18\,
            carryout => \reset_module_System.count_1_cry_19\,
            clk => \N__4787\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_20_LC_12_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5182\,
            in2 => \_gnd_net_\,
            in3 => \N__5168\,
            lcout => \reset_module_System.countZ0Z_20\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_19\,
            carryout => \reset_module_System.count_1_cry_20\,
            clk => \N__4787\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_21_LC_12_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4639\,
            in2 => \_gnd_net_\,
            in3 => \N__5165\,
            lcout => \reset_module_System.countZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4787\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_rdy_RNO_0_LC_12_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5155\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5052\,
            lcout => \uart.data_rdyc_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNO_0_1_LC_13_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4981\,
            in2 => \_gnd_net_\,
            in3 => \N__4958\,
            lcout => \reset_module_System.count_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.source_data_valid_LC_13_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4825\,
            in2 => \_gnd_net_\,
            in3 => \N__4916\,
            lcout => frame_decoder_dv_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4793\,
            ce => 'H',
            sr => \N__4716\
        );

    \reset_module_System.count_RNI34OR1_21_LC_13_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4663\,
            in1 => \N__4652\,
            in2 => \N__4640\,
            in3 => \N__4625\,
            lcout => \reset_module_System.reset6_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
