// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     Mar 12 2019 01:42:22

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "Pc2Drone" view "INTERFACE"

module Pc2Drone (
    debug_state_output,
    uart_input,
    uart_data_rdy,
    debug_sinkdatavalid_output,
    uart_input_debug,
    frame_decoder_dv,
    clk_system);

    output [4:0] debug_state_output;
    input uart_input;
    output uart_data_rdy;
    output debug_sinkdatavalid_output;
    output uart_input_debug;
    output frame_decoder_dv;
    input clk_system;

    wire N__5303;
    wire N__5302;
    wire N__5301;
    wire N__5292;
    wire N__5291;
    wire N__5290;
    wire N__5283;
    wire N__5282;
    wire N__5281;
    wire N__5274;
    wire N__5273;
    wire N__5272;
    wire N__5265;
    wire N__5264;
    wire N__5263;
    wire N__5256;
    wire N__5255;
    wire N__5254;
    wire N__5247;
    wire N__5246;
    wire N__5245;
    wire N__5238;
    wire N__5237;
    wire N__5236;
    wire N__5229;
    wire N__5228;
    wire N__5227;
    wire N__5220;
    wire N__5219;
    wire N__5218;
    wire N__5211;
    wire N__5210;
    wire N__5209;
    wire N__5192;
    wire N__5189;
    wire N__5186;
    wire N__5183;
    wire N__5182;
    wire N__5179;
    wire N__5176;
    wire N__5173;
    wire N__5168;
    wire N__5165;
    wire N__5162;
    wire N__5161;
    wire N__5160;
    wire N__5159;
    wire N__5158;
    wire N__5157;
    wire N__5156;
    wire N__5155;
    wire N__5152;
    wire N__5149;
    wire N__5146;
    wire N__5141;
    wire N__5138;
    wire N__5135;
    wire N__5134;
    wire N__5131;
    wire N__5130;
    wire N__5117;
    wire N__5114;
    wire N__5111;
    wire N__5108;
    wire N__5107;
    wire N__5106;
    wire N__5105;
    wire N__5104;
    wire N__5099;
    wire N__5094;
    wire N__5091;
    wire N__5088;
    wire N__5083;
    wire N__5080;
    wire N__5077;
    wire N__5070;
    wire N__5063;
    wire N__5062;
    wire N__5061;
    wire N__5058;
    wire N__5053;
    wire N__5052;
    wire N__5051;
    wire N__5046;
    wire N__5043;
    wire N__5042;
    wire N__5041;
    wire N__5038;
    wire N__5037;
    wire N__5036;
    wire N__5035;
    wire N__5034;
    wire N__5033;
    wire N__5030;
    wire N__5027;
    wire N__5024;
    wire N__5021;
    wire N__5018;
    wire N__5009;
    wire N__5006;
    wire N__4991;
    wire N__4988;
    wire N__4985;
    wire N__4982;
    wire N__4981;
    wire N__4978;
    wire N__4977;
    wire N__4974;
    wire N__4971;
    wire N__4968;
    wire N__4963;
    wire N__4958;
    wire N__4957;
    wire N__4954;
    wire N__4951;
    wire N__4950;
    wire N__4949;
    wire N__4946;
    wire N__4941;
    wire N__4938;
    wire N__4931;
    wire N__4928;
    wire N__4925;
    wire N__4922;
    wire N__4919;
    wire N__4918;
    wire N__4917;
    wire N__4916;
    wire N__4915;
    wire N__4914;
    wire N__4913;
    wire N__4912;
    wire N__4911;
    wire N__4910;
    wire N__4907;
    wire N__4904;
    wire N__4901;
    wire N__4898;
    wire N__4897;
    wire N__4888;
    wire N__4883;
    wire N__4878;
    wire N__4875;
    wire N__4872;
    wire N__4869;
    wire N__4866;
    wire N__4863;
    wire N__4858;
    wire N__4855;
    wire N__4852;
    wire N__4847;
    wire N__4838;
    wire N__4835;
    wire N__4832;
    wire N__4829;
    wire N__4826;
    wire N__4825;
    wire N__4822;
    wire N__4819;
    wire N__4814;
    wire N__4813;
    wire N__4812;
    wire N__4811;
    wire N__4810;
    wire N__4809;
    wire N__4808;
    wire N__4807;
    wire N__4806;
    wire N__4805;
    wire N__4804;
    wire N__4803;
    wire N__4802;
    wire N__4801;
    wire N__4800;
    wire N__4799;
    wire N__4798;
    wire N__4797;
    wire N__4796;
    wire N__4795;
    wire N__4794;
    wire N__4793;
    wire N__4792;
    wire N__4791;
    wire N__4790;
    wire N__4789;
    wire N__4788;
    wire N__4787;
    wire N__4730;
    wire N__4727;
    wire N__4724;
    wire N__4723;
    wire N__4720;
    wire N__4717;
    wire N__4716;
    wire N__4713;
    wire N__4710;
    wire N__4707;
    wire N__4706;
    wire N__4703;
    wire N__4700;
    wire N__4697;
    wire N__4694;
    wire N__4693;
    wire N__4692;
    wire N__4689;
    wire N__4684;
    wire N__4681;
    wire N__4678;
    wire N__4675;
    wire N__4664;
    wire N__4663;
    wire N__4660;
    wire N__4657;
    wire N__4652;
    wire N__4651;
    wire N__4648;
    wire N__4645;
    wire N__4640;
    wire N__4639;
    wire N__4636;
    wire N__4633;
    wire N__4630;
    wire N__4625;
    wire N__4624;
    wire N__4621;
    wire N__4618;
    wire N__4613;
    wire N__4612;
    wire N__4611;
    wire N__4610;
    wire N__4609;
    wire N__4608;
    wire N__4599;
    wire N__4594;
    wire N__4589;
    wire N__4586;
    wire N__4583;
    wire N__4582;
    wire N__4579;
    wire N__4576;
    wire N__4571;
    wire N__4568;
    wire N__4567;
    wire N__4564;
    wire N__4561;
    wire N__4556;
    wire N__4553;
    wire N__4550;
    wire N__4549;
    wire N__4546;
    wire N__4543;
    wire N__4538;
    wire N__4535;
    wire N__4532;
    wire N__4529;
    wire N__4528;
    wire N__4525;
    wire N__4522;
    wire N__4517;
    wire N__4514;
    wire N__4511;
    wire N__4510;
    wire N__4507;
    wire N__4504;
    wire N__4501;
    wire N__4496;
    wire N__4493;
    wire N__4490;
    wire N__4487;
    wire N__4486;
    wire N__4483;
    wire N__4480;
    wire N__4477;
    wire N__4472;
    wire N__4469;
    wire N__4468;
    wire N__4465;
    wire N__4462;
    wire N__4457;
    wire N__4454;
    wire N__4451;
    wire N__4448;
    wire N__4447;
    wire N__4444;
    wire N__4441;
    wire N__4438;
    wire N__4433;
    wire N__4430;
    wire N__4429;
    wire N__4426;
    wire N__4423;
    wire N__4418;
    wire N__4415;
    wire N__4414;
    wire N__4411;
    wire N__4408;
    wire N__4403;
    wire N__4400;
    wire N__4397;
    wire N__4396;
    wire N__4393;
    wire N__4390;
    wire N__4387;
    wire N__4382;
    wire N__4379;
    wire N__4378;
    wire N__4375;
    wire N__4372;
    wire N__4367;
    wire N__4364;
    wire N__4363;
    wire N__4360;
    wire N__4357;
    wire N__4352;
    wire N__4349;
    wire N__4348;
    wire N__4345;
    wire N__4342;
    wire N__4339;
    wire N__4334;
    wire N__4331;
    wire N__4330;
    wire N__4327;
    wire N__4324;
    wire N__4319;
    wire N__4316;
    wire N__4313;
    wire N__4312;
    wire N__4309;
    wire N__4306;
    wire N__4305;
    wire N__4304;
    wire N__4303;
    wire N__4302;
    wire N__4301;
    wire N__4300;
    wire N__4299;
    wire N__4298;
    wire N__4297;
    wire N__4296;
    wire N__4293;
    wire N__4290;
    wire N__4287;
    wire N__4280;
    wire N__4277;
    wire N__4266;
    wire N__4253;
    wire N__4250;
    wire N__4247;
    wire N__4246;
    wire N__4243;
    wire N__4242;
    wire N__4239;
    wire N__4236;
    wire N__4235;
    wire N__4232;
    wire N__4229;
    wire N__4226;
    wire N__4223;
    wire N__4220;
    wire N__4211;
    wire N__4208;
    wire N__4205;
    wire N__4204;
    wire N__4199;
    wire N__4198;
    wire N__4197;
    wire N__4196;
    wire N__4195;
    wire N__4194;
    wire N__4193;
    wire N__4192;
    wire N__4189;
    wire N__4176;
    wire N__4173;
    wire N__4170;
    wire N__4163;
    wire N__4162;
    wire N__4161;
    wire N__4160;
    wire N__4159;
    wire N__4156;
    wire N__4151;
    wire N__4148;
    wire N__4145;
    wire N__4140;
    wire N__4137;
    wire N__4132;
    wire N__4127;
    wire N__4126;
    wire N__4123;
    wire N__4120;
    wire N__4119;
    wire N__4118;
    wire N__4115;
    wire N__4114;
    wire N__4113;
    wire N__4112;
    wire N__4109;
    wire N__4106;
    wire N__4105;
    wire N__4104;
    wire N__4103;
    wire N__4102;
    wire N__4101;
    wire N__4100;
    wire N__4097;
    wire N__4094;
    wire N__4087;
    wire N__4082;
    wire N__4079;
    wire N__4068;
    wire N__4055;
    wire N__4052;
    wire N__4049;
    wire N__4046;
    wire N__4045;
    wire N__4042;
    wire N__4039;
    wire N__4038;
    wire N__4037;
    wire N__4036;
    wire N__4033;
    wire N__4032;
    wire N__4031;
    wire N__4030;
    wire N__4021;
    wire N__4018;
    wire N__4011;
    wire N__4004;
    wire N__4003;
    wire N__4002;
    wire N__3999;
    wire N__3998;
    wire N__3997;
    wire N__3994;
    wire N__3991;
    wire N__3988;
    wire N__3981;
    wire N__3974;
    wire N__3973;
    wire N__3972;
    wire N__3969;
    wire N__3968;
    wire N__3965;
    wire N__3962;
    wire N__3959;
    wire N__3956;
    wire N__3953;
    wire N__3946;
    wire N__3943;
    wire N__3940;
    wire N__3935;
    wire N__3934;
    wire N__3933;
    wire N__3932;
    wire N__3931;
    wire N__3930;
    wire N__3927;
    wire N__3924;
    wire N__3923;
    wire N__3922;
    wire N__3921;
    wire N__3920;
    wire N__3917;
    wire N__3916;
    wire N__3915;
    wire N__3912;
    wire N__3909;
    wire N__3908;
    wire N__3905;
    wire N__3900;
    wire N__3893;
    wire N__3890;
    wire N__3885;
    wire N__3882;
    wire N__3875;
    wire N__3860;
    wire N__3857;
    wire N__3854;
    wire N__3853;
    wire N__3852;
    wire N__3849;
    wire N__3846;
    wire N__3843;
    wire N__3836;
    wire N__3833;
    wire N__3830;
    wire N__3829;
    wire N__3828;
    wire N__3827;
    wire N__3824;
    wire N__3821;
    wire N__3816;
    wire N__3809;
    wire N__3806;
    wire N__3803;
    wire N__3800;
    wire N__3799;
    wire N__3798;
    wire N__3797;
    wire N__3792;
    wire N__3789;
    wire N__3786;
    wire N__3783;
    wire N__3776;
    wire N__3775;
    wire N__3774;
    wire N__3773;
    wire N__3770;
    wire N__3763;
    wire N__3762;
    wire N__3759;
    wire N__3756;
    wire N__3753;
    wire N__3748;
    wire N__3743;
    wire N__3742;
    wire N__3739;
    wire N__3736;
    wire N__3735;
    wire N__3734;
    wire N__3729;
    wire N__3724;
    wire N__3719;
    wire N__3716;
    wire N__3713;
    wire N__3710;
    wire N__3707;
    wire N__3704;
    wire N__3703;
    wire N__3702;
    wire N__3701;
    wire N__3700;
    wire N__3691;
    wire N__3688;
    wire N__3683;
    wire N__3682;
    wire N__3679;
    wire N__3678;
    wire N__3675;
    wire N__3668;
    wire N__3667;
    wire N__3666;
    wire N__3663;
    wire N__3658;
    wire N__3653;
    wire N__3650;
    wire N__3647;
    wire N__3644;
    wire N__3641;
    wire N__3640;
    wire N__3639;
    wire N__3638;
    wire N__3635;
    wire N__3632;
    wire N__3629;
    wire N__3626;
    wire N__3625;
    wire N__3624;
    wire N__3621;
    wire N__3616;
    wire N__3615;
    wire N__3612;
    wire N__3611;
    wire N__3608;
    wire N__3607;
    wire N__3606;
    wire N__3603;
    wire N__3602;
    wire N__3601;
    wire N__3600;
    wire N__3595;
    wire N__3592;
    wire N__3589;
    wire N__3578;
    wire N__3571;
    wire N__3560;
    wire N__3557;
    wire N__3554;
    wire N__3551;
    wire N__3550;
    wire N__3549;
    wire N__3546;
    wire N__3543;
    wire N__3540;
    wire N__3539;
    wire N__3536;
    wire N__3533;
    wire N__3532;
    wire N__3531;
    wire N__3530;
    wire N__3527;
    wire N__3524;
    wire N__3519;
    wire N__3512;
    wire N__3509;
    wire N__3506;
    wire N__3497;
    wire N__3494;
    wire N__3491;
    wire N__3488;
    wire N__3485;
    wire N__3482;
    wire N__3479;
    wire N__3478;
    wire N__3477;
    wire N__3474;
    wire N__3473;
    wire N__3472;
    wire N__3467;
    wire N__3464;
    wire N__3459;
    wire N__3452;
    wire N__3449;
    wire N__3446;
    wire N__3443;
    wire N__3442;
    wire N__3441;
    wire N__3438;
    wire N__3433;
    wire N__3428;
    wire N__3427;
    wire N__3424;
    wire N__3421;
    wire N__3418;
    wire N__3415;
    wire N__3410;
    wire N__3407;
    wire N__3404;
    wire N__3401;
    wire N__3400;
    wire N__3397;
    wire N__3394;
    wire N__3391;
    wire N__3386;
    wire N__3385;
    wire N__3382;
    wire N__3381;
    wire N__3380;
    wire N__3379;
    wire N__3376;
    wire N__3373;
    wire N__3368;
    wire N__3365;
    wire N__3364;
    wire N__3363;
    wire N__3362;
    wire N__3357;
    wire N__3352;
    wire N__3351;
    wire N__3350;
    wire N__3345;
    wire N__3344;
    wire N__3343;
    wire N__3340;
    wire N__3335;
    wire N__3330;
    wire N__3327;
    wire N__3322;
    wire N__3311;
    wire N__3308;
    wire N__3305;
    wire N__3302;
    wire N__3301;
    wire N__3300;
    wire N__3297;
    wire N__3294;
    wire N__3291;
    wire N__3286;
    wire N__3281;
    wire N__3278;
    wire N__3277;
    wire N__3276;
    wire N__3275;
    wire N__3272;
    wire N__3269;
    wire N__3266;
    wire N__3261;
    wire N__3258;
    wire N__3255;
    wire N__3252;
    wire N__3245;
    wire N__3242;
    wire N__3239;
    wire N__3236;
    wire N__3233;
    wire N__3232;
    wire N__3231;
    wire N__3228;
    wire N__3221;
    wire N__3218;
    wire N__3215;
    wire N__3212;
    wire N__3209;
    wire N__3206;
    wire N__3203;
    wire N__3202;
    wire N__3201;
    wire N__3196;
    wire N__3195;
    wire N__3192;
    wire N__3189;
    wire N__3184;
    wire N__3179;
    wire N__3176;
    wire N__3173;
    wire N__3172;
    wire N__3171;
    wire N__3168;
    wire N__3165;
    wire N__3162;
    wire N__3161;
    wire N__3160;
    wire N__3159;
    wire N__3158;
    wire N__3153;
    wire N__3150;
    wire N__3149;
    wire N__3148;
    wire N__3147;
    wire N__3146;
    wire N__3143;
    wire N__3140;
    wire N__3139;
    wire N__3136;
    wire N__3135;
    wire N__3132;
    wire N__3129;
    wire N__3126;
    wire N__3123;
    wire N__3120;
    wire N__3115;
    wire N__3106;
    wire N__3103;
    wire N__3098;
    wire N__3083;
    wire N__3080;
    wire N__3077;
    wire N__3076;
    wire N__3075;
    wire N__3074;
    wire N__3073;
    wire N__3070;
    wire N__3067;
    wire N__3062;
    wire N__3061;
    wire N__3060;
    wire N__3059;
    wire N__3056;
    wire N__3053;
    wire N__3048;
    wire N__3045;
    wire N__3040;
    wire N__3029;
    wire N__3026;
    wire N__3025;
    wire N__3024;
    wire N__3023;
    wire N__3020;
    wire N__3017;
    wire N__3012;
    wire N__3011;
    wire N__3010;
    wire N__3009;
    wire N__3008;
    wire N__3007;
    wire N__3004;
    wire N__2999;
    wire N__2994;
    wire N__2987;
    wire N__2978;
    wire N__2975;
    wire N__2972;
    wire N__2969;
    wire N__2966;
    wire N__2963;
    wire N__2962;
    wire N__2961;
    wire N__2958;
    wire N__2957;
    wire N__2954;
    wire N__2947;
    wire N__2942;
    wire N__2939;
    wire N__2936;
    wire N__2933;
    wire N__2930;
    wire N__2927;
    wire N__2924;
    wire N__2923;
    wire N__2922;
    wire N__2919;
    wire N__2918;
    wire N__2917;
    wire N__2914;
    wire N__2911;
    wire N__2908;
    wire N__2901;
    wire N__2894;
    wire N__2891;
    wire N__2888;
    wire N__2885;
    wire N__2884;
    wire N__2883;
    wire N__2880;
    wire N__2877;
    wire N__2874;
    wire N__2871;
    wire N__2868;
    wire N__2863;
    wire N__2858;
    wire N__2855;
    wire N__2852;
    wire N__2849;
    wire N__2848;
    wire N__2847;
    wire N__2842;
    wire N__2841;
    wire N__2838;
    wire N__2837;
    wire N__2836;
    wire N__2835;
    wire N__2834;
    wire N__2831;
    wire N__2828;
    wire N__2825;
    wire N__2816;
    wire N__2807;
    wire N__2804;
    wire N__2801;
    wire N__2798;
    wire N__2797;
    wire N__2794;
    wire N__2791;
    wire N__2786;
    wire N__2783;
    wire N__2780;
    wire N__2777;
    wire N__2774;
    wire N__2771;
    wire N__2768;
    wire N__2765;
    wire N__2762;
    wire N__2759;
    wire N__2756;
    wire N__2753;
    wire N__2750;
    wire N__2747;
    wire N__2744;
    wire N__2743;
    wire N__2742;
    wire N__2741;
    wire N__2740;
    wire N__2739;
    wire N__2736;
    wire N__2733;
    wire N__2730;
    wire N__2729;
    wire N__2728;
    wire N__2727;
    wire N__2726;
    wire N__2723;
    wire N__2720;
    wire N__2717;
    wire N__2716;
    wire N__2713;
    wire N__2708;
    wire N__2705;
    wire N__2704;
    wire N__2697;
    wire N__2696;
    wire N__2695;
    wire N__2694;
    wire N__2689;
    wire N__2686;
    wire N__2683;
    wire N__2682;
    wire N__2679;
    wire N__2676;
    wire N__2673;
    wire N__2670;
    wire N__2667;
    wire N__2660;
    wire N__2653;
    wire N__2650;
    wire N__2633;
    wire N__2632;
    wire N__2629;
    wire N__2628;
    wire N__2627;
    wire N__2626;
    wire N__2623;
    wire N__2622;
    wire N__2621;
    wire N__2620;
    wire N__2615;
    wire N__2602;
    wire N__2597;
    wire N__2594;
    wire N__2593;
    wire N__2590;
    wire N__2587;
    wire N__2582;
    wire N__2579;
    wire N__2576;
    wire N__2573;
    wire N__2570;
    wire N__2567;
    wire N__2564;
    wire N__2561;
    wire N__2558;
    wire N__2557;
    wire N__2554;
    wire N__2551;
    wire N__2546;
    wire N__2543;
    wire N__2540;
    wire N__2537;
    wire N__2534;
    wire N__2531;
    wire N__2528;
    wire N__2525;
    wire N__2522;
    wire N__2519;
    wire N__2518;
    wire N__2513;
    wire N__2510;
    wire N__2507;
    wire N__2504;
    wire N__2501;
    wire N__2498;
    wire N__2497;
    wire N__2494;
    wire N__2491;
    wire N__2486;
    wire N__2485;
    wire N__2480;
    wire N__2477;
    wire N__2476;
    wire N__2475;
    wire N__2474;
    wire N__2469;
    wire N__2466;
    wire N__2465;
    wire N__2464;
    wire N__2463;
    wire N__2460;
    wire N__2457;
    wire N__2448;
    wire N__2441;
    wire N__2438;
    wire N__2435;
    wire N__2432;
    wire N__2429;
    wire N__2426;
    wire N__2423;
    wire N__2420;
    wire N__2417;
    wire N__2414;
    wire N__2411;
    wire N__2408;
    wire N__2405;
    wire N__2402;
    wire N__2399;
    wire N__2396;
    wire N__2393;
    wire N__2392;
    wire N__2389;
    wire N__2386;
    wire N__2381;
    wire N__2378;
    wire N__2375;
    wire N__2372;
    wire N__2369;
    wire N__2366;
    wire N__2363;
    wire N__2360;
    wire N__2357;
    wire N__2354;
    wire N__2351;
    wire N__2348;
    wire N__2345;
    wire N__2342;
    wire N__2341;
    wire N__2338;
    wire N__2335;
    wire N__2330;
    wire N__2327;
    wire N__2324;
    wire N__2321;
    wire N__2318;
    wire N__2315;
    wire N__2312;
    wire N__2309;
    wire N__2306;
    wire N__2303;
    wire N__2302;
    wire N__2299;
    wire N__2296;
    wire N__2293;
    wire N__2288;
    wire N__2285;
    wire N__2282;
    wire N__2279;
    wire N__2276;
    wire N__2273;
    wire N__2270;
    wire N__2267;
    wire N__2266;
    wire N__2265;
    wire N__2262;
    wire N__2261;
    wire N__2260;
    wire N__2255;
    wire N__2248;
    wire N__2243;
    wire N__2240;
    wire N__2237;
    wire N__2234;
    wire N__2233;
    wire N__2228;
    wire N__2225;
    wire N__2222;
    wire N__2219;
    wire N__2216;
    wire N__2215;
    wire N__2212;
    wire N__2209;
    wire N__2204;
    wire N__2201;
    wire N__2198;
    wire N__2195;
    wire N__2194;
    wire N__2191;
    wire N__2188;
    wire N__2183;
    wire N__2180;
    wire N__2177;
    wire N__2174;
    wire N__2171;
    wire N__2168;
    wire N__2167;
    wire N__2164;
    wire N__2161;
    wire N__2156;
    wire N__2153;
    wire N__2150;
    wire N__2147;
    wire N__2144;
    wire N__2141;
    wire N__2138;
    wire N__2135;
    wire N__2132;
    wire N__2129;
    wire N__2126;
    wire N__2123;
    wire N__2120;
    wire N__2117;
    wire N__2114;
    wire N__2111;
    wire N__2108;
    wire N__2105;
    wire N__2102;
    wire N__2099;
    wire N__2096;
    wire N__2093;
    wire N__2090;
    wire N__2087;
    wire N__2084;
    wire N__2081;
    wire N__2078;
    wire N__2075;
    wire N__2072;
    wire N__2069;
    wire N__2066;
    wire GNDG0;
    wire VCCG0;
    wire \uart_frame_decoder.N_43_cascade_ ;
    wire \uart_frame_decoder.state_1_srsts_i_i_0_0_cascade_ ;
    wire uart_frame_decoder_N_131_i;
    wire \uart_frame_decoder.state_1Z0Z_0 ;
    wire \uart_frame_decoder.state_1_srsts_0_i_1_1 ;
    wire \uart_frame_decoder.N_58_4 ;
    wire \uart_frame_decoder.N_58_4_cascade_ ;
    wire \uart_frame_decoder.N_32_i_1 ;
    wire \uart.state_0_sqmuxa_1_d_cascade_ ;
    wire \uart.m13_0_0_o2_2_cascade_ ;
    wire \uart.N_10_cascade_ ;
    wire \uart.data_Auxce_0_2_cascade_ ;
    wire \uart.data_Aux_esr_RNO_0Z0Z_2_cascade_ ;
    wire \uart.N_118_0 ;
    wire \uart_frame_decoder.state_1_srsts_0_i_a2_0_0_1Z0Z_2_cascade_ ;
    wire \uart_frame_decoder.N_49 ;
    wire \uart_frame_decoder.state_1Z0Z_1 ;
    wire uart_frame_decoder_N_129_i;
    wire \uart_frame_decoder.state_1_srsts_i_i_a2_3_0Z0Z_0_cascade_ ;
    wire \uart_frame_decoder.N_67 ;
    wire \uart_frame_decoder.N_61 ;
    wire \uart_frame_decoder.N_67_cascade_ ;
    wire \uart_frame_decoder.state_1_srsts_0_i_a2_0_0_2 ;
    wire \uart.data_AuxZ0Z_0 ;
    wire uart_data_0;
    wire uart_data_1;
    wire \uart.data_AuxZ0Z_2 ;
    wire uart_data_2;
    wire uart_data_3;
    wire uart_data_4;
    wire uart_data_5;
    wire \uart.data_AuxZ0Z_6 ;
    wire uart_data_6;
    wire \uart.data_AuxZ0Z_7 ;
    wire uart_data_7;
    wire \uart.N_147_0_0_cascade_ ;
    wire \uart.g3_1_0_cascade_ ;
    wire \uart.g0_4_0 ;
    wire \uart.N_175_cascade_ ;
    wire \uart.data_Aux_esr_RNO_0Z0Z_0_cascade_ ;
    wire \uart.N_120_0 ;
    wire \uart.data_Auxce_0_0 ;
    wire \uart.data_Aux_esr_RNO_0Z0Z_1_cascade_ ;
    wire \uart.data_AuxZ0Z_1 ;
    wire \uart.N_119_0 ;
    wire \uart.data_Auxce_0_2 ;
    wire \uart.data_Aux_esr_RNO_0Z0Z_3_cascade_ ;
    wire \uart.data_Aux_esr_RNO_0Z0Z_4_cascade_ ;
    wire \uart.data_Auxce_0_4 ;
    wire \uart.N_113_0 ;
    wire \uart.N_133_0 ;
    wire \uart.stateZ0Z_0 ;
    wire \uart.N_175 ;
    wire \uart.data_Auxce_0_6_cascade_ ;
    wire \uart.N_114_0 ;
    wire \uart.data_Aux_esr_RNO_0Z0Z_5 ;
    wire \uart.data_AuxZ0Z_5 ;
    wire \uart.N_115_0 ;
    wire \uart.un4_timer_Count_1_c2_cascade_ ;
    wire \uart.state_srsts_0_a3_1_4_cascade_ ;
    wire \uart.timer_Count_fastZ0Z_4 ;
    wire \uart.timer_Count10lto4_0 ;
    wire \uart.timer_Count10lto4_0_cascade_ ;
    wire \uart.N_51_cascade_ ;
    wire \uart.N_146_0 ;
    wire \uart.data_14_1_cascade_ ;
    wire \uart.state_RNILS533Z0Z_4 ;
    wire \uart.state_RNILS533Z0Z_4_cascade_ ;
    wire \uart.state_1_sqmuxa_0 ;
    wire \uart.stateZ0Z_1 ;
    wire \uart.N_151 ;
    wire \uart.N_174 ;
    wire \uart.state_srsts_0_a3_2_0_4 ;
    wire \uart.state_1_sqmuxa ;
    wire \uart.data_AuxZ0Z_3 ;
    wire \uart.N_117_0 ;
    wire \uart.data_AuxZ0Z_4 ;
    wire \uart.N_116_0 ;
    wire \uart.state_RNIAFHLZ0Z_4 ;
    wire \uart.timer_CountZ0Z_2 ;
    wire \uart.timer_Count_fastZ0Z_2 ;
    wire \reset_module_System.reset6_11_cascade_ ;
    wire \reset_module_System.reset6_19_cascade_ ;
    wire \uart.N_66 ;
    wire \uart.N_51 ;
    wire \uart.timer_Count_fastZ0Z_3 ;
    wire \uart.N_5 ;
    wire \uart.timer_Count_RNI3B101Z0Z_6 ;
    wire \uart.un4_timer_Count_1_c5 ;
    wire \uart.un1_state_2_0_a3_2 ;
    wire \uart.timer_CountZ0Z_0 ;
    wire \uart.timer_Count_RNI22NA1Z0Z_4 ;
    wire \uart.bit_CountZ0Z_0 ;
    wire \uart.bit_CountZ0Z_2 ;
    wire \uart.bit_CountZ0Z_1 ;
    wire \uart.g1_4_cascade_ ;
    wire \uart.g1_0 ;
    wire \uart.g1_3 ;
    wire \uart.stateZ0Z_2 ;
    wire \uart.un1_state_5 ;
    wire \uart.N_177 ;
    wire reset_system;
    wire \uart.N_28_mux ;
    wire \uart.N_8_cascade_ ;
    wire \uart_frame_decoder.state_1Z0Z_4 ;
    wire \uart_frame_decoder.state_1Z0Z_5 ;
    wire \reset_module_System.reset6_3 ;
    wire \reset_module_System.reset6_14_cascade_ ;
    wire \reset_module_System.reset6_19 ;
    wire \reset_module_System.reset6_14 ;
    wire \reset_module_System.reset6_19_1 ;
    wire \reset_module_System.reset6_13 ;
    wire \uart.stateZ0Z_3 ;
    wire \uart.g3_0_0 ;
    wire \uart.timer_CountZ0Z_4 ;
    wire \uart.state_0_sqmuxa_1_d_0 ;
    wire \uart.timer_CountZ0Z_1 ;
    wire \uart.g3_cascade_ ;
    wire \uart.timer_CountZ0Z_6 ;
    wire \uart.N_167_0 ;
    wire reset_module_System_reset_fast;
    wire \uart.g0_3_1 ;
    wire \uart.timer_CountZ0Z_3 ;
    wire \uart.timer_Count_4_repZ0Z1 ;
    wire \uart.timer_CountZ0Z_5 ;
    wire \uart.state_RNO_2Z0Z_3 ;
    wire \uart.un4_timer_Count_1_c2 ;
    wire \uart.timer_Count_2_repZ0Z1 ;
    wire \uart.state_RNI38F97Z0Z_2 ;
    wire \uart.timer_CountZ0Z_7 ;
    wire \uart.N_41 ;
    wire \uart.state_srsts_0_o4_0_a2_0_4 ;
    wire \uart_frame_decoder.uart_data_rdy_c_0 ;
    wire \uart_frame_decoder.state_1Z0Z_3 ;
    wire \uart_frame_decoder.state_1Z0Z_6 ;
    wire \uart_frame_decoder.state_1Z0Z_2 ;
    wire uart_frame_decoder_N_130_i;
    wire bfn_12_2_0_;
    wire \reset_module_System.countZ0Z_2 ;
    wire \reset_module_System.count_1_2 ;
    wire \reset_module_System.count_1_cry_1 ;
    wire \reset_module_System.countZ0Z_3 ;
    wire \reset_module_System.count_1_cry_2 ;
    wire \reset_module_System.countZ0Z_4 ;
    wire \reset_module_System.count_1_cry_3 ;
    wire \reset_module_System.countZ0Z_5 ;
    wire \reset_module_System.count_1_cry_4 ;
    wire \reset_module_System.countZ0Z_6 ;
    wire \reset_module_System.count_1_cry_5 ;
    wire \reset_module_System.countZ0Z_7 ;
    wire \reset_module_System.count_1_cry_6 ;
    wire \reset_module_System.countZ0Z_8 ;
    wire \reset_module_System.count_1_cry_7 ;
    wire \reset_module_System.count_1_cry_8 ;
    wire \reset_module_System.countZ0Z_9 ;
    wire bfn_12_3_0_;
    wire \reset_module_System.countZ0Z_10 ;
    wire \reset_module_System.count_1_cry_9 ;
    wire \reset_module_System.countZ0Z_11 ;
    wire \reset_module_System.count_1_cry_10 ;
    wire \reset_module_System.countZ0Z_12 ;
    wire \reset_module_System.count_1_cry_11 ;
    wire \reset_module_System.count_1_cry_12 ;
    wire \reset_module_System.countZ0Z_14 ;
    wire \reset_module_System.count_1_cry_13 ;
    wire \reset_module_System.count_1_cry_14 ;
    wire \reset_module_System.countZ0Z_16 ;
    wire \reset_module_System.count_1_cry_15 ;
    wire \reset_module_System.count_1_cry_16 ;
    wire \reset_module_System.countZ0Z_17 ;
    wire bfn_12_4_0_;
    wire \reset_module_System.countZ0Z_18 ;
    wire \reset_module_System.count_1_cry_17 ;
    wire \reset_module_System.count_1_cry_18 ;
    wire \reset_module_System.countZ0Z_20 ;
    wire \reset_module_System.count_1_cry_19 ;
    wire \reset_module_System.count_1_cry_20 ;
    wire uart_input_c;
    wire \uart.stateZ0Z_4 ;
    wire \uart.data_rdyc_0 ;
    wire \reset_module_System.countZ0Z_1 ;
    wire \reset_module_System.countZ0Z_0 ;
    wire \reset_module_System.count_1_1 ;
    wire uart_data_rdy_c;
    wire frame_decoder_dv_c;
    wire clk_system_c_g;
    wire reset_module_System_reset_iso;
    wire \reset_module_System.countZ0Z_19 ;
    wire \reset_module_System.countZ0Z_15 ;
    wire \reset_module_System.countZ0Z_21 ;
    wire \reset_module_System.countZ0Z_13 ;
    wire \reset_module_System.reset6_15 ;
    wire _gnd_net_;

    PRE_IO_GBUF clk_system_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__5301),
            .GLOBALBUFFEROUTPUT(clk_system_c_g));
    defparam clk_system_ibuf_gb_io_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD clk_system_ibuf_gb_io_iopad (
            .OE(N__5303),
            .DIN(N__5302),
            .DOUT(N__5301),
            .PACKAGEPIN(clk_system));
    defparam clk_system_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam clk_system_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_system_ibuf_gb_io_preio (
            .PADOEN(N__5303),
            .PADOUT(N__5302),
            .PADIN(N__5301),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD debug_state_output_obuf_4_iopad (
            .OE(N__5292),
            .DIN(N__5291),
            .DOUT(N__5290),
            .PACKAGEPIN(debug_state_output[4]));
    defparam debug_state_output_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam debug_state_output_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_state_output_obuf_4_preio (
            .PADOEN(N__5292),
            .PADOUT(N__5291),
            .PADIN(N__5290),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_state_output_obuf_1_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_state_output_obuf_1_iopad (
            .OE(N__5283),
            .DIN(N__5282),
            .DOUT(N__5281),
            .PACKAGEPIN(debug_state_output[1]));
    defparam debug_state_output_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam debug_state_output_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_state_output_obuf_1_preio (
            .PADOEN(N__5283),
            .PADOUT(N__5282),
            .PADIN(N__5281),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3719),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam uart_data_rdy_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD uart_data_rdy_obuf_iopad (
            .OE(N__5274),
            .DIN(N__5273),
            .DOUT(N__5272),
            .PACKAGEPIN(uart_data_rdy));
    defparam uart_data_rdy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam uart_data_rdy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO uart_data_rdy_obuf_preio (
            .PADOEN(N__5274),
            .PADOUT(N__5273),
            .PADIN(N__5272),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4922),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_state_output_obuf_3_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_state_output_obuf_3_iopad (
            .OE(N__5265),
            .DIN(N__5264),
            .DOUT(N__5263),
            .PACKAGEPIN(debug_state_output[3]));
    defparam debug_state_output_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam debug_state_output_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_state_output_obuf_3_preio (
            .PADOEN(N__5265),
            .PADOUT(N__5264),
            .PADIN(N__5263),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_sinkdatavalid_output_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_sinkdatavalid_output_obuf_iopad (
            .OE(N__5256),
            .DIN(N__5255),
            .DOUT(N__5254),
            .PACKAGEPIN(debug_sinkdatavalid_output));
    defparam debug_sinkdatavalid_output_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_sinkdatavalid_output_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_sinkdatavalid_output_obuf_preio (
            .PADOEN(N__5256),
            .PADOUT(N__5255),
            .PADIN(N__5254),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4918),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam frame_decoder_dv_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD frame_decoder_dv_obuf_iopad (
            .OE(N__5247),
            .DIN(N__5246),
            .DOUT(N__5245),
            .PACKAGEPIN(frame_decoder_dv));
    defparam frame_decoder_dv_obuf_preio.NEG_TRIGGER=1'b0;
    defparam frame_decoder_dv_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO frame_decoder_dv_obuf_preio (
            .PADOEN(N__5247),
            .PADOUT(N__5246),
            .PADIN(N__5245),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4838),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam uart_input_ibuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD uart_input_ibuf_iopad (
            .OE(N__5238),
            .DIN(N__5237),
            .DOUT(N__5236),
            .PACKAGEPIN(uart_input));
    defparam uart_input_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam uart_input_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO uart_input_ibuf_preio (
            .PADOEN(N__5238),
            .PADOUT(N__5237),
            .PADIN(N__5236),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(uart_input_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_state_output_obuf_0_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_state_output_obuf_0_iopad (
            .OE(N__5229),
            .DIN(N__5228),
            .DOUT(N__5227),
            .PACKAGEPIN(debug_state_output[0]));
    defparam debug_state_output_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam debug_state_output_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_state_output_obuf_0_preio (
            .PADOEN(N__5229),
            .PADOUT(N__5228),
            .PADIN(N__5227),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2243),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_state_output_obuf_2_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_state_output_obuf_2_iopad (
            .OE(N__5220),
            .DIN(N__5219),
            .DOUT(N__5218),
            .PACKAGEPIN(debug_state_output[2]));
    defparam debug_state_output_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam debug_state_output_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_state_output_obuf_2_preio (
            .PADOEN(N__5220),
            .PADOUT(N__5219),
            .PADIN(N__5218),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2096),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam uart_input_debug_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD uart_input_debug_obuf_iopad (
            .OE(N__5211),
            .DIN(N__5210),
            .DOUT(N__5209),
            .PACKAGEPIN(uart_input_debug));
    defparam uart_input_debug_obuf_preio.NEG_TRIGGER=1'b0;
    defparam uart_input_debug_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO uart_input_debug_obuf_preio (
            .PADOEN(N__5211),
            .PADOUT(N__5210),
            .PADIN(N__5209),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5130),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__1217 (
            .O(N__5192),
            .I(\reset_module_System.count_1_cry_18 ));
    CascadeMux I__1216 (
            .O(N__5189),
            .I(N__5186));
    InMux I__1215 (
            .O(N__5186),
            .I(N__5183));
    LocalMux I__1214 (
            .O(N__5183),
            .I(N__5179));
    InMux I__1213 (
            .O(N__5182),
            .I(N__5176));
    Span4Mux_s3_v I__1212 (
            .O(N__5179),
            .I(N__5173));
    LocalMux I__1211 (
            .O(N__5176),
            .I(\reset_module_System.countZ0Z_20 ));
    Odrv4 I__1210 (
            .O(N__5173),
            .I(\reset_module_System.countZ0Z_20 ));
    InMux I__1209 (
            .O(N__5168),
            .I(\reset_module_System.count_1_cry_19 ));
    InMux I__1208 (
            .O(N__5165),
            .I(\reset_module_System.count_1_cry_20 ));
    InMux I__1207 (
            .O(N__5162),
            .I(N__5152));
    InMux I__1206 (
            .O(N__5161),
            .I(N__5149));
    InMux I__1205 (
            .O(N__5160),
            .I(N__5146));
    InMux I__1204 (
            .O(N__5159),
            .I(N__5141));
    InMux I__1203 (
            .O(N__5158),
            .I(N__5141));
    InMux I__1202 (
            .O(N__5157),
            .I(N__5138));
    InMux I__1201 (
            .O(N__5156),
            .I(N__5135));
    InMux I__1200 (
            .O(N__5155),
            .I(N__5131));
    LocalMux I__1199 (
            .O(N__5152),
            .I(N__5117));
    LocalMux I__1198 (
            .O(N__5149),
            .I(N__5117));
    LocalMux I__1197 (
            .O(N__5146),
            .I(N__5117));
    LocalMux I__1196 (
            .O(N__5141),
            .I(N__5117));
    LocalMux I__1195 (
            .O(N__5138),
            .I(N__5117));
    LocalMux I__1194 (
            .O(N__5135),
            .I(N__5117));
    InMux I__1193 (
            .O(N__5134),
            .I(N__5114));
    LocalMux I__1192 (
            .O(N__5131),
            .I(N__5111));
    IoInMux I__1191 (
            .O(N__5130),
            .I(N__5108));
    Span4Mux_v I__1190 (
            .O(N__5117),
            .I(N__5099));
    LocalMux I__1189 (
            .O(N__5114),
            .I(N__5099));
    Span4Mux_v I__1188 (
            .O(N__5111),
            .I(N__5094));
    LocalMux I__1187 (
            .O(N__5108),
            .I(N__5094));
    InMux I__1186 (
            .O(N__5107),
            .I(N__5091));
    InMux I__1185 (
            .O(N__5106),
            .I(N__5088));
    InMux I__1184 (
            .O(N__5105),
            .I(N__5083));
    InMux I__1183 (
            .O(N__5104),
            .I(N__5083));
    IoSpan4Mux I__1182 (
            .O(N__5099),
            .I(N__5080));
    IoSpan4Mux I__1181 (
            .O(N__5094),
            .I(N__5077));
    LocalMux I__1180 (
            .O(N__5091),
            .I(N__5070));
    LocalMux I__1179 (
            .O(N__5088),
            .I(N__5070));
    LocalMux I__1178 (
            .O(N__5083),
            .I(N__5070));
    Odrv4 I__1177 (
            .O(N__5080),
            .I(uart_input_c));
    Odrv4 I__1176 (
            .O(N__5077),
            .I(uart_input_c));
    Odrv12 I__1175 (
            .O(N__5070),
            .I(uart_input_c));
    InMux I__1174 (
            .O(N__5063),
            .I(N__5058));
    InMux I__1173 (
            .O(N__5062),
            .I(N__5053));
    InMux I__1172 (
            .O(N__5061),
            .I(N__5053));
    LocalMux I__1171 (
            .O(N__5058),
            .I(N__5046));
    LocalMux I__1170 (
            .O(N__5053),
            .I(N__5046));
    InMux I__1169 (
            .O(N__5052),
            .I(N__5043));
    InMux I__1168 (
            .O(N__5051),
            .I(N__5038));
    Span4Mux_s3_v I__1167 (
            .O(N__5046),
            .I(N__5030));
    LocalMux I__1166 (
            .O(N__5043),
            .I(N__5027));
    InMux I__1165 (
            .O(N__5042),
            .I(N__5024));
    InMux I__1164 (
            .O(N__5041),
            .I(N__5021));
    LocalMux I__1163 (
            .O(N__5038),
            .I(N__5018));
    InMux I__1162 (
            .O(N__5037),
            .I(N__5009));
    InMux I__1161 (
            .O(N__5036),
            .I(N__5009));
    InMux I__1160 (
            .O(N__5035),
            .I(N__5009));
    InMux I__1159 (
            .O(N__5034),
            .I(N__5009));
    InMux I__1158 (
            .O(N__5033),
            .I(N__5006));
    Odrv4 I__1157 (
            .O(N__5030),
            .I(\uart.stateZ0Z_4 ));
    Odrv4 I__1156 (
            .O(N__5027),
            .I(\uart.stateZ0Z_4 ));
    LocalMux I__1155 (
            .O(N__5024),
            .I(\uart.stateZ0Z_4 ));
    LocalMux I__1154 (
            .O(N__5021),
            .I(\uart.stateZ0Z_4 ));
    Odrv4 I__1153 (
            .O(N__5018),
            .I(\uart.stateZ0Z_4 ));
    LocalMux I__1152 (
            .O(N__5009),
            .I(\uart.stateZ0Z_4 ));
    LocalMux I__1151 (
            .O(N__5006),
            .I(\uart.stateZ0Z_4 ));
    CascadeMux I__1150 (
            .O(N__4991),
            .I(N__4988));
    InMux I__1149 (
            .O(N__4988),
            .I(N__4985));
    LocalMux I__1148 (
            .O(N__4985),
            .I(\uart.data_rdyc_0 ));
    CascadeMux I__1147 (
            .O(N__4982),
            .I(N__4978));
    InMux I__1146 (
            .O(N__4981),
            .I(N__4974));
    InMux I__1145 (
            .O(N__4978),
            .I(N__4971));
    InMux I__1144 (
            .O(N__4977),
            .I(N__4968));
    LocalMux I__1143 (
            .O(N__4974),
            .I(N__4963));
    LocalMux I__1142 (
            .O(N__4971),
            .I(N__4963));
    LocalMux I__1141 (
            .O(N__4968),
            .I(\reset_module_System.countZ0Z_1 ));
    Odrv4 I__1140 (
            .O(N__4963),
            .I(\reset_module_System.countZ0Z_1 ));
    InMux I__1139 (
            .O(N__4958),
            .I(N__4954));
    CascadeMux I__1138 (
            .O(N__4957),
            .I(N__4951));
    LocalMux I__1137 (
            .O(N__4954),
            .I(N__4946));
    InMux I__1136 (
            .O(N__4951),
            .I(N__4941));
    InMux I__1135 (
            .O(N__4950),
            .I(N__4941));
    InMux I__1134 (
            .O(N__4949),
            .I(N__4938));
    Odrv4 I__1133 (
            .O(N__4946),
            .I(\reset_module_System.countZ0Z_0 ));
    LocalMux I__1132 (
            .O(N__4941),
            .I(\reset_module_System.countZ0Z_0 ));
    LocalMux I__1131 (
            .O(N__4938),
            .I(\reset_module_System.countZ0Z_0 ));
    InMux I__1130 (
            .O(N__4931),
            .I(N__4928));
    LocalMux I__1129 (
            .O(N__4928),
            .I(N__4925));
    Odrv4 I__1128 (
            .O(N__4925),
            .I(\reset_module_System.count_1_1 ));
    IoInMux I__1127 (
            .O(N__4922),
            .I(N__4919));
    LocalMux I__1126 (
            .O(N__4919),
            .I(N__4907));
    IoInMux I__1125 (
            .O(N__4918),
            .I(N__4904));
    CascadeMux I__1124 (
            .O(N__4917),
            .I(N__4901));
    InMux I__1123 (
            .O(N__4916),
            .I(N__4898));
    InMux I__1122 (
            .O(N__4915),
            .I(N__4888));
    InMux I__1121 (
            .O(N__4914),
            .I(N__4888));
    InMux I__1120 (
            .O(N__4913),
            .I(N__4888));
    InMux I__1119 (
            .O(N__4912),
            .I(N__4888));
    InMux I__1118 (
            .O(N__4911),
            .I(N__4883));
    InMux I__1117 (
            .O(N__4910),
            .I(N__4883));
    IoSpan4Mux I__1116 (
            .O(N__4907),
            .I(N__4878));
    LocalMux I__1115 (
            .O(N__4904),
            .I(N__4878));
    InMux I__1114 (
            .O(N__4901),
            .I(N__4875));
    LocalMux I__1113 (
            .O(N__4898),
            .I(N__4872));
    InMux I__1112 (
            .O(N__4897),
            .I(N__4869));
    LocalMux I__1111 (
            .O(N__4888),
            .I(N__4866));
    LocalMux I__1110 (
            .O(N__4883),
            .I(N__4863));
    IoSpan4Mux I__1109 (
            .O(N__4878),
            .I(N__4858));
    LocalMux I__1108 (
            .O(N__4875),
            .I(N__4858));
    Span4Mux_s3_v I__1107 (
            .O(N__4872),
            .I(N__4855));
    LocalMux I__1106 (
            .O(N__4869),
            .I(N__4852));
    Span4Mux_h I__1105 (
            .O(N__4866),
            .I(N__4847));
    Span4Mux_h I__1104 (
            .O(N__4863),
            .I(N__4847));
    Odrv4 I__1103 (
            .O(N__4858),
            .I(uart_data_rdy_c));
    Odrv4 I__1102 (
            .O(N__4855),
            .I(uart_data_rdy_c));
    Odrv4 I__1101 (
            .O(N__4852),
            .I(uart_data_rdy_c));
    Odrv4 I__1100 (
            .O(N__4847),
            .I(uart_data_rdy_c));
    IoInMux I__1099 (
            .O(N__4838),
            .I(N__4835));
    LocalMux I__1098 (
            .O(N__4835),
            .I(N__4832));
    IoSpan4Mux I__1097 (
            .O(N__4832),
            .I(N__4829));
    Span4Mux_s2_v I__1096 (
            .O(N__4829),
            .I(N__4826));
    Span4Mux_h I__1095 (
            .O(N__4826),
            .I(N__4822));
    InMux I__1094 (
            .O(N__4825),
            .I(N__4819));
    Odrv4 I__1093 (
            .O(N__4822),
            .I(frame_decoder_dv_c));
    LocalMux I__1092 (
            .O(N__4819),
            .I(frame_decoder_dv_c));
    ClkMux I__1091 (
            .O(N__4814),
            .I(N__4730));
    ClkMux I__1090 (
            .O(N__4813),
            .I(N__4730));
    ClkMux I__1089 (
            .O(N__4812),
            .I(N__4730));
    ClkMux I__1088 (
            .O(N__4811),
            .I(N__4730));
    ClkMux I__1087 (
            .O(N__4810),
            .I(N__4730));
    ClkMux I__1086 (
            .O(N__4809),
            .I(N__4730));
    ClkMux I__1085 (
            .O(N__4808),
            .I(N__4730));
    ClkMux I__1084 (
            .O(N__4807),
            .I(N__4730));
    ClkMux I__1083 (
            .O(N__4806),
            .I(N__4730));
    ClkMux I__1082 (
            .O(N__4805),
            .I(N__4730));
    ClkMux I__1081 (
            .O(N__4804),
            .I(N__4730));
    ClkMux I__1080 (
            .O(N__4803),
            .I(N__4730));
    ClkMux I__1079 (
            .O(N__4802),
            .I(N__4730));
    ClkMux I__1078 (
            .O(N__4801),
            .I(N__4730));
    ClkMux I__1077 (
            .O(N__4800),
            .I(N__4730));
    ClkMux I__1076 (
            .O(N__4799),
            .I(N__4730));
    ClkMux I__1075 (
            .O(N__4798),
            .I(N__4730));
    ClkMux I__1074 (
            .O(N__4797),
            .I(N__4730));
    ClkMux I__1073 (
            .O(N__4796),
            .I(N__4730));
    ClkMux I__1072 (
            .O(N__4795),
            .I(N__4730));
    ClkMux I__1071 (
            .O(N__4794),
            .I(N__4730));
    ClkMux I__1070 (
            .O(N__4793),
            .I(N__4730));
    ClkMux I__1069 (
            .O(N__4792),
            .I(N__4730));
    ClkMux I__1068 (
            .O(N__4791),
            .I(N__4730));
    ClkMux I__1067 (
            .O(N__4790),
            .I(N__4730));
    ClkMux I__1066 (
            .O(N__4789),
            .I(N__4730));
    ClkMux I__1065 (
            .O(N__4788),
            .I(N__4730));
    ClkMux I__1064 (
            .O(N__4787),
            .I(N__4730));
    GlobalMux I__1063 (
            .O(N__4730),
            .I(N__4727));
    gio2CtrlBuf I__1062 (
            .O(N__4727),
            .I(clk_system_c_g));
    SRMux I__1061 (
            .O(N__4724),
            .I(N__4720));
    SRMux I__1060 (
            .O(N__4723),
            .I(N__4717));
    LocalMux I__1059 (
            .O(N__4720),
            .I(N__4713));
    LocalMux I__1058 (
            .O(N__4717),
            .I(N__4710));
    SRMux I__1057 (
            .O(N__4716),
            .I(N__4707));
    Span4Mux_v I__1056 (
            .O(N__4713),
            .I(N__4703));
    Span4Mux_v I__1055 (
            .O(N__4710),
            .I(N__4700));
    LocalMux I__1054 (
            .O(N__4707),
            .I(N__4697));
    SRMux I__1053 (
            .O(N__4706),
            .I(N__4694));
    Span4Mux_h I__1052 (
            .O(N__4703),
            .I(N__4689));
    Span4Mux_s1_v I__1051 (
            .O(N__4700),
            .I(N__4684));
    Span4Mux_v I__1050 (
            .O(N__4697),
            .I(N__4684));
    LocalMux I__1049 (
            .O(N__4694),
            .I(N__4681));
    SRMux I__1048 (
            .O(N__4693),
            .I(N__4678));
    InMux I__1047 (
            .O(N__4692),
            .I(N__4675));
    Odrv4 I__1046 (
            .O(N__4689),
            .I(reset_module_System_reset_iso));
    Odrv4 I__1045 (
            .O(N__4684),
            .I(reset_module_System_reset_iso));
    Odrv12 I__1044 (
            .O(N__4681),
            .I(reset_module_System_reset_iso));
    LocalMux I__1043 (
            .O(N__4678),
            .I(reset_module_System_reset_iso));
    LocalMux I__1042 (
            .O(N__4675),
            .I(reset_module_System_reset_iso));
    InMux I__1041 (
            .O(N__4664),
            .I(N__4660));
    InMux I__1040 (
            .O(N__4663),
            .I(N__4657));
    LocalMux I__1039 (
            .O(N__4660),
            .I(\reset_module_System.countZ0Z_19 ));
    LocalMux I__1038 (
            .O(N__4657),
            .I(\reset_module_System.countZ0Z_19 ));
    InMux I__1037 (
            .O(N__4652),
            .I(N__4648));
    InMux I__1036 (
            .O(N__4651),
            .I(N__4645));
    LocalMux I__1035 (
            .O(N__4648),
            .I(\reset_module_System.countZ0Z_15 ));
    LocalMux I__1034 (
            .O(N__4645),
            .I(\reset_module_System.countZ0Z_15 ));
    CascadeMux I__1033 (
            .O(N__4640),
            .I(N__4636));
    InMux I__1032 (
            .O(N__4639),
            .I(N__4633));
    InMux I__1031 (
            .O(N__4636),
            .I(N__4630));
    LocalMux I__1030 (
            .O(N__4633),
            .I(\reset_module_System.countZ0Z_21 ));
    LocalMux I__1029 (
            .O(N__4630),
            .I(\reset_module_System.countZ0Z_21 ));
    InMux I__1028 (
            .O(N__4625),
            .I(N__4621));
    InMux I__1027 (
            .O(N__4624),
            .I(N__4618));
    LocalMux I__1026 (
            .O(N__4621),
            .I(\reset_module_System.countZ0Z_13 ));
    LocalMux I__1025 (
            .O(N__4618),
            .I(\reset_module_System.countZ0Z_13 ));
    InMux I__1024 (
            .O(N__4613),
            .I(N__4599));
    InMux I__1023 (
            .O(N__4612),
            .I(N__4599));
    InMux I__1022 (
            .O(N__4611),
            .I(N__4599));
    InMux I__1021 (
            .O(N__4610),
            .I(N__4599));
    InMux I__1020 (
            .O(N__4609),
            .I(N__4594));
    InMux I__1019 (
            .O(N__4608),
            .I(N__4594));
    LocalMux I__1018 (
            .O(N__4599),
            .I(N__4589));
    LocalMux I__1017 (
            .O(N__4594),
            .I(N__4589));
    Span4Mux_h I__1016 (
            .O(N__4589),
            .I(N__4586));
    Odrv4 I__1015 (
            .O(N__4586),
            .I(\reset_module_System.reset6_15 ));
    InMux I__1014 (
            .O(N__4583),
            .I(N__4579));
    InMux I__1013 (
            .O(N__4582),
            .I(N__4576));
    LocalMux I__1012 (
            .O(N__4579),
            .I(\reset_module_System.countZ0Z_11 ));
    LocalMux I__1011 (
            .O(N__4576),
            .I(\reset_module_System.countZ0Z_11 ));
    InMux I__1010 (
            .O(N__4571),
            .I(\reset_module_System.count_1_cry_10 ));
    InMux I__1009 (
            .O(N__4568),
            .I(N__4564));
    InMux I__1008 (
            .O(N__4567),
            .I(N__4561));
    LocalMux I__1007 (
            .O(N__4564),
            .I(\reset_module_System.countZ0Z_12 ));
    LocalMux I__1006 (
            .O(N__4561),
            .I(\reset_module_System.countZ0Z_12 ));
    InMux I__1005 (
            .O(N__4556),
            .I(\reset_module_System.count_1_cry_11 ));
    InMux I__1004 (
            .O(N__4553),
            .I(\reset_module_System.count_1_cry_12 ));
    InMux I__1003 (
            .O(N__4550),
            .I(N__4546));
    InMux I__1002 (
            .O(N__4549),
            .I(N__4543));
    LocalMux I__1001 (
            .O(N__4546),
            .I(\reset_module_System.countZ0Z_14 ));
    LocalMux I__1000 (
            .O(N__4543),
            .I(\reset_module_System.countZ0Z_14 ));
    InMux I__999 (
            .O(N__4538),
            .I(\reset_module_System.count_1_cry_13 ));
    InMux I__998 (
            .O(N__4535),
            .I(\reset_module_System.count_1_cry_14 ));
    InMux I__997 (
            .O(N__4532),
            .I(N__4529));
    LocalMux I__996 (
            .O(N__4529),
            .I(N__4525));
    InMux I__995 (
            .O(N__4528),
            .I(N__4522));
    Odrv4 I__994 (
            .O(N__4525),
            .I(\reset_module_System.countZ0Z_16 ));
    LocalMux I__993 (
            .O(N__4522),
            .I(\reset_module_System.countZ0Z_16 ));
    InMux I__992 (
            .O(N__4517),
            .I(\reset_module_System.count_1_cry_15 ));
    CascadeMux I__991 (
            .O(N__4514),
            .I(N__4511));
    InMux I__990 (
            .O(N__4511),
            .I(N__4507));
    InMux I__989 (
            .O(N__4510),
            .I(N__4504));
    LocalMux I__988 (
            .O(N__4507),
            .I(N__4501));
    LocalMux I__987 (
            .O(N__4504),
            .I(\reset_module_System.countZ0Z_17 ));
    Odrv4 I__986 (
            .O(N__4501),
            .I(\reset_module_System.countZ0Z_17 ));
    InMux I__985 (
            .O(N__4496),
            .I(bfn_12_4_0_));
    CascadeMux I__984 (
            .O(N__4493),
            .I(N__4490));
    InMux I__983 (
            .O(N__4490),
            .I(N__4487));
    LocalMux I__982 (
            .O(N__4487),
            .I(N__4483));
    InMux I__981 (
            .O(N__4486),
            .I(N__4480));
    Span4Mux_s1_v I__980 (
            .O(N__4483),
            .I(N__4477));
    LocalMux I__979 (
            .O(N__4480),
            .I(\reset_module_System.countZ0Z_18 ));
    Odrv4 I__978 (
            .O(N__4477),
            .I(\reset_module_System.countZ0Z_18 ));
    InMux I__977 (
            .O(N__4472),
            .I(\reset_module_System.count_1_cry_17 ));
    InMux I__976 (
            .O(N__4469),
            .I(N__4465));
    InMux I__975 (
            .O(N__4468),
            .I(N__4462));
    LocalMux I__974 (
            .O(N__4465),
            .I(\reset_module_System.countZ0Z_2 ));
    LocalMux I__973 (
            .O(N__4462),
            .I(\reset_module_System.countZ0Z_2 ));
    InMux I__972 (
            .O(N__4457),
            .I(N__4454));
    LocalMux I__971 (
            .O(N__4454),
            .I(\reset_module_System.count_1_2 ));
    InMux I__970 (
            .O(N__4451),
            .I(\reset_module_System.count_1_cry_1 ));
    InMux I__969 (
            .O(N__4448),
            .I(N__4444));
    InMux I__968 (
            .O(N__4447),
            .I(N__4441));
    LocalMux I__967 (
            .O(N__4444),
            .I(N__4438));
    LocalMux I__966 (
            .O(N__4441),
            .I(\reset_module_System.countZ0Z_3 ));
    Odrv4 I__965 (
            .O(N__4438),
            .I(\reset_module_System.countZ0Z_3 ));
    InMux I__964 (
            .O(N__4433),
            .I(\reset_module_System.count_1_cry_2 ));
    InMux I__963 (
            .O(N__4430),
            .I(N__4426));
    InMux I__962 (
            .O(N__4429),
            .I(N__4423));
    LocalMux I__961 (
            .O(N__4426),
            .I(\reset_module_System.countZ0Z_4 ));
    LocalMux I__960 (
            .O(N__4423),
            .I(\reset_module_System.countZ0Z_4 ));
    InMux I__959 (
            .O(N__4418),
            .I(\reset_module_System.count_1_cry_3 ));
    InMux I__958 (
            .O(N__4415),
            .I(N__4411));
    InMux I__957 (
            .O(N__4414),
            .I(N__4408));
    LocalMux I__956 (
            .O(N__4411),
            .I(\reset_module_System.countZ0Z_5 ));
    LocalMux I__955 (
            .O(N__4408),
            .I(\reset_module_System.countZ0Z_5 ));
    InMux I__954 (
            .O(N__4403),
            .I(\reset_module_System.count_1_cry_4 ));
    InMux I__953 (
            .O(N__4400),
            .I(N__4397));
    LocalMux I__952 (
            .O(N__4397),
            .I(N__4393));
    InMux I__951 (
            .O(N__4396),
            .I(N__4390));
    Span4Mux_s1_v I__950 (
            .O(N__4393),
            .I(N__4387));
    LocalMux I__949 (
            .O(N__4390),
            .I(\reset_module_System.countZ0Z_6 ));
    Odrv4 I__948 (
            .O(N__4387),
            .I(\reset_module_System.countZ0Z_6 ));
    InMux I__947 (
            .O(N__4382),
            .I(\reset_module_System.count_1_cry_5 ));
    InMux I__946 (
            .O(N__4379),
            .I(N__4375));
    InMux I__945 (
            .O(N__4378),
            .I(N__4372));
    LocalMux I__944 (
            .O(N__4375),
            .I(\reset_module_System.countZ0Z_7 ));
    LocalMux I__943 (
            .O(N__4372),
            .I(\reset_module_System.countZ0Z_7 ));
    InMux I__942 (
            .O(N__4367),
            .I(\reset_module_System.count_1_cry_6 ));
    InMux I__941 (
            .O(N__4364),
            .I(N__4360));
    InMux I__940 (
            .O(N__4363),
            .I(N__4357));
    LocalMux I__939 (
            .O(N__4360),
            .I(\reset_module_System.countZ0Z_8 ));
    LocalMux I__938 (
            .O(N__4357),
            .I(\reset_module_System.countZ0Z_8 ));
    InMux I__937 (
            .O(N__4352),
            .I(\reset_module_System.count_1_cry_7 ));
    CascadeMux I__936 (
            .O(N__4349),
            .I(N__4345));
    InMux I__935 (
            .O(N__4348),
            .I(N__4342));
    InMux I__934 (
            .O(N__4345),
            .I(N__4339));
    LocalMux I__933 (
            .O(N__4342),
            .I(\reset_module_System.countZ0Z_9 ));
    LocalMux I__932 (
            .O(N__4339),
            .I(\reset_module_System.countZ0Z_9 ));
    InMux I__931 (
            .O(N__4334),
            .I(bfn_12_3_0_));
    InMux I__930 (
            .O(N__4331),
            .I(N__4327));
    InMux I__929 (
            .O(N__4330),
            .I(N__4324));
    LocalMux I__928 (
            .O(N__4327),
            .I(\reset_module_System.countZ0Z_10 ));
    LocalMux I__927 (
            .O(N__4324),
            .I(\reset_module_System.countZ0Z_10 ));
    InMux I__926 (
            .O(N__4319),
            .I(\reset_module_System.count_1_cry_9 ));
    CascadeMux I__925 (
            .O(N__4316),
            .I(\uart.g3_cascade_ ));
    InMux I__924 (
            .O(N__4313),
            .I(N__4309));
    InMux I__923 (
            .O(N__4312),
            .I(N__4306));
    LocalMux I__922 (
            .O(N__4309),
            .I(N__4293));
    LocalMux I__921 (
            .O(N__4306),
            .I(N__4290));
    InMux I__920 (
            .O(N__4305),
            .I(N__4287));
    InMux I__919 (
            .O(N__4304),
            .I(N__4280));
    InMux I__918 (
            .O(N__4303),
            .I(N__4280));
    InMux I__917 (
            .O(N__4302),
            .I(N__4280));
    InMux I__916 (
            .O(N__4301),
            .I(N__4277));
    InMux I__915 (
            .O(N__4300),
            .I(N__4266));
    InMux I__914 (
            .O(N__4299),
            .I(N__4266));
    InMux I__913 (
            .O(N__4298),
            .I(N__4266));
    InMux I__912 (
            .O(N__4297),
            .I(N__4266));
    InMux I__911 (
            .O(N__4296),
            .I(N__4266));
    Odrv4 I__910 (
            .O(N__4293),
            .I(\uart.timer_CountZ0Z_6 ));
    Odrv4 I__909 (
            .O(N__4290),
            .I(\uart.timer_CountZ0Z_6 ));
    LocalMux I__908 (
            .O(N__4287),
            .I(\uart.timer_CountZ0Z_6 ));
    LocalMux I__907 (
            .O(N__4280),
            .I(\uart.timer_CountZ0Z_6 ));
    LocalMux I__906 (
            .O(N__4277),
            .I(\uart.timer_CountZ0Z_6 ));
    LocalMux I__905 (
            .O(N__4266),
            .I(\uart.timer_CountZ0Z_6 ));
    InMux I__904 (
            .O(N__4253),
            .I(N__4250));
    LocalMux I__903 (
            .O(N__4250),
            .I(\uart.N_167_0 ));
    InMux I__902 (
            .O(N__4247),
            .I(N__4243));
    InMux I__901 (
            .O(N__4246),
            .I(N__4239));
    LocalMux I__900 (
            .O(N__4243),
            .I(N__4236));
    CascadeMux I__899 (
            .O(N__4242),
            .I(N__4232));
    LocalMux I__898 (
            .O(N__4239),
            .I(N__4229));
    Span4Mux_s1_v I__897 (
            .O(N__4236),
            .I(N__4226));
    InMux I__896 (
            .O(N__4235),
            .I(N__4223));
    InMux I__895 (
            .O(N__4232),
            .I(N__4220));
    Odrv4 I__894 (
            .O(N__4229),
            .I(reset_module_System_reset_fast));
    Odrv4 I__893 (
            .O(N__4226),
            .I(reset_module_System_reset_fast));
    LocalMux I__892 (
            .O(N__4223),
            .I(reset_module_System_reset_fast));
    LocalMux I__891 (
            .O(N__4220),
            .I(reset_module_System_reset_fast));
    InMux I__890 (
            .O(N__4211),
            .I(N__4208));
    LocalMux I__889 (
            .O(N__4208),
            .I(\uart.g0_3_1 ));
    InMux I__888 (
            .O(N__4205),
            .I(N__4199));
    InMux I__887 (
            .O(N__4204),
            .I(N__4199));
    LocalMux I__886 (
            .O(N__4199),
            .I(N__4189));
    InMux I__885 (
            .O(N__4198),
            .I(N__4176));
    InMux I__884 (
            .O(N__4197),
            .I(N__4176));
    InMux I__883 (
            .O(N__4196),
            .I(N__4176));
    InMux I__882 (
            .O(N__4195),
            .I(N__4176));
    InMux I__881 (
            .O(N__4194),
            .I(N__4176));
    InMux I__880 (
            .O(N__4193),
            .I(N__4176));
    InMux I__879 (
            .O(N__4192),
            .I(N__4173));
    Span4Mux_h I__878 (
            .O(N__4189),
            .I(N__4170));
    LocalMux I__877 (
            .O(N__4176),
            .I(\uart.timer_CountZ0Z_3 ));
    LocalMux I__876 (
            .O(N__4173),
            .I(\uart.timer_CountZ0Z_3 ));
    Odrv4 I__875 (
            .O(N__4170),
            .I(\uart.timer_CountZ0Z_3 ));
    InMux I__874 (
            .O(N__4163),
            .I(N__4156));
    InMux I__873 (
            .O(N__4162),
            .I(N__4151));
    InMux I__872 (
            .O(N__4161),
            .I(N__4151));
    CascadeMux I__871 (
            .O(N__4160),
            .I(N__4148));
    InMux I__870 (
            .O(N__4159),
            .I(N__4145));
    LocalMux I__869 (
            .O(N__4156),
            .I(N__4140));
    LocalMux I__868 (
            .O(N__4151),
            .I(N__4140));
    InMux I__867 (
            .O(N__4148),
            .I(N__4137));
    LocalMux I__866 (
            .O(N__4145),
            .I(N__4132));
    Span4Mux_h I__865 (
            .O(N__4140),
            .I(N__4132));
    LocalMux I__864 (
            .O(N__4137),
            .I(\uart.timer_Count_4_repZ0Z1 ));
    Odrv4 I__863 (
            .O(N__4132),
            .I(\uart.timer_Count_4_repZ0Z1 ));
    CascadeMux I__862 (
            .O(N__4127),
            .I(N__4123));
    InMux I__861 (
            .O(N__4126),
            .I(N__4120));
    InMux I__860 (
            .O(N__4123),
            .I(N__4115));
    LocalMux I__859 (
            .O(N__4120),
            .I(N__4109));
    InMux I__858 (
            .O(N__4119),
            .I(N__4106));
    InMux I__857 (
            .O(N__4118),
            .I(N__4097));
    LocalMux I__856 (
            .O(N__4115),
            .I(N__4094));
    InMux I__855 (
            .O(N__4114),
            .I(N__4087));
    InMux I__854 (
            .O(N__4113),
            .I(N__4087));
    InMux I__853 (
            .O(N__4112),
            .I(N__4087));
    Span4Mux_h I__852 (
            .O(N__4109),
            .I(N__4082));
    LocalMux I__851 (
            .O(N__4106),
            .I(N__4082));
    InMux I__850 (
            .O(N__4105),
            .I(N__4079));
    InMux I__849 (
            .O(N__4104),
            .I(N__4068));
    InMux I__848 (
            .O(N__4103),
            .I(N__4068));
    InMux I__847 (
            .O(N__4102),
            .I(N__4068));
    InMux I__846 (
            .O(N__4101),
            .I(N__4068));
    InMux I__845 (
            .O(N__4100),
            .I(N__4068));
    LocalMux I__844 (
            .O(N__4097),
            .I(\uart.timer_CountZ0Z_5 ));
    Odrv4 I__843 (
            .O(N__4094),
            .I(\uart.timer_CountZ0Z_5 ));
    LocalMux I__842 (
            .O(N__4087),
            .I(\uart.timer_CountZ0Z_5 ));
    Odrv4 I__841 (
            .O(N__4082),
            .I(\uart.timer_CountZ0Z_5 ));
    LocalMux I__840 (
            .O(N__4079),
            .I(\uart.timer_CountZ0Z_5 ));
    LocalMux I__839 (
            .O(N__4068),
            .I(\uart.timer_CountZ0Z_5 ));
    CascadeMux I__838 (
            .O(N__4055),
            .I(N__4052));
    InMux I__837 (
            .O(N__4052),
            .I(N__4049));
    LocalMux I__836 (
            .O(N__4049),
            .I(\uart.state_RNO_2Z0Z_3 ));
    InMux I__835 (
            .O(N__4046),
            .I(N__4042));
    CascadeMux I__834 (
            .O(N__4045),
            .I(N__4039));
    LocalMux I__833 (
            .O(N__4042),
            .I(N__4033));
    InMux I__832 (
            .O(N__4039),
            .I(N__4021));
    InMux I__831 (
            .O(N__4038),
            .I(N__4021));
    InMux I__830 (
            .O(N__4037),
            .I(N__4021));
    InMux I__829 (
            .O(N__4036),
            .I(N__4021));
    Span4Mux_h I__828 (
            .O(N__4033),
            .I(N__4018));
    InMux I__827 (
            .O(N__4032),
            .I(N__4011));
    InMux I__826 (
            .O(N__4031),
            .I(N__4011));
    InMux I__825 (
            .O(N__4030),
            .I(N__4011));
    LocalMux I__824 (
            .O(N__4021),
            .I(\uart.un4_timer_Count_1_c2 ));
    Odrv4 I__823 (
            .O(N__4018),
            .I(\uart.un4_timer_Count_1_c2 ));
    LocalMux I__822 (
            .O(N__4011),
            .I(\uart.un4_timer_Count_1_c2 ));
    CascadeMux I__821 (
            .O(N__4004),
            .I(N__3999));
    CascadeMux I__820 (
            .O(N__4003),
            .I(N__3994));
    InMux I__819 (
            .O(N__4002),
            .I(N__3991));
    InMux I__818 (
            .O(N__3999),
            .I(N__3988));
    InMux I__817 (
            .O(N__3998),
            .I(N__3981));
    InMux I__816 (
            .O(N__3997),
            .I(N__3981));
    InMux I__815 (
            .O(N__3994),
            .I(N__3981));
    LocalMux I__814 (
            .O(N__3991),
            .I(\uart.timer_Count_2_repZ0Z1 ));
    LocalMux I__813 (
            .O(N__3988),
            .I(\uart.timer_Count_2_repZ0Z1 ));
    LocalMux I__812 (
            .O(N__3981),
            .I(\uart.timer_Count_2_repZ0Z1 ));
    SRMux I__811 (
            .O(N__3974),
            .I(N__3969));
    SRMux I__810 (
            .O(N__3973),
            .I(N__3965));
    SRMux I__809 (
            .O(N__3972),
            .I(N__3962));
    LocalMux I__808 (
            .O(N__3969),
            .I(N__3959));
    SRMux I__807 (
            .O(N__3968),
            .I(N__3956));
    LocalMux I__806 (
            .O(N__3965),
            .I(N__3953));
    LocalMux I__805 (
            .O(N__3962),
            .I(N__3946));
    Span4Mux_v I__804 (
            .O(N__3959),
            .I(N__3946));
    LocalMux I__803 (
            .O(N__3956),
            .I(N__3946));
    Span4Mux_v I__802 (
            .O(N__3953),
            .I(N__3943));
    Span4Mux_s0_v I__801 (
            .O(N__3946),
            .I(N__3940));
    Odrv4 I__800 (
            .O(N__3943),
            .I(\uart.state_RNI38F97Z0Z_2 ));
    Odrv4 I__799 (
            .O(N__3940),
            .I(\uart.state_RNI38F97Z0Z_2 ));
    InMux I__798 (
            .O(N__3935),
            .I(N__3927));
    InMux I__797 (
            .O(N__3934),
            .I(N__3924));
    CascadeMux I__796 (
            .O(N__3933),
            .I(N__3917));
    CascadeMux I__795 (
            .O(N__3932),
            .I(N__3912));
    CascadeMux I__794 (
            .O(N__3931),
            .I(N__3909));
    InMux I__793 (
            .O(N__3930),
            .I(N__3905));
    LocalMux I__792 (
            .O(N__3927),
            .I(N__3900));
    LocalMux I__791 (
            .O(N__3924),
            .I(N__3900));
    InMux I__790 (
            .O(N__3923),
            .I(N__3893));
    InMux I__789 (
            .O(N__3922),
            .I(N__3893));
    InMux I__788 (
            .O(N__3921),
            .I(N__3893));
    InMux I__787 (
            .O(N__3920),
            .I(N__3890));
    InMux I__786 (
            .O(N__3917),
            .I(N__3885));
    InMux I__785 (
            .O(N__3916),
            .I(N__3885));
    InMux I__784 (
            .O(N__3915),
            .I(N__3882));
    InMux I__783 (
            .O(N__3912),
            .I(N__3875));
    InMux I__782 (
            .O(N__3909),
            .I(N__3875));
    InMux I__781 (
            .O(N__3908),
            .I(N__3875));
    LocalMux I__780 (
            .O(N__3905),
            .I(\uart.timer_CountZ0Z_7 ));
    Odrv4 I__779 (
            .O(N__3900),
            .I(\uart.timer_CountZ0Z_7 ));
    LocalMux I__778 (
            .O(N__3893),
            .I(\uart.timer_CountZ0Z_7 ));
    LocalMux I__777 (
            .O(N__3890),
            .I(\uart.timer_CountZ0Z_7 ));
    LocalMux I__776 (
            .O(N__3885),
            .I(\uart.timer_CountZ0Z_7 ));
    LocalMux I__775 (
            .O(N__3882),
            .I(\uart.timer_CountZ0Z_7 ));
    LocalMux I__774 (
            .O(N__3875),
            .I(\uart.timer_CountZ0Z_7 ));
    InMux I__773 (
            .O(N__3860),
            .I(N__3857));
    LocalMux I__772 (
            .O(N__3857),
            .I(N__3854));
    Span4Mux_h I__771 (
            .O(N__3854),
            .I(N__3849));
    InMux I__770 (
            .O(N__3853),
            .I(N__3846));
    InMux I__769 (
            .O(N__3852),
            .I(N__3843));
    Odrv4 I__768 (
            .O(N__3849),
            .I(\uart.N_41 ));
    LocalMux I__767 (
            .O(N__3846),
            .I(\uart.N_41 ));
    LocalMux I__766 (
            .O(N__3843),
            .I(\uart.N_41 ));
    InMux I__765 (
            .O(N__3836),
            .I(N__3833));
    LocalMux I__764 (
            .O(N__3833),
            .I(N__3830));
    Span4Mux_h I__763 (
            .O(N__3830),
            .I(N__3824));
    InMux I__762 (
            .O(N__3829),
            .I(N__3821));
    InMux I__761 (
            .O(N__3828),
            .I(N__3816));
    InMux I__760 (
            .O(N__3827),
            .I(N__3816));
    Odrv4 I__759 (
            .O(N__3824),
            .I(\uart.state_srsts_0_o4_0_a2_0_4 ));
    LocalMux I__758 (
            .O(N__3821),
            .I(\uart.state_srsts_0_o4_0_a2_0_4 ));
    LocalMux I__757 (
            .O(N__3816),
            .I(\uart.state_srsts_0_o4_0_a2_0_4 ));
    CEMux I__756 (
            .O(N__3809),
            .I(N__3806));
    LocalMux I__755 (
            .O(N__3806),
            .I(N__3803));
    Odrv4 I__754 (
            .O(N__3803),
            .I(\uart_frame_decoder.uart_data_rdy_c_0 ));
    InMux I__753 (
            .O(N__3800),
            .I(N__3792));
    InMux I__752 (
            .O(N__3799),
            .I(N__3792));
    InMux I__751 (
            .O(N__3798),
            .I(N__3789));
    InMux I__750 (
            .O(N__3797),
            .I(N__3786));
    LocalMux I__749 (
            .O(N__3792),
            .I(N__3783));
    LocalMux I__748 (
            .O(N__3789),
            .I(\uart_frame_decoder.state_1Z0Z_3 ));
    LocalMux I__747 (
            .O(N__3786),
            .I(\uart_frame_decoder.state_1Z0Z_3 ));
    Odrv12 I__746 (
            .O(N__3783),
            .I(\uart_frame_decoder.state_1Z0Z_3 ));
    InMux I__745 (
            .O(N__3776),
            .I(N__3770));
    InMux I__744 (
            .O(N__3775),
            .I(N__3763));
    InMux I__743 (
            .O(N__3774),
            .I(N__3763));
    InMux I__742 (
            .O(N__3773),
            .I(N__3763));
    LocalMux I__741 (
            .O(N__3770),
            .I(N__3759));
    LocalMux I__740 (
            .O(N__3763),
            .I(N__3756));
    InMux I__739 (
            .O(N__3762),
            .I(N__3753));
    Span4Mux_s1_v I__738 (
            .O(N__3759),
            .I(N__3748));
    Span4Mux_s1_v I__737 (
            .O(N__3756),
            .I(N__3748));
    LocalMux I__736 (
            .O(N__3753),
            .I(\uart_frame_decoder.state_1Z0Z_6 ));
    Odrv4 I__735 (
            .O(N__3748),
            .I(\uart_frame_decoder.state_1Z0Z_6 ));
    InMux I__734 (
            .O(N__3743),
            .I(N__3739));
    InMux I__733 (
            .O(N__3742),
            .I(N__3736));
    LocalMux I__732 (
            .O(N__3739),
            .I(N__3729));
    LocalMux I__731 (
            .O(N__3736),
            .I(N__3729));
    InMux I__730 (
            .O(N__3735),
            .I(N__3724));
    InMux I__729 (
            .O(N__3734),
            .I(N__3724));
    Odrv12 I__728 (
            .O(N__3729),
            .I(\uart_frame_decoder.state_1Z0Z_2 ));
    LocalMux I__727 (
            .O(N__3724),
            .I(\uart_frame_decoder.state_1Z0Z_2 ));
    IoInMux I__726 (
            .O(N__3719),
            .I(N__3716));
    LocalMux I__725 (
            .O(N__3716),
            .I(N__3713));
    IoSpan4Mux I__724 (
            .O(N__3713),
            .I(N__3710));
    Odrv4 I__723 (
            .O(N__3710),
            .I(uart_frame_decoder_N_130_i));
    CascadeMux I__722 (
            .O(N__3707),
            .I(\reset_module_System.reset6_14_cascade_ ));
    InMux I__721 (
            .O(N__3704),
            .I(N__3691));
    InMux I__720 (
            .O(N__3703),
            .I(N__3691));
    InMux I__719 (
            .O(N__3702),
            .I(N__3691));
    InMux I__718 (
            .O(N__3701),
            .I(N__3691));
    InMux I__717 (
            .O(N__3700),
            .I(N__3688));
    LocalMux I__716 (
            .O(N__3691),
            .I(\reset_module_System.reset6_19 ));
    LocalMux I__715 (
            .O(N__3688),
            .I(\reset_module_System.reset6_19 ));
    CascadeMux I__714 (
            .O(N__3683),
            .I(N__3679));
    CascadeMux I__713 (
            .O(N__3682),
            .I(N__3675));
    InMux I__712 (
            .O(N__3679),
            .I(N__3668));
    InMux I__711 (
            .O(N__3678),
            .I(N__3668));
    InMux I__710 (
            .O(N__3675),
            .I(N__3668));
    LocalMux I__709 (
            .O(N__3668),
            .I(N__3663));
    InMux I__708 (
            .O(N__3667),
            .I(N__3658));
    InMux I__707 (
            .O(N__3666),
            .I(N__3658));
    Odrv4 I__706 (
            .O(N__3663),
            .I(\reset_module_System.reset6_14 ));
    LocalMux I__705 (
            .O(N__3658),
            .I(\reset_module_System.reset6_14 ));
    InMux I__704 (
            .O(N__3653),
            .I(N__3650));
    LocalMux I__703 (
            .O(N__3650),
            .I(\reset_module_System.reset6_19_1 ));
    InMux I__702 (
            .O(N__3647),
            .I(N__3644));
    LocalMux I__701 (
            .O(N__3644),
            .I(\reset_module_System.reset6_13 ));
    InMux I__700 (
            .O(N__3641),
            .I(N__3635));
    InMux I__699 (
            .O(N__3640),
            .I(N__3632));
    InMux I__698 (
            .O(N__3639),
            .I(N__3629));
    InMux I__697 (
            .O(N__3638),
            .I(N__3626));
    LocalMux I__696 (
            .O(N__3635),
            .I(N__3621));
    LocalMux I__695 (
            .O(N__3632),
            .I(N__3616));
    LocalMux I__694 (
            .O(N__3629),
            .I(N__3616));
    LocalMux I__693 (
            .O(N__3626),
            .I(N__3612));
    CascadeMux I__692 (
            .O(N__3625),
            .I(N__3608));
    CascadeMux I__691 (
            .O(N__3624),
            .I(N__3603));
    Span4Mux_h I__690 (
            .O(N__3621),
            .I(N__3595));
    Span4Mux_h I__689 (
            .O(N__3616),
            .I(N__3595));
    InMux I__688 (
            .O(N__3615),
            .I(N__3592));
    Span4Mux_h I__687 (
            .O(N__3612),
            .I(N__3589));
    InMux I__686 (
            .O(N__3611),
            .I(N__3578));
    InMux I__685 (
            .O(N__3608),
            .I(N__3578));
    InMux I__684 (
            .O(N__3607),
            .I(N__3578));
    InMux I__683 (
            .O(N__3606),
            .I(N__3578));
    InMux I__682 (
            .O(N__3603),
            .I(N__3578));
    InMux I__681 (
            .O(N__3602),
            .I(N__3571));
    InMux I__680 (
            .O(N__3601),
            .I(N__3571));
    InMux I__679 (
            .O(N__3600),
            .I(N__3571));
    Odrv4 I__678 (
            .O(N__3595),
            .I(\uart.stateZ0Z_3 ));
    LocalMux I__677 (
            .O(N__3592),
            .I(\uart.stateZ0Z_3 ));
    Odrv4 I__676 (
            .O(N__3589),
            .I(\uart.stateZ0Z_3 ));
    LocalMux I__675 (
            .O(N__3578),
            .I(\uart.stateZ0Z_3 ));
    LocalMux I__674 (
            .O(N__3571),
            .I(\uart.stateZ0Z_3 ));
    CascadeMux I__673 (
            .O(N__3560),
            .I(N__3557));
    InMux I__672 (
            .O(N__3557),
            .I(N__3554));
    LocalMux I__671 (
            .O(N__3554),
            .I(\uart.g3_0_0 ));
    InMux I__670 (
            .O(N__3551),
            .I(N__3546));
    InMux I__669 (
            .O(N__3550),
            .I(N__3543));
    CascadeMux I__668 (
            .O(N__3549),
            .I(N__3540));
    LocalMux I__667 (
            .O(N__3546),
            .I(N__3536));
    LocalMux I__666 (
            .O(N__3543),
            .I(N__3533));
    InMux I__665 (
            .O(N__3540),
            .I(N__3527));
    InMux I__664 (
            .O(N__3539),
            .I(N__3524));
    Span4Mux_v I__663 (
            .O(N__3536),
            .I(N__3519));
    Span4Mux_v I__662 (
            .O(N__3533),
            .I(N__3519));
    InMux I__661 (
            .O(N__3532),
            .I(N__3512));
    InMux I__660 (
            .O(N__3531),
            .I(N__3512));
    InMux I__659 (
            .O(N__3530),
            .I(N__3512));
    LocalMux I__658 (
            .O(N__3527),
            .I(N__3509));
    LocalMux I__657 (
            .O(N__3524),
            .I(N__3506));
    Odrv4 I__656 (
            .O(N__3519),
            .I(\uart.timer_CountZ0Z_4 ));
    LocalMux I__655 (
            .O(N__3512),
            .I(\uart.timer_CountZ0Z_4 ));
    Odrv4 I__654 (
            .O(N__3509),
            .I(\uart.timer_CountZ0Z_4 ));
    Odrv4 I__653 (
            .O(N__3506),
            .I(\uart.timer_CountZ0Z_4 ));
    InMux I__652 (
            .O(N__3497),
            .I(N__3494));
    LocalMux I__651 (
            .O(N__3494),
            .I(N__3491));
    Span4Mux_h I__650 (
            .O(N__3491),
            .I(N__3488));
    Odrv4 I__649 (
            .O(N__3488),
            .I(\uart.state_0_sqmuxa_1_d_0 ));
    CascadeMux I__648 (
            .O(N__3485),
            .I(N__3482));
    InMux I__647 (
            .O(N__3482),
            .I(N__3479));
    LocalMux I__646 (
            .O(N__3479),
            .I(N__3474));
    InMux I__645 (
            .O(N__3478),
            .I(N__3467));
    InMux I__644 (
            .O(N__3477),
            .I(N__3467));
    Span4Mux_h I__643 (
            .O(N__3474),
            .I(N__3464));
    InMux I__642 (
            .O(N__3473),
            .I(N__3459));
    InMux I__641 (
            .O(N__3472),
            .I(N__3459));
    LocalMux I__640 (
            .O(N__3467),
            .I(\uart.timer_CountZ0Z_1 ));
    Odrv4 I__639 (
            .O(N__3464),
            .I(\uart.timer_CountZ0Z_1 ));
    LocalMux I__638 (
            .O(N__3459),
            .I(\uart.timer_CountZ0Z_1 ));
    InMux I__637 (
            .O(N__3452),
            .I(N__3449));
    LocalMux I__636 (
            .O(N__3449),
            .I(\uart.g1_3 ));
    InMux I__635 (
            .O(N__3446),
            .I(N__3443));
    LocalMux I__634 (
            .O(N__3443),
            .I(N__3438));
    InMux I__633 (
            .O(N__3442),
            .I(N__3433));
    InMux I__632 (
            .O(N__3441),
            .I(N__3433));
    Odrv4 I__631 (
            .O(N__3438),
            .I(\uart.stateZ0Z_2 ));
    LocalMux I__630 (
            .O(N__3433),
            .I(\uart.stateZ0Z_2 ));
    InMux I__629 (
            .O(N__3428),
            .I(N__3424));
    InMux I__628 (
            .O(N__3427),
            .I(N__3421));
    LocalMux I__627 (
            .O(N__3424),
            .I(N__3418));
    LocalMux I__626 (
            .O(N__3421),
            .I(N__3415));
    Span4Mux_s3_v I__625 (
            .O(N__3418),
            .I(N__3410));
    Span4Mux_v I__624 (
            .O(N__3415),
            .I(N__3410));
    Odrv4 I__623 (
            .O(N__3410),
            .I(\uart.un1_state_5 ));
    InMux I__622 (
            .O(N__3407),
            .I(N__3404));
    LocalMux I__621 (
            .O(N__3404),
            .I(N__3401));
    Span4Mux_v I__620 (
            .O(N__3401),
            .I(N__3397));
    InMux I__619 (
            .O(N__3400),
            .I(N__3394));
    Span4Mux_h I__618 (
            .O(N__3397),
            .I(N__3391));
    LocalMux I__617 (
            .O(N__3394),
            .I(\uart.N_177 ));
    Odrv4 I__616 (
            .O(N__3391),
            .I(\uart.N_177 ));
    CascadeMux I__615 (
            .O(N__3386),
            .I(N__3382));
    InMux I__614 (
            .O(N__3385),
            .I(N__3376));
    InMux I__613 (
            .O(N__3382),
            .I(N__3373));
    InMux I__612 (
            .O(N__3381),
            .I(N__3368));
    InMux I__611 (
            .O(N__3380),
            .I(N__3368));
    InMux I__610 (
            .O(N__3379),
            .I(N__3365));
    LocalMux I__609 (
            .O(N__3376),
            .I(N__3357));
    LocalMux I__608 (
            .O(N__3373),
            .I(N__3357));
    LocalMux I__607 (
            .O(N__3368),
            .I(N__3352));
    LocalMux I__606 (
            .O(N__3365),
            .I(N__3352));
    InMux I__605 (
            .O(N__3364),
            .I(N__3345));
    InMux I__604 (
            .O(N__3363),
            .I(N__3345));
    InMux I__603 (
            .O(N__3362),
            .I(N__3340));
    Span4Mux_v I__602 (
            .O(N__3357),
            .I(N__3335));
    Span4Mux_s1_v I__601 (
            .O(N__3352),
            .I(N__3335));
    InMux I__600 (
            .O(N__3351),
            .I(N__3330));
    InMux I__599 (
            .O(N__3350),
            .I(N__3330));
    LocalMux I__598 (
            .O(N__3345),
            .I(N__3327));
    InMux I__597 (
            .O(N__3344),
            .I(N__3322));
    InMux I__596 (
            .O(N__3343),
            .I(N__3322));
    LocalMux I__595 (
            .O(N__3340),
            .I(reset_system));
    Odrv4 I__594 (
            .O(N__3335),
            .I(reset_system));
    LocalMux I__593 (
            .O(N__3330),
            .I(reset_system));
    Odrv12 I__592 (
            .O(N__3327),
            .I(reset_system));
    LocalMux I__591 (
            .O(N__3322),
            .I(reset_system));
    InMux I__590 (
            .O(N__3311),
            .I(N__3308));
    LocalMux I__589 (
            .O(N__3308),
            .I(\uart.N_28_mux ));
    CascadeMux I__588 (
            .O(N__3305),
            .I(\uart.N_8_cascade_ ));
    InMux I__587 (
            .O(N__3302),
            .I(N__3297));
    InMux I__586 (
            .O(N__3301),
            .I(N__3294));
    InMux I__585 (
            .O(N__3300),
            .I(N__3291));
    LocalMux I__584 (
            .O(N__3297),
            .I(N__3286));
    LocalMux I__583 (
            .O(N__3294),
            .I(N__3286));
    LocalMux I__582 (
            .O(N__3291),
            .I(N__3281));
    Span4Mux_h I__581 (
            .O(N__3286),
            .I(N__3281));
    Odrv4 I__580 (
            .O(N__3281),
            .I(\uart_frame_decoder.state_1Z0Z_4 ));
    CascadeMux I__579 (
            .O(N__3278),
            .I(N__3272));
    InMux I__578 (
            .O(N__3277),
            .I(N__3269));
    InMux I__577 (
            .O(N__3276),
            .I(N__3266));
    InMux I__576 (
            .O(N__3275),
            .I(N__3261));
    InMux I__575 (
            .O(N__3272),
            .I(N__3261));
    LocalMux I__574 (
            .O(N__3269),
            .I(N__3258));
    LocalMux I__573 (
            .O(N__3266),
            .I(N__3255));
    LocalMux I__572 (
            .O(N__3261),
            .I(N__3252));
    Odrv12 I__571 (
            .O(N__3258),
            .I(\uart_frame_decoder.state_1Z0Z_5 ));
    Odrv4 I__570 (
            .O(N__3255),
            .I(\uart_frame_decoder.state_1Z0Z_5 ));
    Odrv4 I__569 (
            .O(N__3252),
            .I(\uart_frame_decoder.state_1Z0Z_5 ));
    InMux I__568 (
            .O(N__3245),
            .I(N__3242));
    LocalMux I__567 (
            .O(N__3242),
            .I(\reset_module_System.reset6_3 ));
    InMux I__566 (
            .O(N__3239),
            .I(N__3236));
    LocalMux I__565 (
            .O(N__3236),
            .I(\uart.timer_Count_RNI3B101Z0Z_6 ));
    CascadeMux I__564 (
            .O(N__3233),
            .I(N__3228));
    InMux I__563 (
            .O(N__3232),
            .I(N__3221));
    InMux I__562 (
            .O(N__3231),
            .I(N__3221));
    InMux I__561 (
            .O(N__3228),
            .I(N__3221));
    LocalMux I__560 (
            .O(N__3221),
            .I(N__3218));
    Odrv4 I__559 (
            .O(N__3218),
            .I(\uart.un4_timer_Count_1_c5 ));
    InMux I__558 (
            .O(N__3215),
            .I(N__3212));
    LocalMux I__557 (
            .O(N__3212),
            .I(N__3209));
    Odrv4 I__556 (
            .O(N__3209),
            .I(\uart.un1_state_2_0_a3_2 ));
    CascadeMux I__555 (
            .O(N__3206),
            .I(N__3203));
    InMux I__554 (
            .O(N__3203),
            .I(N__3196));
    InMux I__553 (
            .O(N__3202),
            .I(N__3196));
    CascadeMux I__552 (
            .O(N__3201),
            .I(N__3192));
    LocalMux I__551 (
            .O(N__3196),
            .I(N__3189));
    InMux I__550 (
            .O(N__3195),
            .I(N__3184));
    InMux I__549 (
            .O(N__3192),
            .I(N__3184));
    Odrv4 I__548 (
            .O(N__3189),
            .I(\uart.timer_CountZ0Z_0 ));
    LocalMux I__547 (
            .O(N__3184),
            .I(\uart.timer_CountZ0Z_0 ));
    InMux I__546 (
            .O(N__3179),
            .I(N__3176));
    LocalMux I__545 (
            .O(N__3176),
            .I(\uart.timer_Count_RNI22NA1Z0Z_4 ));
    CascadeMux I__544 (
            .O(N__3173),
            .I(N__3168));
    CascadeMux I__543 (
            .O(N__3172),
            .I(N__3165));
    InMux I__542 (
            .O(N__3171),
            .I(N__3162));
    InMux I__541 (
            .O(N__3168),
            .I(N__3153));
    InMux I__540 (
            .O(N__3165),
            .I(N__3153));
    LocalMux I__539 (
            .O(N__3162),
            .I(N__3150));
    CascadeMux I__538 (
            .O(N__3161),
            .I(N__3143));
    CascadeMux I__537 (
            .O(N__3160),
            .I(N__3140));
    CascadeMux I__536 (
            .O(N__3159),
            .I(N__3136));
    InMux I__535 (
            .O(N__3158),
            .I(N__3132));
    LocalMux I__534 (
            .O(N__3153),
            .I(N__3129));
    Span4Mux_h I__533 (
            .O(N__3150),
            .I(N__3126));
    InMux I__532 (
            .O(N__3149),
            .I(N__3123));
    InMux I__531 (
            .O(N__3148),
            .I(N__3120));
    InMux I__530 (
            .O(N__3147),
            .I(N__3115));
    InMux I__529 (
            .O(N__3146),
            .I(N__3115));
    InMux I__528 (
            .O(N__3143),
            .I(N__3106));
    InMux I__527 (
            .O(N__3140),
            .I(N__3106));
    InMux I__526 (
            .O(N__3139),
            .I(N__3106));
    InMux I__525 (
            .O(N__3136),
            .I(N__3106));
    InMux I__524 (
            .O(N__3135),
            .I(N__3103));
    LocalMux I__523 (
            .O(N__3132),
            .I(N__3098));
    Span4Mux_h I__522 (
            .O(N__3129),
            .I(N__3098));
    Odrv4 I__521 (
            .O(N__3126),
            .I(\uart.bit_CountZ0Z_0 ));
    LocalMux I__520 (
            .O(N__3123),
            .I(\uart.bit_CountZ0Z_0 ));
    LocalMux I__519 (
            .O(N__3120),
            .I(\uart.bit_CountZ0Z_0 ));
    LocalMux I__518 (
            .O(N__3115),
            .I(\uart.bit_CountZ0Z_0 ));
    LocalMux I__517 (
            .O(N__3106),
            .I(\uart.bit_CountZ0Z_0 ));
    LocalMux I__516 (
            .O(N__3103),
            .I(\uart.bit_CountZ0Z_0 ));
    Odrv4 I__515 (
            .O(N__3098),
            .I(\uart.bit_CountZ0Z_0 ));
    CascadeMux I__514 (
            .O(N__3083),
            .I(N__3080));
    InMux I__513 (
            .O(N__3080),
            .I(N__3077));
    LocalMux I__512 (
            .O(N__3077),
            .I(N__3070));
    InMux I__511 (
            .O(N__3076),
            .I(N__3067));
    InMux I__510 (
            .O(N__3075),
            .I(N__3062));
    InMux I__509 (
            .O(N__3074),
            .I(N__3062));
    InMux I__508 (
            .O(N__3073),
            .I(N__3056));
    Span4Mux_v I__507 (
            .O(N__3070),
            .I(N__3053));
    LocalMux I__506 (
            .O(N__3067),
            .I(N__3048));
    LocalMux I__505 (
            .O(N__3062),
            .I(N__3048));
    InMux I__504 (
            .O(N__3061),
            .I(N__3045));
    InMux I__503 (
            .O(N__3060),
            .I(N__3040));
    InMux I__502 (
            .O(N__3059),
            .I(N__3040));
    LocalMux I__501 (
            .O(N__3056),
            .I(\uart.bit_CountZ0Z_2 ));
    Odrv4 I__500 (
            .O(N__3053),
            .I(\uart.bit_CountZ0Z_2 ));
    Odrv4 I__499 (
            .O(N__3048),
            .I(\uart.bit_CountZ0Z_2 ));
    LocalMux I__498 (
            .O(N__3045),
            .I(\uart.bit_CountZ0Z_2 ));
    LocalMux I__497 (
            .O(N__3040),
            .I(\uart.bit_CountZ0Z_2 ));
    InMux I__496 (
            .O(N__3029),
            .I(N__3026));
    LocalMux I__495 (
            .O(N__3026),
            .I(N__3020));
    InMux I__494 (
            .O(N__3025),
            .I(N__3017));
    InMux I__493 (
            .O(N__3024),
            .I(N__3012));
    InMux I__492 (
            .O(N__3023),
            .I(N__3012));
    Span4Mux_h I__491 (
            .O(N__3020),
            .I(N__3004));
    LocalMux I__490 (
            .O(N__3017),
            .I(N__2999));
    LocalMux I__489 (
            .O(N__3012),
            .I(N__2999));
    InMux I__488 (
            .O(N__3011),
            .I(N__2994));
    InMux I__487 (
            .O(N__3010),
            .I(N__2994));
    InMux I__486 (
            .O(N__3009),
            .I(N__2987));
    InMux I__485 (
            .O(N__3008),
            .I(N__2987));
    InMux I__484 (
            .O(N__3007),
            .I(N__2987));
    Odrv4 I__483 (
            .O(N__3004),
            .I(\uart.bit_CountZ0Z_1 ));
    Odrv4 I__482 (
            .O(N__2999),
            .I(\uart.bit_CountZ0Z_1 ));
    LocalMux I__481 (
            .O(N__2994),
            .I(\uart.bit_CountZ0Z_1 ));
    LocalMux I__480 (
            .O(N__2987),
            .I(\uart.bit_CountZ0Z_1 ));
    CascadeMux I__479 (
            .O(N__2978),
            .I(\uart.g1_4_cascade_ ));
    InMux I__478 (
            .O(N__2975),
            .I(N__2972));
    LocalMux I__477 (
            .O(N__2972),
            .I(N__2969));
    Span4Mux_v I__476 (
            .O(N__2969),
            .I(N__2966));
    Odrv4 I__475 (
            .O(N__2966),
            .I(\uart.g1_0 ));
    CascadeMux I__474 (
            .O(N__2963),
            .I(N__2958));
    InMux I__473 (
            .O(N__2962),
            .I(N__2954));
    InMux I__472 (
            .O(N__2961),
            .I(N__2947));
    InMux I__471 (
            .O(N__2958),
            .I(N__2947));
    InMux I__470 (
            .O(N__2957),
            .I(N__2947));
    LocalMux I__469 (
            .O(N__2954),
            .I(\uart.timer_Count_fastZ0Z_2 ));
    LocalMux I__468 (
            .O(N__2947),
            .I(\uart.timer_Count_fastZ0Z_2 ));
    CascadeMux I__467 (
            .O(N__2942),
            .I(\reset_module_System.reset6_11_cascade_ ));
    CascadeMux I__466 (
            .O(N__2939),
            .I(\reset_module_System.reset6_19_cascade_ ));
    InMux I__465 (
            .O(N__2936),
            .I(N__2933));
    LocalMux I__464 (
            .O(N__2933),
            .I(\uart.N_66 ));
    InMux I__463 (
            .O(N__2930),
            .I(N__2927));
    LocalMux I__462 (
            .O(N__2927),
            .I(\uart.N_51 ));
    InMux I__461 (
            .O(N__2924),
            .I(N__2919));
    CascadeMux I__460 (
            .O(N__2923),
            .I(N__2914));
    InMux I__459 (
            .O(N__2922),
            .I(N__2911));
    LocalMux I__458 (
            .O(N__2919),
            .I(N__2908));
    InMux I__457 (
            .O(N__2918),
            .I(N__2901));
    InMux I__456 (
            .O(N__2917),
            .I(N__2901));
    InMux I__455 (
            .O(N__2914),
            .I(N__2901));
    LocalMux I__454 (
            .O(N__2911),
            .I(\uart.timer_Count_fastZ0Z_3 ));
    Odrv4 I__453 (
            .O(N__2908),
            .I(\uart.timer_Count_fastZ0Z_3 ));
    LocalMux I__452 (
            .O(N__2901),
            .I(\uart.timer_Count_fastZ0Z_3 ));
    InMux I__451 (
            .O(N__2894),
            .I(N__2891));
    LocalMux I__450 (
            .O(N__2891),
            .I(N__2888));
    Odrv12 I__449 (
            .O(N__2888),
            .I(\uart.N_5 ));
    CascadeMux I__448 (
            .O(N__2885),
            .I(N__2880));
    CascadeMux I__447 (
            .O(N__2884),
            .I(N__2877));
    InMux I__446 (
            .O(N__2883),
            .I(N__2874));
    InMux I__445 (
            .O(N__2880),
            .I(N__2871));
    InMux I__444 (
            .O(N__2877),
            .I(N__2868));
    LocalMux I__443 (
            .O(N__2874),
            .I(N__2863));
    LocalMux I__442 (
            .O(N__2871),
            .I(N__2863));
    LocalMux I__441 (
            .O(N__2868),
            .I(\uart.stateZ0Z_1 ));
    Odrv4 I__440 (
            .O(N__2863),
            .I(\uart.stateZ0Z_1 ));
    InMux I__439 (
            .O(N__2858),
            .I(N__2855));
    LocalMux I__438 (
            .O(N__2855),
            .I(\uart.N_151 ));
    CascadeMux I__437 (
            .O(N__2852),
            .I(N__2849));
    InMux I__436 (
            .O(N__2849),
            .I(N__2842));
    InMux I__435 (
            .O(N__2848),
            .I(N__2842));
    InMux I__434 (
            .O(N__2847),
            .I(N__2838));
    LocalMux I__433 (
            .O(N__2842),
            .I(N__2831));
    InMux I__432 (
            .O(N__2841),
            .I(N__2828));
    LocalMux I__431 (
            .O(N__2838),
            .I(N__2825));
    InMux I__430 (
            .O(N__2837),
            .I(N__2816));
    InMux I__429 (
            .O(N__2836),
            .I(N__2816));
    InMux I__428 (
            .O(N__2835),
            .I(N__2816));
    InMux I__427 (
            .O(N__2834),
            .I(N__2816));
    Odrv4 I__426 (
            .O(N__2831),
            .I(\uart.N_174 ));
    LocalMux I__425 (
            .O(N__2828),
            .I(\uart.N_174 ));
    Odrv4 I__424 (
            .O(N__2825),
            .I(\uart.N_174 ));
    LocalMux I__423 (
            .O(N__2816),
            .I(\uart.N_174 ));
    InMux I__422 (
            .O(N__2807),
            .I(N__2804));
    LocalMux I__421 (
            .O(N__2804),
            .I(\uart.state_srsts_0_a3_2_0_4 ));
    InMux I__420 (
            .O(N__2801),
            .I(N__2798));
    LocalMux I__419 (
            .O(N__2798),
            .I(N__2794));
    InMux I__418 (
            .O(N__2797),
            .I(N__2791));
    Odrv4 I__417 (
            .O(N__2794),
            .I(\uart.state_1_sqmuxa ));
    LocalMux I__416 (
            .O(N__2791),
            .I(\uart.state_1_sqmuxa ));
    InMux I__415 (
            .O(N__2786),
            .I(N__2783));
    LocalMux I__414 (
            .O(N__2783),
            .I(N__2780));
    Odrv4 I__413 (
            .O(N__2780),
            .I(\uart.data_AuxZ0Z_3 ));
    CEMux I__412 (
            .O(N__2777),
            .I(N__2774));
    LocalMux I__411 (
            .O(N__2774),
            .I(N__2771));
    Odrv12 I__410 (
            .O(N__2771),
            .I(\uart.N_117_0 ));
    InMux I__409 (
            .O(N__2768),
            .I(N__2765));
    LocalMux I__408 (
            .O(N__2765),
            .I(N__2762));
    Span4Mux_h I__407 (
            .O(N__2762),
            .I(N__2759));
    Odrv4 I__406 (
            .O(N__2759),
            .I(\uart.data_AuxZ0Z_4 ));
    CEMux I__405 (
            .O(N__2756),
            .I(N__2753));
    LocalMux I__404 (
            .O(N__2753),
            .I(N__2750));
    Span4Mux_h I__403 (
            .O(N__2750),
            .I(N__2747));
    Odrv4 I__402 (
            .O(N__2747),
            .I(\uart.N_116_0 ));
    SRMux I__401 (
            .O(N__2744),
            .I(N__2736));
    SRMux I__400 (
            .O(N__2743),
            .I(N__2733));
    SRMux I__399 (
            .O(N__2742),
            .I(N__2730));
    SRMux I__398 (
            .O(N__2741),
            .I(N__2723));
    SRMux I__397 (
            .O(N__2740),
            .I(N__2720));
    SRMux I__396 (
            .O(N__2739),
            .I(N__2717));
    LocalMux I__395 (
            .O(N__2736),
            .I(N__2713));
    LocalMux I__394 (
            .O(N__2733),
            .I(N__2708));
    LocalMux I__393 (
            .O(N__2730),
            .I(N__2708));
    SRMux I__392 (
            .O(N__2729),
            .I(N__2705));
    InMux I__391 (
            .O(N__2728),
            .I(N__2697));
    InMux I__390 (
            .O(N__2727),
            .I(N__2697));
    InMux I__389 (
            .O(N__2726),
            .I(N__2697));
    LocalMux I__388 (
            .O(N__2723),
            .I(N__2689));
    LocalMux I__387 (
            .O(N__2720),
            .I(N__2689));
    LocalMux I__386 (
            .O(N__2717),
            .I(N__2686));
    InMux I__385 (
            .O(N__2716),
            .I(N__2683));
    Span4Mux_h I__384 (
            .O(N__2713),
            .I(N__2679));
    Span4Mux_v I__383 (
            .O(N__2708),
            .I(N__2676));
    LocalMux I__382 (
            .O(N__2705),
            .I(N__2673));
    SRMux I__381 (
            .O(N__2704),
            .I(N__2670));
    LocalMux I__380 (
            .O(N__2697),
            .I(N__2667));
    InMux I__379 (
            .O(N__2696),
            .I(N__2660));
    InMux I__378 (
            .O(N__2695),
            .I(N__2660));
    InMux I__377 (
            .O(N__2694),
            .I(N__2660));
    Span4Mux_v I__376 (
            .O(N__2689),
            .I(N__2653));
    Span4Mux_s2_v I__375 (
            .O(N__2686),
            .I(N__2653));
    LocalMux I__374 (
            .O(N__2683),
            .I(N__2653));
    InMux I__373 (
            .O(N__2682),
            .I(N__2650));
    Odrv4 I__372 (
            .O(N__2679),
            .I(\uart.state_RNIAFHLZ0Z_4 ));
    Odrv4 I__371 (
            .O(N__2676),
            .I(\uart.state_RNIAFHLZ0Z_4 ));
    Odrv12 I__370 (
            .O(N__2673),
            .I(\uart.state_RNIAFHLZ0Z_4 ));
    LocalMux I__369 (
            .O(N__2670),
            .I(\uart.state_RNIAFHLZ0Z_4 ));
    Odrv4 I__368 (
            .O(N__2667),
            .I(\uart.state_RNIAFHLZ0Z_4 ));
    LocalMux I__367 (
            .O(N__2660),
            .I(\uart.state_RNIAFHLZ0Z_4 ));
    Odrv4 I__366 (
            .O(N__2653),
            .I(\uart.state_RNIAFHLZ0Z_4 ));
    LocalMux I__365 (
            .O(N__2650),
            .I(\uart.state_RNIAFHLZ0Z_4 ));
    CascadeMux I__364 (
            .O(N__2633),
            .I(N__2629));
    CascadeMux I__363 (
            .O(N__2632),
            .I(N__2623));
    InMux I__362 (
            .O(N__2629),
            .I(N__2615));
    InMux I__361 (
            .O(N__2628),
            .I(N__2615));
    InMux I__360 (
            .O(N__2627),
            .I(N__2602));
    InMux I__359 (
            .O(N__2626),
            .I(N__2602));
    InMux I__358 (
            .O(N__2623),
            .I(N__2602));
    InMux I__357 (
            .O(N__2622),
            .I(N__2602));
    InMux I__356 (
            .O(N__2621),
            .I(N__2602));
    InMux I__355 (
            .O(N__2620),
            .I(N__2602));
    LocalMux I__354 (
            .O(N__2615),
            .I(\uart.timer_CountZ0Z_2 ));
    LocalMux I__353 (
            .O(N__2602),
            .I(\uart.timer_CountZ0Z_2 ));
    CascadeMux I__352 (
            .O(N__2597),
            .I(\uart.state_srsts_0_a3_1_4_cascade_ ));
    InMux I__351 (
            .O(N__2594),
            .I(N__2590));
    InMux I__350 (
            .O(N__2593),
            .I(N__2587));
    LocalMux I__349 (
            .O(N__2590),
            .I(\uart.timer_Count_fastZ0Z_4 ));
    LocalMux I__348 (
            .O(N__2587),
            .I(\uart.timer_Count_fastZ0Z_4 ));
    CascadeMux I__347 (
            .O(N__2582),
            .I(N__2579));
    InMux I__346 (
            .O(N__2579),
            .I(N__2576));
    LocalMux I__345 (
            .O(N__2576),
            .I(N__2573));
    Span4Mux_v I__344 (
            .O(N__2573),
            .I(N__2570));
    Odrv4 I__343 (
            .O(N__2570),
            .I(\uart.timer_Count10lto4_0 ));
    CascadeMux I__342 (
            .O(N__2567),
            .I(\uart.timer_Count10lto4_0_cascade_ ));
    CascadeMux I__341 (
            .O(N__2564),
            .I(\uart.N_51_cascade_ ));
    CascadeMux I__340 (
            .O(N__2561),
            .I(N__2558));
    InMux I__339 (
            .O(N__2558),
            .I(N__2554));
    InMux I__338 (
            .O(N__2557),
            .I(N__2551));
    LocalMux I__337 (
            .O(N__2554),
            .I(\uart.N_146_0 ));
    LocalMux I__336 (
            .O(N__2551),
            .I(\uart.N_146_0 ));
    CascadeMux I__335 (
            .O(N__2546),
            .I(\uart.data_14_1_cascade_ ));
    SRMux I__334 (
            .O(N__2543),
            .I(N__2540));
    LocalMux I__333 (
            .O(N__2540),
            .I(N__2537));
    Span4Mux_s2_v I__332 (
            .O(N__2537),
            .I(N__2534));
    Odrv4 I__331 (
            .O(N__2534),
            .I(\uart.state_RNILS533Z0Z_4 ));
    CascadeMux I__330 (
            .O(N__2531),
            .I(\uart.state_RNILS533Z0Z_4_cascade_ ));
    CEMux I__329 (
            .O(N__2528),
            .I(N__2525));
    LocalMux I__328 (
            .O(N__2525),
            .I(\uart.state_1_sqmuxa_0 ));
    CascadeMux I__327 (
            .O(N__2522),
            .I(\uart.un4_timer_Count_1_c2_cascade_ ));
    InMux I__326 (
            .O(N__2519),
            .I(N__2513));
    InMux I__325 (
            .O(N__2518),
            .I(N__2513));
    LocalMux I__324 (
            .O(N__2513),
            .I(\uart.data_Auxce_0_4 ));
    CEMux I__323 (
            .O(N__2510),
            .I(N__2507));
    LocalMux I__322 (
            .O(N__2507),
            .I(N__2504));
    Odrv4 I__321 (
            .O(N__2504),
            .I(\uart.N_113_0 ));
    InMux I__320 (
            .O(N__2501),
            .I(N__2498));
    LocalMux I__319 (
            .O(N__2498),
            .I(N__2494));
    InMux I__318 (
            .O(N__2497),
            .I(N__2491));
    Odrv4 I__317 (
            .O(N__2494),
            .I(\uart.N_133_0 ));
    LocalMux I__316 (
            .O(N__2491),
            .I(\uart.N_133_0 ));
    InMux I__315 (
            .O(N__2486),
            .I(N__2480));
    InMux I__314 (
            .O(N__2485),
            .I(N__2480));
    LocalMux I__313 (
            .O(N__2480),
            .I(\uart.stateZ0Z_0 ));
    InMux I__312 (
            .O(N__2477),
            .I(N__2469));
    InMux I__311 (
            .O(N__2476),
            .I(N__2469));
    CascadeMux I__310 (
            .O(N__2475),
            .I(N__2466));
    InMux I__309 (
            .O(N__2474),
            .I(N__2460));
    LocalMux I__308 (
            .O(N__2469),
            .I(N__2457));
    InMux I__307 (
            .O(N__2466),
            .I(N__2448));
    InMux I__306 (
            .O(N__2465),
            .I(N__2448));
    InMux I__305 (
            .O(N__2464),
            .I(N__2448));
    InMux I__304 (
            .O(N__2463),
            .I(N__2448));
    LocalMux I__303 (
            .O(N__2460),
            .I(\uart.N_175 ));
    Odrv4 I__302 (
            .O(N__2457),
            .I(\uart.N_175 ));
    LocalMux I__301 (
            .O(N__2448),
            .I(\uart.N_175 ));
    CascadeMux I__300 (
            .O(N__2441),
            .I(\uart.data_Auxce_0_6_cascade_ ));
    CEMux I__299 (
            .O(N__2438),
            .I(N__2435));
    LocalMux I__298 (
            .O(N__2435),
            .I(N__2432));
    Odrv4 I__297 (
            .O(N__2432),
            .I(\uart.N_114_0 ));
    InMux I__296 (
            .O(N__2429),
            .I(N__2426));
    LocalMux I__295 (
            .O(N__2426),
            .I(\uart.data_Aux_esr_RNO_0Z0Z_5 ));
    InMux I__294 (
            .O(N__2423),
            .I(N__2420));
    LocalMux I__293 (
            .O(N__2420),
            .I(N__2417));
    Odrv12 I__292 (
            .O(N__2417),
            .I(\uart.data_AuxZ0Z_5 ));
    CEMux I__291 (
            .O(N__2414),
            .I(N__2411));
    LocalMux I__290 (
            .O(N__2411),
            .I(N__2408));
    Odrv4 I__289 (
            .O(N__2408),
            .I(\uart.N_115_0 ));
    CascadeMux I__288 (
            .O(N__2405),
            .I(\uart.data_Aux_esr_RNO_0Z0Z_0_cascade_ ));
    CEMux I__287 (
            .O(N__2402),
            .I(N__2399));
    LocalMux I__286 (
            .O(N__2399),
            .I(N__2396));
    Odrv4 I__285 (
            .O(N__2396),
            .I(\uart.N_120_0 ));
    InMux I__284 (
            .O(N__2393),
            .I(N__2389));
    InMux I__283 (
            .O(N__2392),
            .I(N__2386));
    LocalMux I__282 (
            .O(N__2389),
            .I(\uart.data_Auxce_0_0 ));
    LocalMux I__281 (
            .O(N__2386),
            .I(\uart.data_Auxce_0_0 ));
    CascadeMux I__280 (
            .O(N__2381),
            .I(\uart.data_Aux_esr_RNO_0Z0Z_1_cascade_ ));
    InMux I__279 (
            .O(N__2378),
            .I(N__2375));
    LocalMux I__278 (
            .O(N__2375),
            .I(N__2372));
    Odrv4 I__277 (
            .O(N__2372),
            .I(\uart.data_AuxZ0Z_1 ));
    CEMux I__276 (
            .O(N__2369),
            .I(N__2366));
    LocalMux I__275 (
            .O(N__2366),
            .I(N__2363));
    Odrv4 I__274 (
            .O(N__2363),
            .I(\uart.N_119_0 ));
    InMux I__273 (
            .O(N__2360),
            .I(N__2357));
    LocalMux I__272 (
            .O(N__2357),
            .I(\uart.data_Auxce_0_2 ));
    CascadeMux I__271 (
            .O(N__2354),
            .I(\uart.data_Aux_esr_RNO_0Z0Z_3_cascade_ ));
    CascadeMux I__270 (
            .O(N__2351),
            .I(\uart.data_Aux_esr_RNO_0Z0Z_4_cascade_ ));
    InMux I__269 (
            .O(N__2348),
            .I(N__2345));
    LocalMux I__268 (
            .O(N__2345),
            .I(uart_data_4));
    InMux I__267 (
            .O(N__2342),
            .I(N__2338));
    InMux I__266 (
            .O(N__2341),
            .I(N__2335));
    LocalMux I__265 (
            .O(N__2338),
            .I(uart_data_5));
    LocalMux I__264 (
            .O(N__2335),
            .I(uart_data_5));
    InMux I__263 (
            .O(N__2330),
            .I(N__2327));
    LocalMux I__262 (
            .O(N__2327),
            .I(N__2324));
    Span4Mux_s2_v I__261 (
            .O(N__2324),
            .I(N__2321));
    Odrv4 I__260 (
            .O(N__2321),
            .I(\uart.data_AuxZ0Z_6 ));
    InMux I__259 (
            .O(N__2318),
            .I(N__2315));
    LocalMux I__258 (
            .O(N__2315),
            .I(uart_data_6));
    InMux I__257 (
            .O(N__2312),
            .I(N__2309));
    LocalMux I__256 (
            .O(N__2309),
            .I(N__2306));
    Odrv4 I__255 (
            .O(N__2306),
            .I(\uart.data_AuxZ0Z_7 ));
    CascadeMux I__254 (
            .O(N__2303),
            .I(N__2299));
    InMux I__253 (
            .O(N__2302),
            .I(N__2296));
    InMux I__252 (
            .O(N__2299),
            .I(N__2293));
    LocalMux I__251 (
            .O(N__2296),
            .I(uart_data_7));
    LocalMux I__250 (
            .O(N__2293),
            .I(uart_data_7));
    CascadeMux I__249 (
            .O(N__2288),
            .I(\uart.N_147_0_0_cascade_ ));
    CascadeMux I__248 (
            .O(N__2285),
            .I(\uart.g3_1_0_cascade_ ));
    InMux I__247 (
            .O(N__2282),
            .I(N__2279));
    LocalMux I__246 (
            .O(N__2279),
            .I(N__2276));
    Span4Mux_s2_v I__245 (
            .O(N__2276),
            .I(N__2273));
    Odrv4 I__244 (
            .O(N__2273),
            .I(\uart.g0_4_0 ));
    CascadeMux I__243 (
            .O(N__2270),
            .I(\uart.N_175_cascade_ ));
    CascadeMux I__242 (
            .O(N__2267),
            .I(N__2262));
    InMux I__241 (
            .O(N__2266),
            .I(N__2255));
    InMux I__240 (
            .O(N__2265),
            .I(N__2255));
    InMux I__239 (
            .O(N__2262),
            .I(N__2248));
    InMux I__238 (
            .O(N__2261),
            .I(N__2248));
    InMux I__237 (
            .O(N__2260),
            .I(N__2248));
    LocalMux I__236 (
            .O(N__2255),
            .I(\uart_frame_decoder.state_1Z0Z_1 ));
    LocalMux I__235 (
            .O(N__2248),
            .I(\uart_frame_decoder.state_1Z0Z_1 ));
    IoInMux I__234 (
            .O(N__2243),
            .I(N__2240));
    LocalMux I__233 (
            .O(N__2240),
            .I(uart_frame_decoder_N_129_i));
    CascadeMux I__232 (
            .O(N__2237),
            .I(\uart_frame_decoder.state_1_srsts_i_i_a2_3_0Z0Z_0_cascade_ ));
    InMux I__231 (
            .O(N__2234),
            .I(N__2228));
    InMux I__230 (
            .O(N__2233),
            .I(N__2228));
    LocalMux I__229 (
            .O(N__2228),
            .I(\uart_frame_decoder.N_67 ));
    InMux I__228 (
            .O(N__2225),
            .I(N__2222));
    LocalMux I__227 (
            .O(N__2222),
            .I(\uart_frame_decoder.N_61 ));
    CascadeMux I__226 (
            .O(N__2219),
            .I(\uart_frame_decoder.N_67_cascade_ ));
    InMux I__225 (
            .O(N__2216),
            .I(N__2212));
    InMux I__224 (
            .O(N__2215),
            .I(N__2209));
    LocalMux I__223 (
            .O(N__2212),
            .I(\uart_frame_decoder.state_1_srsts_0_i_a2_0_0_2 ));
    LocalMux I__222 (
            .O(N__2209),
            .I(\uart_frame_decoder.state_1_srsts_0_i_a2_0_0_2 ));
    InMux I__221 (
            .O(N__2204),
            .I(N__2201));
    LocalMux I__220 (
            .O(N__2201),
            .I(N__2198));
    Odrv4 I__219 (
            .O(N__2198),
            .I(\uart.data_AuxZ0Z_0 ));
    InMux I__218 (
            .O(N__2195),
            .I(N__2191));
    InMux I__217 (
            .O(N__2194),
            .I(N__2188));
    LocalMux I__216 (
            .O(N__2191),
            .I(uart_data_0));
    LocalMux I__215 (
            .O(N__2188),
            .I(uart_data_0));
    InMux I__214 (
            .O(N__2183),
            .I(N__2180));
    LocalMux I__213 (
            .O(N__2180),
            .I(N__2177));
    Odrv4 I__212 (
            .O(N__2177),
            .I(uart_data_1));
    InMux I__211 (
            .O(N__2174),
            .I(N__2171));
    LocalMux I__210 (
            .O(N__2171),
            .I(\uart.data_AuxZ0Z_2 ));
    InMux I__209 (
            .O(N__2168),
            .I(N__2164));
    InMux I__208 (
            .O(N__2167),
            .I(N__2161));
    LocalMux I__207 (
            .O(N__2164),
            .I(uart_data_2));
    LocalMux I__206 (
            .O(N__2161),
            .I(uart_data_2));
    InMux I__205 (
            .O(N__2156),
            .I(N__2153));
    LocalMux I__204 (
            .O(N__2153),
            .I(N__2150));
    Odrv4 I__203 (
            .O(N__2150),
            .I(uart_data_3));
    CascadeMux I__202 (
            .O(N__2147),
            .I(\uart.data_Aux_esr_RNO_0Z0Z_2_cascade_ ));
    CEMux I__201 (
            .O(N__2144),
            .I(N__2141));
    LocalMux I__200 (
            .O(N__2141),
            .I(N__2138));
    Odrv4 I__199 (
            .O(N__2138),
            .I(\uart.N_118_0 ));
    CascadeMux I__198 (
            .O(N__2135),
            .I(\uart_frame_decoder.state_1_srsts_0_i_a2_0_0_1Z0Z_2_cascade_ ));
    InMux I__197 (
            .O(N__2132),
            .I(N__2129));
    LocalMux I__196 (
            .O(N__2129),
            .I(\uart_frame_decoder.N_49 ));
    CascadeMux I__195 (
            .O(N__2126),
            .I(\uart_frame_decoder.N_58_4_cascade_ ));
    InMux I__194 (
            .O(N__2123),
            .I(N__2120));
    LocalMux I__193 (
            .O(N__2120),
            .I(N__2117));
    Odrv4 I__192 (
            .O(N__2117),
            .I(\uart_frame_decoder.N_32_i_1 ));
    CascadeMux I__191 (
            .O(N__2114),
            .I(\uart.state_0_sqmuxa_1_d_cascade_ ));
    CascadeMux I__190 (
            .O(N__2111),
            .I(\uart.m13_0_0_o2_2_cascade_ ));
    CascadeMux I__189 (
            .O(N__2108),
            .I(\uart.N_10_cascade_ ));
    CascadeMux I__188 (
            .O(N__2105),
            .I(\uart.data_Auxce_0_2_cascade_ ));
    CascadeMux I__187 (
            .O(N__2102),
            .I(\uart_frame_decoder.N_43_cascade_ ));
    CascadeMux I__186 (
            .O(N__2099),
            .I(\uart_frame_decoder.state_1_srsts_i_i_0_0_cascade_ ));
    IoInMux I__185 (
            .O(N__2096),
            .I(N__2093));
    LocalMux I__184 (
            .O(N__2093),
            .I(N__2090));
    Span4Mux_s0_v I__183 (
            .O(N__2090),
            .I(N__2087));
    Odrv4 I__182 (
            .O(N__2087),
            .I(uart_frame_decoder_N_131_i));
    CascadeMux I__181 (
            .O(N__2084),
            .I(N__2081));
    InMux I__180 (
            .O(N__2081),
            .I(N__2078));
    LocalMux I__179 (
            .O(N__2078),
            .I(\uart_frame_decoder.state_1Z0Z_0 ));
    InMux I__178 (
            .O(N__2075),
            .I(N__2072));
    LocalMux I__177 (
            .O(N__2072),
            .I(\uart_frame_decoder.state_1_srsts_0_i_1_1 ));
    InMux I__176 (
            .O(N__2069),
            .I(N__2066));
    LocalMux I__175 (
            .O(N__2066),
            .I(\uart_frame_decoder.N_58_4 ));
    defparam IN_MUX_bfv_12_2_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_2_0_));
    defparam IN_MUX_bfv_12_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_3_0_ (
            .carryinitin(\reset_module_System.count_1_cry_8 ),
            .carryinitout(bfn_12_3_0_));
    defparam IN_MUX_bfv_12_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_4_0_ (
            .carryinitin(\reset_module_System.count_1_cry_16 ),
            .carryinitout(bfn_12_4_0_));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNO_2_0_LC_7_1_0 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNO_2_0_LC_7_1_0 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNO_2_0_LC_7_1_0 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \uart_frame_decoder.state_1_RNO_2_0_LC_7_1_0  (
            .in0(N__3773),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2260),
            .lcout(),
            .ltout(\uart_frame_decoder.N_43_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNO_1_0_LC_7_1_1 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNO_1_0_LC_7_1_1 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNO_1_0_LC_7_1_1 .LUT_INIT=16'b0101010100010000;
    LogicCell40 \uart_frame_decoder.state_1_RNO_1_0_LC_7_1_1  (
            .in0(N__3381),
            .in1(N__4914),
            .in2(N__2102),
            .in3(N__2132),
            .lcout(),
            .ltout(\uart_frame_decoder.state_1_srsts_i_i_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_0_LC_7_1_2 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_0_LC_7_1_2 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.state_1_0_LC_7_1_2 .LUT_INIT=16'b0000001100000111;
    LogicCell40 \uart_frame_decoder.state_1_0_LC_7_1_2  (
            .in0(N__2215),
            .in1(N__2233),
            .in2(N__2099),
            .in3(N__2123),
            .lcout(\uart_frame_decoder.state_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4814),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_1_LC_7_1_3 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_1_LC_7_1_3 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.state_1_1_LC_7_1_3 .LUT_INIT=16'b0011000010001000;
    LogicCell40 \uart_frame_decoder.state_1_1_LC_7_1_3  (
            .in0(N__2234),
            .in1(N__4915),
            .in2(N__2267),
            .in3(N__2075),
            .lcout(\uart_frame_decoder.state_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4814),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_esr_RNI7FFE_4_LC_7_1_4 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_esr_RNI7FFE_4_LC_7_1_4 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_esr_RNI7FFE_4_LC_7_1_4 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \uart_frame_decoder.state_1_esr_RNI7FFE_4_LC_7_1_4  (
            .in0(N__3775),
            .in1(N__3302),
            .in2(_gnd_net_),
            .in3(N__3277),
            .lcout(uart_frame_decoder_N_131_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNO_0_1_LC_7_1_5 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNO_0_1_LC_7_1_5 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNO_0_1_LC_7_1_5 .LUT_INIT=16'b0001110111011101;
    LogicCell40 \uart_frame_decoder.state_1_RNO_0_1_LC_7_1_5  (
            .in0(N__3380),
            .in1(N__4913),
            .in2(N__2084),
            .in3(N__2069),
            .lcout(\uart_frame_decoder.state_1_srsts_0_i_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_srsts_0_i_a2_0_4_1_LC_7_1_6 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_srsts_0_i_a2_0_4_1_LC_7_1_6 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_srsts_0_i_a2_0_4_1_LC_7_1_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uart_frame_decoder.state_1_srsts_0_i_a2_0_4_1_LC_7_1_6  (
            .in0(N__2341),
            .in1(N__2167),
            .in2(N__2303),
            .in3(N__2194),
            .lcout(\uart_frame_decoder.N_58_4 ),
            .ltout(\uart_frame_decoder.N_58_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNO_0_0_LC_7_1_7 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNO_0_0_LC_7_1_7 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNO_0_0_LC_7_1_7 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \uart_frame_decoder.state_1_RNO_0_0_LC_7_1_7  (
            .in0(N__2261),
            .in1(N__4912),
            .in2(N__2126),
            .in3(N__3774),
            .lcout(\uart_frame_decoder.N_32_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_esr_2_LC_7_2_0 .C_ON=1'b0;
    defparam \uart.data_Aux_esr_2_LC_7_2_0 .SEQ_MODE=4'b1000;
    defparam \uart.data_Aux_esr_2_LC_7_2_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart.data_Aux_esr_2_LC_7_2_0  (
            .in0(N__5134),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uart.data_AuxZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4812),
            .ce(N__2144),
            .sr(N__2739));
    defparam \uart.bit_Count_RNO_0_0_LC_7_3_0 .C_ON=1'b0;
    defparam \uart.bit_Count_RNO_0_0_LC_7_3_0 .SEQ_MODE=4'b0000;
    defparam \uart.bit_Count_RNO_0_0_LC_7_3_0 .LUT_INIT=16'b1111111111010101;
    LogicCell40 \uart.bit_Count_RNO_0_0_LC_7_3_0  (
            .in0(N__3639),
            .in1(N__3551),
            .in2(N__2582),
            .in3(N__4126),
            .lcout(),
            .ltout(\uart.state_0_sqmuxa_1_d_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.bit_Count_0_LC_7_3_1 .C_ON=1'b0;
    defparam \uart.bit_Count_0_LC_7_3_1 .SEQ_MODE=4'b1000;
    defparam \uart.bit_Count_0_LC_7_3_1 .LUT_INIT=16'b0110110001001100;
    LogicCell40 \uart.bit_Count_0_LC_7_3_1  (
            .in0(N__3428),
            .in1(N__3147),
            .in2(N__2114),
            .in3(N__2501),
            .lcout(\uart.bit_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4809),
            .ce(),
            .sr(N__4724));
    defparam \uart.bit_Count_RNO_2_2_LC_7_3_2 .C_ON=1'b0;
    defparam \uart.bit_Count_RNO_2_2_LC_7_3_2 .SEQ_MODE=4'b0000;
    defparam \uart.bit_Count_RNO_2_2_LC_7_3_2 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \uart.bit_Count_RNO_2_2_LC_7_3_2  (
            .in0(N__3011),
            .in1(N__3135),
            .in2(_gnd_net_),
            .in3(N__4313),
            .lcout(),
            .ltout(\uart.m13_0_0_o2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.bit_Count_RNO_0_2_LC_7_3_3 .C_ON=1'b0;
    defparam \uart.bit_Count_RNO_0_2_LC_7_3_3 .SEQ_MODE=4'b0000;
    defparam \uart.bit_Count_RNO_0_2_LC_7_3_3 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \uart.bit_Count_RNO_0_2_LC_7_3_3  (
            .in0(N__2894),
            .in1(N__3935),
            .in2(N__2111),
            .in3(N__5061),
            .lcout(),
            .ltout(\uart.N_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.bit_Count_2_LC_7_3_4 .C_ON=1'b0;
    defparam \uart.bit_Count_2_LC_7_3_4 .SEQ_MODE=4'b1000;
    defparam \uart.bit_Count_2_LC_7_3_4 .LUT_INIT=16'b1110000000001110;
    LogicCell40 \uart.bit_Count_2_LC_7_3_4  (
            .in0(N__5062),
            .in1(N__3641),
            .in2(N__2108),
            .in3(N__3073),
            .lcout(\uart.bit_CountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4809),
            .ce(),
            .sr(N__4724));
    defparam \uart.bit_Count_RNILKM9_0_2_LC_7_3_5 .C_ON=1'b0;
    defparam \uart.bit_Count_RNILKM9_0_2_LC_7_3_5 .SEQ_MODE=4'b0000;
    defparam \uart.bit_Count_RNILKM9_0_2_LC_7_3_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uart.bit_Count_RNILKM9_0_2_LC_7_3_5  (
            .in0(_gnd_net_),
            .in1(N__3061),
            .in2(_gnd_net_),
            .in3(N__3010),
            .lcout(\uart.data_Auxce_0_2 ),
            .ltout(\uart.data_Auxce_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_esr_RNO_0_2_LC_7_3_6 .C_ON=1'b0;
    defparam \uart.data_Aux_esr_RNO_0_2_LC_7_3_6 .SEQ_MODE=4'b0000;
    defparam \uart.data_Aux_esr_RNO_0_2_LC_7_3_6 .LUT_INIT=16'b0101000001000000;
    LogicCell40 \uart.data_Aux_esr_RNO_0_2_LC_7_3_6  (
            .in0(N__3146),
            .in1(N__2847),
            .in2(N__2105),
            .in3(N__2474),
            .lcout(),
            .ltout(\uart.data_Aux_esr_RNO_0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_esr_RNO_2_LC_7_3_7 .C_ON=1'b0;
    defparam \uart.data_Aux_esr_RNO_2_LC_7_3_7 .SEQ_MODE=4'b0000;
    defparam \uart.data_Aux_esr_RNO_2_LC_7_3_7 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \uart.data_Aux_esr_RNO_2_LC_7_3_7  (
            .in0(N__2716),
            .in1(_gnd_net_),
            .in2(N__2147),
            .in3(_gnd_net_),
            .lcout(\uart.N_118_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_esr_0_LC_7_4_0 .C_ON=1'b0;
    defparam \uart.data_Aux_esr_0_LC_7_4_0 .SEQ_MODE=4'b1000;
    defparam \uart.data_Aux_esr_0_LC_7_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart.data_Aux_esr_0_LC_7_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5157),
            .lcout(\uart.data_AuxZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4806),
            .ce(N__2402),
            .sr(N__2740));
    defparam \uart.bit_Count_RNIETHE_2_LC_7_5_1 .C_ON=1'b0;
    defparam \uart.bit_Count_RNIETHE_2_LC_7_5_1 .SEQ_MODE=4'b0000;
    defparam \uart.bit_Count_RNIETHE_2_LC_7_5_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uart.bit_Count_RNIETHE_2_LC_7_5_1  (
            .in0(N__3158),
            .in1(N__3076),
            .in2(_gnd_net_),
            .in3(N__3025),
            .lcout(\uart.N_177 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_esr_7_LC_7_5_3 .C_ON=1'b0;
    defparam \uart.data_Aux_esr_7_LC_7_5_3 .SEQ_MODE=4'b1000;
    defparam \uart.data_Aux_esr_7_LC_7_5_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart.data_Aux_esr_7_LC_7_5_3  (
            .in0(N__5161),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uart.data_AuxZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4803),
            .ce(N__2510),
            .sr(N__2744));
    defparam \uart.bit_Count_RNO_0_1_LC_7_5_6 .C_ON=1'b0;
    defparam \uart.bit_Count_RNO_0_1_LC_7_5_6 .SEQ_MODE=4'b0000;
    defparam \uart.bit_Count_RNO_0_1_LC_7_5_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \uart.bit_Count_RNO_0_1_LC_7_5_6  (
            .in0(_gnd_net_),
            .in1(N__3427),
            .in2(_gnd_net_),
            .in3(N__2497),
            .lcout(\uart.g0_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_esr_6_LC_7_6_0 .C_ON=1'b0;
    defparam \uart.data_Aux_esr_6_LC_7_6_0 .SEQ_MODE=4'b1000;
    defparam \uart.data_Aux_esr_6_LC_7_6_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart.data_Aux_esr_6_LC_7_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5162),
            .lcout(\uart.data_AuxZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4798),
            .ce(N__2438),
            .sr(N__2741));
    defparam \uart_frame_decoder.state_1_srsts_0_i_a2_0_0_1_2_LC_8_1_0 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_srsts_0_i_a2_0_0_1_2_LC_8_1_0 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_srsts_0_i_a2_0_0_1_2_LC_8_1_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \uart_frame_decoder.state_1_srsts_0_i_a2_0_0_1_2_LC_8_1_0  (
            .in0(_gnd_net_),
            .in1(N__2342),
            .in2(_gnd_net_),
            .in3(N__2168),
            .lcout(),
            .ltout(\uart_frame_decoder.state_1_srsts_0_i_a2_0_0_1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNI5BVV_1_LC_8_1_1 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNI5BVV_1_LC_8_1_1 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNI5BVV_1_LC_8_1_1 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \uart_frame_decoder.state_1_RNI5BVV_1_LC_8_1_1  (
            .in0(N__2265),
            .in1(N__2195),
            .in2(N__2135),
            .in3(N__2302),
            .lcout(\uart_frame_decoder.state_1_srsts_0_i_a2_0_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNO_0_2_LC_8_1_2 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNO_0_2_LC_8_1_2 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNO_0_2_LC_8_1_2 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \uart_frame_decoder.state_1_RNO_0_2_LC_8_1_2  (
            .in0(N__3735),
            .in1(N__4910),
            .in2(_gnd_net_),
            .in3(N__3379),
            .lcout(\uart_frame_decoder.N_61 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNO_3_0_LC_8_1_3 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNO_3_0_LC_8_1_3 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNO_3_0_LC_8_1_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \uart_frame_decoder.state_1_RNO_3_0_LC_8_1_3  (
            .in0(N__3301),
            .in1(N__3799),
            .in2(N__3278),
            .in3(N__3734),
            .lcout(\uart_frame_decoder.N_49 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_esr_RNI19FE_3_LC_8_1_4 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_esr_RNI19FE_3_LC_8_1_4 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_esr_RNI19FE_3_LC_8_1_4 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \uart_frame_decoder.state_1_esr_RNI19FE_3_LC_8_1_4  (
            .in0(N__3800),
            .in1(N__3275),
            .in2(_gnd_net_),
            .in3(N__2266),
            .lcout(uart_frame_decoder_N_129_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_srsts_i_i_a2_3_0_0_LC_8_1_5 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_srsts_i_i_a2_3_0_0_LC_8_1_5 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_srsts_i_i_a2_3_0_0_LC_8_1_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \uart_frame_decoder.state_1_srsts_i_i_a2_3_0_0_LC_8_1_5  (
            .in0(_gnd_net_),
            .in1(N__2348),
            .in2(_gnd_net_),
            .in3(N__4247),
            .lcout(),
            .ltout(\uart_frame_decoder.state_1_srsts_i_i_a2_3_0Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_srsts_i_i_a2_3_0_LC_8_1_6 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_srsts_i_i_a2_3_0_LC_8_1_6 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_srsts_i_i_a2_3_0_LC_8_1_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uart_frame_decoder.state_1_srsts_i_i_a2_3_0_LC_8_1_6  (
            .in0(N__2156),
            .in1(N__2318),
            .in2(N__2237),
            .in3(N__2183),
            .lcout(\uart_frame_decoder.N_67 ),
            .ltout(\uart_frame_decoder.N_67_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_2_LC_8_1_7 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_2_LC_8_1_7 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.state_1_2_LC_8_1_7 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \uart_frame_decoder.state_1_2_LC_8_1_7  (
            .in0(N__4911),
            .in1(N__2225),
            .in2(N__2219),
            .in3(N__2216),
            .lcout(\uart_frame_decoder.state_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4813),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_esr_0_LC_8_2_0 .C_ON=1'b0;
    defparam \uart.data_esr_0_LC_8_2_0 .SEQ_MODE=4'b1000;
    defparam \uart.data_esr_0_LC_8_2_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart.data_esr_0_LC_8_2_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2204),
            .lcout(uart_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4810),
            .ce(N__2528),
            .sr(N__2543));
    defparam \uart.data_esr_1_LC_8_2_1 .C_ON=1'b0;
    defparam \uart.data_esr_1_LC_8_2_1 .SEQ_MODE=4'b1000;
    defparam \uart.data_esr_1_LC_8_2_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart.data_esr_1_LC_8_2_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2378),
            .lcout(uart_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4810),
            .ce(N__2528),
            .sr(N__2543));
    defparam \uart.data_esr_2_LC_8_2_2 .C_ON=1'b0;
    defparam \uart.data_esr_2_LC_8_2_2 .SEQ_MODE=4'b1000;
    defparam \uart.data_esr_2_LC_8_2_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart.data_esr_2_LC_8_2_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2174),
            .lcout(uart_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4810),
            .ce(N__2528),
            .sr(N__2543));
    defparam \uart.data_esr_3_LC_8_2_3 .C_ON=1'b0;
    defparam \uart.data_esr_3_LC_8_2_3 .SEQ_MODE=4'b1000;
    defparam \uart.data_esr_3_LC_8_2_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart.data_esr_3_LC_8_2_3  (
            .in0(N__2786),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(uart_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4810),
            .ce(N__2528),
            .sr(N__2543));
    defparam \uart.data_esr_4_LC_8_2_4 .C_ON=1'b0;
    defparam \uart.data_esr_4_LC_8_2_4 .SEQ_MODE=4'b1000;
    defparam \uart.data_esr_4_LC_8_2_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart.data_esr_4_LC_8_2_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2768),
            .lcout(uart_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4810),
            .ce(N__2528),
            .sr(N__2543));
    defparam \uart.data_esr_5_LC_8_2_5 .C_ON=1'b0;
    defparam \uart.data_esr_5_LC_8_2_5 .SEQ_MODE=4'b1000;
    defparam \uart.data_esr_5_LC_8_2_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart.data_esr_5_LC_8_2_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2423),
            .lcout(uart_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4810),
            .ce(N__2528),
            .sr(N__2543));
    defparam \uart.data_esr_6_LC_8_2_6 .C_ON=1'b0;
    defparam \uart.data_esr_6_LC_8_2_6 .SEQ_MODE=4'b1000;
    defparam \uart.data_esr_6_LC_8_2_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart.data_esr_6_LC_8_2_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2330),
            .lcout(uart_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4810),
            .ce(N__2528),
            .sr(N__2543));
    defparam \uart.data_esr_7_LC_8_2_7 .C_ON=1'b0;
    defparam \uart.data_esr_7_LC_8_2_7 .SEQ_MODE=4'b1000;
    defparam \uart.data_esr_7_LC_8_2_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart.data_esr_7_LC_8_2_7  (
            .in0(N__2312),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(uart_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4810),
            .ce(N__2528),
            .sr(N__2543));
    defparam \uart.bit_Count_RNO_3_1_LC_8_3_0 .C_ON=1'b0;
    defparam \uart.bit_Count_RNO_3_1_LC_8_3_0 .SEQ_MODE=4'b0000;
    defparam \uart.bit_Count_RNO_3_1_LC_8_3_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart.bit_Count_RNO_3_1_LC_8_3_0  (
            .in0(_gnd_net_),
            .in1(N__3934),
            .in2(_gnd_net_),
            .in3(N__4312),
            .lcout(),
            .ltout(\uart.N_147_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.bit_Count_RNO_1_1_LC_8_3_1 .C_ON=1'b0;
    defparam \uart.bit_Count_RNO_1_1_LC_8_3_1 .SEQ_MODE=4'b0000;
    defparam \uart.bit_Count_RNO_1_1_LC_8_3_1 .LUT_INIT=16'b0000000010100010;
    LogicCell40 \uart.bit_Count_RNO_1_1_LC_8_3_1  (
            .in0(N__3149),
            .in1(N__3640),
            .in2(N__2288),
            .in3(N__5063),
            .lcout(),
            .ltout(\uart.g3_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.bit_Count_1_LC_8_3_2 .C_ON=1'b0;
    defparam \uart.bit_Count_1_LC_8_3_2 .SEQ_MODE=4'b1000;
    defparam \uart.bit_Count_1_LC_8_3_2 .LUT_INIT=16'b0010001001101010;
    LogicCell40 \uart.bit_Count_1_LC_8_3_2  (
            .in0(N__3009),
            .in1(N__3497),
            .in2(N__2285),
            .in3(N__2282),
            .lcout(\uart.bit_CountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4807),
            .ce(),
            .sr(N__4723));
    defparam \uart.bit_Count_RNILKM9_2_LC_8_3_3 .C_ON=1'b0;
    defparam \uart.bit_Count_RNILKM9_2_LC_8_3_3 .SEQ_MODE=4'b0000;
    defparam \uart.bit_Count_RNILKM9_2_LC_8_3_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \uart.bit_Count_RNILKM9_2_LC_8_3_3  (
            .in0(_gnd_net_),
            .in1(N__3059),
            .in2(_gnd_net_),
            .in3(N__3007),
            .lcout(\uart.data_Auxce_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_RNI3UCP2_4_LC_8_3_4 .C_ON=1'b0;
    defparam \uart.timer_Count_RNI3UCP2_4_LC_8_3_4 .SEQ_MODE=4'b0000;
    defparam \uart.timer_Count_RNI3UCP2_4_LC_8_3_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \uart.timer_Count_RNI3UCP2_4_LC_8_3_4  (
            .in0(N__4119),
            .in1(N__2557),
            .in2(N__3549),
            .in3(N__3215),
            .lcout(\uart.N_175 ),
            .ltout(\uart.N_175_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_esr_RNO_0_0_LC_8_3_5 .C_ON=1'b0;
    defparam \uart.data_Aux_esr_RNO_0_0_LC_8_3_5 .SEQ_MODE=4'b0000;
    defparam \uart.data_Aux_esr_RNO_0_0_LC_8_3_5 .LUT_INIT=16'b0011001000000000;
    LogicCell40 \uart.data_Aux_esr_RNO_0_0_LC_8_3_5  (
            .in0(N__2841),
            .in1(N__3148),
            .in2(N__2270),
            .in3(N__2392),
            .lcout(),
            .ltout(\uart.data_Aux_esr_RNO_0Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_esr_RNO_0_LC_8_3_6 .C_ON=1'b0;
    defparam \uart.data_Aux_esr_RNO_0_LC_8_3_6 .SEQ_MODE=4'b0000;
    defparam \uart.data_Aux_esr_RNO_0_LC_8_3_6 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \uart.data_Aux_esr_RNO_0_LC_8_3_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2405),
            .in3(N__2682),
            .lcout(\uart.N_120_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.bit_Count_RNILKM9_1_2_LC_8_3_7 .C_ON=1'b0;
    defparam \uart.bit_Count_RNILKM9_1_2_LC_8_3_7 .SEQ_MODE=4'b0000;
    defparam \uart.bit_Count_RNILKM9_1_2_LC_8_3_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \uart.bit_Count_RNILKM9_1_2_LC_8_3_7  (
            .in0(_gnd_net_),
            .in1(N__3060),
            .in2(_gnd_net_),
            .in3(N__3008),
            .lcout(\uart.data_Auxce_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_esr_RNO_0_1_LC_8_4_0 .C_ON=1'b0;
    defparam \uart.data_Aux_esr_RNO_0_1_LC_8_4_0 .SEQ_MODE=4'b0000;
    defparam \uart.data_Aux_esr_RNO_0_1_LC_8_4_0 .LUT_INIT=16'b1100100000000000;
    LogicCell40 \uart.data_Aux_esr_RNO_0_1_LC_8_4_0  (
            .in0(N__2837),
            .in1(N__3139),
            .in2(N__2475),
            .in3(N__2393),
            .lcout(),
            .ltout(\uart.data_Aux_esr_RNO_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_esr_RNO_1_LC_8_4_1 .C_ON=1'b0;
    defparam \uart.data_Aux_esr_RNO_1_LC_8_4_1 .SEQ_MODE=4'b0000;
    defparam \uart.data_Aux_esr_RNO_1_LC_8_4_1 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \uart.data_Aux_esr_RNO_1_LC_8_4_1  (
            .in0(N__2694),
            .in1(_gnd_net_),
            .in2(N__2381),
            .in3(_gnd_net_),
            .lcout(\uart.N_119_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_esr_1_LC_8_4_2 .C_ON=1'b0;
    defparam \uart.data_Aux_esr_1_LC_8_4_2 .SEQ_MODE=4'b1000;
    defparam \uart.data_Aux_esr_1_LC_8_4_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart.data_Aux_esr_1_LC_8_4_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5156),
            .lcout(\uart.data_AuxZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4804),
            .ce(N__2369),
            .sr(N__2742));
    defparam \uart.data_Aux_esr_RNO_0_3_LC_8_4_3 .C_ON=1'b0;
    defparam \uart.data_Aux_esr_RNO_0_3_LC_8_4_3 .SEQ_MODE=4'b0000;
    defparam \uart.data_Aux_esr_RNO_0_3_LC_8_4_3 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \uart.data_Aux_esr_RNO_0_3_LC_8_4_3  (
            .in0(N__2360),
            .in1(N__2836),
            .in2(N__3160),
            .in3(N__2465),
            .lcout(),
            .ltout(\uart.data_Aux_esr_RNO_0Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_esr_RNO_3_LC_8_4_4 .C_ON=1'b0;
    defparam \uart.data_Aux_esr_RNO_3_LC_8_4_4 .SEQ_MODE=4'b0000;
    defparam \uart.data_Aux_esr_RNO_3_LC_8_4_4 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \uart.data_Aux_esr_RNO_3_LC_8_4_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2354),
            .in3(N__2695),
            .lcout(\uart.N_117_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_esr_RNO_0_4_LC_8_4_5 .C_ON=1'b0;
    defparam \uart.data_Aux_esr_RNO_0_4_LC_8_4_5 .SEQ_MODE=4'b0000;
    defparam \uart.data_Aux_esr_RNO_0_4_LC_8_4_5 .LUT_INIT=16'b0000101000001000;
    LogicCell40 \uart.data_Aux_esr_RNO_0_4_LC_8_4_5  (
            .in0(N__2519),
            .in1(N__2835),
            .in2(N__3161),
            .in3(N__2464),
            .lcout(),
            .ltout(\uart.data_Aux_esr_RNO_0Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_esr_RNO_4_LC_8_4_6 .C_ON=1'b0;
    defparam \uart.data_Aux_esr_RNO_4_LC_8_4_6 .SEQ_MODE=4'b0000;
    defparam \uart.data_Aux_esr_RNO_4_LC_8_4_6 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \uart.data_Aux_esr_RNO_4_LC_8_4_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2351),
            .in3(N__2696),
            .lcout(\uart.N_116_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_esr_RNO_0_5_LC_8_4_7 .C_ON=1'b0;
    defparam \uart.data_Aux_esr_RNO_0_5_LC_8_4_7 .SEQ_MODE=4'b0000;
    defparam \uart.data_Aux_esr_RNO_0_5_LC_8_4_7 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \uart.data_Aux_esr_RNO_0_5_LC_8_4_7  (
            .in0(N__2518),
            .in1(N__2834),
            .in2(N__3159),
            .in3(N__2463),
            .lcout(\uart.data_Aux_esr_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_0_LC_8_5_0 .C_ON=1'b0;
    defparam \uart.state_0_LC_8_5_0 .SEQ_MODE=4'b1000;
    defparam \uart.state_0_LC_8_5_0 .LUT_INIT=16'b1111111111110010;
    LogicCell40 \uart.state_0_LC_8_5_0  (
            .in0(N__2485),
            .in1(N__5158),
            .in2(N__3386),
            .in3(N__2801),
            .lcout(\uart.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4799),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_esr_RNO_7_LC_8_5_1 .C_ON=1'b0;
    defparam \uart.data_Aux_esr_RNO_7_LC_8_5_1 .SEQ_MODE=4'b0000;
    defparam \uart.data_Aux_esr_RNO_7_LC_8_5_1 .LUT_INIT=16'b1111111010101010;
    LogicCell40 \uart.data_Aux_esr_RNO_7_LC_8_5_1  (
            .in0(N__2728),
            .in1(N__2476),
            .in2(N__2852),
            .in3(N__3400),
            .lcout(\uart.N_113_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.bit_Count_RNI4ENK_2_LC_8_5_3 .C_ON=1'b0;
    defparam \uart.bit_Count_RNI4ENK_2_LC_8_5_3 .SEQ_MODE=4'b0000;
    defparam \uart.bit_Count_RNI4ENK_2_LC_8_5_3 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \uart.bit_Count_RNI4ENK_2_LC_8_5_3  (
            .in0(N__3074),
            .in1(N__3023),
            .in2(N__3172),
            .in3(N__3638),
            .lcout(\uart.N_133_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_1_LC_8_5_4 .C_ON=1'b0;
    defparam \uart.state_1_LC_8_5_4 .SEQ_MODE=4'b1000;
    defparam \uart.state_1_LC_8_5_4 .LUT_INIT=16'b0000000011001000;
    LogicCell40 \uart.state_1_LC_8_5_4  (
            .in0(N__2486),
            .in1(N__5159),
            .in2(N__2884),
            .in3(N__3385),
            .lcout(\uart.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4799),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_esr_RNO_0_6_LC_8_5_5 .C_ON=1'b0;
    defparam \uart.data_Aux_esr_RNO_0_6_LC_8_5_5 .SEQ_MODE=4'b0000;
    defparam \uart.data_Aux_esr_RNO_0_6_LC_8_5_5 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \uart.data_Aux_esr_RNO_0_6_LC_8_5_5  (
            .in0(N__3075),
            .in1(_gnd_net_),
            .in2(N__3173),
            .in3(N__3024),
            .lcout(),
            .ltout(\uart.data_Auxce_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_esr_RNO_6_LC_8_5_6 .C_ON=1'b0;
    defparam \uart.data_Aux_esr_RNO_6_LC_8_5_6 .SEQ_MODE=4'b0000;
    defparam \uart.data_Aux_esr_RNO_6_LC_8_5_6 .LUT_INIT=16'b1111110011101100;
    LogicCell40 \uart.data_Aux_esr_RNO_6_LC_8_5_6  (
            .in0(N__2477),
            .in1(N__2727),
            .in2(N__2441),
            .in3(N__2848),
            .lcout(\uart.N_114_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_esr_RNO_5_LC_8_5_7 .C_ON=1'b0;
    defparam \uart.data_Aux_esr_RNO_5_LC_8_5_7 .SEQ_MODE=4'b0000;
    defparam \uart.data_Aux_esr_RNO_5_LC_8_5_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \uart.data_Aux_esr_RNO_5_LC_8_5_7  (
            .in0(N__2726),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2429),
            .lcout(\uart.N_115_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_esr_5_LC_8_6_0 .C_ON=1'b0;
    defparam \uart.data_Aux_esr_5_LC_8_6_0 .SEQ_MODE=4'b1000;
    defparam \uart.data_Aux_esr_5_LC_8_6_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart.data_Aux_esr_5_LC_8_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5160),
            .lcout(\uart.data_AuxZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4794),
            .ce(N__2414),
            .sr(N__2743));
    defparam \uart.state_RNO_1_4_LC_9_1_0 .C_ON=1'b0;
    defparam \uart.state_RNO_1_4_LC_9_1_0 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNO_1_4_LC_9_1_0 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \uart.state_RNO_1_4_LC_9_1_0  (
            .in0(N__4193),
            .in1(N__3530),
            .in2(N__4127),
            .in3(N__2620),
            .lcout(\uart.g1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_RNIN6BL_0_LC_9_1_1 .C_ON=1'b0;
    defparam \uart.timer_Count_RNIN6BL_0_LC_9_1_1 .SEQ_MODE=4'b0000;
    defparam \uart.timer_Count_RNIN6BL_0_LC_9_1_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart.timer_Count_RNIN6BL_0_LC_9_1_1  (
            .in0(_gnd_net_),
            .in1(N__3202),
            .in2(_gnd_net_),
            .in3(N__3477),
            .lcout(\uart.un4_timer_Count_1_c2 ),
            .ltout(\uart.un4_timer_Count_1_c2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_RNIH8CL1_4_LC_9_1_2 .C_ON=1'b0;
    defparam \uart.timer_Count_RNIH8CL1_4_LC_9_1_2 .SEQ_MODE=4'b0000;
    defparam \uart.timer_Count_RNIH8CL1_4_LC_9_1_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uart.timer_Count_RNIH8CL1_4_LC_9_1_2  (
            .in0(N__4194),
            .in1(N__2621),
            .in2(N__2522),
            .in3(N__3531),
            .lcout(\uart.un4_timer_Count_1_c5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_4_LC_9_1_3 .C_ON=1'b0;
    defparam \uart.timer_Count_4_LC_9_1_3 .SEQ_MODE=4'b1000;
    defparam \uart.timer_Count_4_LC_9_1_3 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \uart.timer_Count_4_LC_9_1_3  (
            .in0(N__3532),
            .in1(N__4037),
            .in2(N__2632),
            .in3(N__4196),
            .lcout(\uart.timer_CountZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4811),
            .ce(),
            .sr(N__3972));
    defparam \uart.timer_Count_1_LC_9_1_4 .C_ON=1'b0;
    defparam \uart.timer_Count_1_LC_9_1_4 .SEQ_MODE=4'b1000;
    defparam \uart.timer_Count_1_LC_9_1_4 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \uart.timer_Count_1_LC_9_1_4  (
            .in0(N__3478),
            .in1(_gnd_net_),
            .in2(N__3206),
            .in3(_gnd_net_),
            .lcout(\uart.timer_CountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4811),
            .ce(),
            .sr(N__3972));
    defparam \uart.timer_Count_3_LC_9_1_5 .C_ON=1'b0;
    defparam \uart.timer_Count_3_LC_9_1_5 .SEQ_MODE=4'b1000;
    defparam \uart.timer_Count_3_LC_9_1_5 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \uart.timer_Count_3_LC_9_1_5  (
            .in0(N__2622),
            .in1(N__4036),
            .in2(_gnd_net_),
            .in3(N__4195),
            .lcout(\uart.timer_CountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4811),
            .ce(),
            .sr(N__3972));
    defparam \uart.timer_Count_fast_4_LC_9_1_6 .C_ON=1'b0;
    defparam \uart.timer_Count_fast_4_LC_9_1_6 .SEQ_MODE=4'b1000;
    defparam \uart.timer_Count_fast_4_LC_9_1_6 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uart.timer_Count_fast_4_LC_9_1_6  (
            .in0(N__4198),
            .in1(N__2627),
            .in2(N__4045),
            .in3(N__2594),
            .lcout(\uart.timer_Count_fastZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4811),
            .ce(),
            .sr(N__3972));
    defparam \uart.timer_Count_4_rep1_LC_9_1_7 .C_ON=1'b0;
    defparam \uart.timer_Count_4_rep1_LC_9_1_7 .SEQ_MODE=4'b1000;
    defparam \uart.timer_Count_4_rep1_LC_9_1_7 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uart.timer_Count_4_rep1_LC_9_1_7  (
            .in0(N__2626),
            .in1(N__4197),
            .in2(N__4160),
            .in3(N__4038),
            .lcout(\uart.timer_Count_4_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4811),
            .ce(),
            .sr(N__3972));
    defparam \uart.timer_Count_RNI1HBL_6_LC_9_2_0 .C_ON=1'b0;
    defparam \uart.timer_Count_RNI1HBL_6_LC_9_2_0 .SEQ_MODE=4'b0000;
    defparam \uart.timer_Count_RNI1HBL_6_LC_9_2_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart.timer_Count_RNI1HBL_6_LC_9_2_0  (
            .in0(_gnd_net_),
            .in1(N__4301),
            .in2(_gnd_net_),
            .in3(N__4105),
            .lcout(\uart.state_srsts_0_o4_0_a2_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNI3TGU_4_LC_9_2_1 .C_ON=1'b0;
    defparam \uart.state_RNI3TGU_4_LC_9_2_1 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNI3TGU_4_LC_9_2_1 .LUT_INIT=16'b0000000000001010;
    LogicCell40 \uart.state_RNI3TGU_4_LC_9_2_1  (
            .in0(N__5051),
            .in1(_gnd_net_),
            .in2(N__4242),
            .in3(N__3915),
            .lcout(),
            .ltout(\uart.state_srsts_0_a3_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNICGLN3_2_LC_9_2_2 .C_ON=1'b0;
    defparam \uart.state_RNICGLN3_2_LC_9_2_2 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNICGLN3_2_LC_9_2_2 .LUT_INIT=16'b1000101000001010;
    LogicCell40 \uart.state_RNICGLN3_2_LC_9_2_2  (
            .in0(N__2807),
            .in1(N__3852),
            .in2(N__2597),
            .in3(N__3829),
            .lcout(\uart.N_66 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_fast_RNIHHG81_2_LC_9_2_3 .C_ON=1'b0;
    defparam \uart.timer_Count_fast_RNIHHG81_2_LC_9_2_3 .SEQ_MODE=4'b0000;
    defparam \uart.timer_Count_fast_RNIHHG81_2_LC_9_2_3 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \uart.timer_Count_fast_RNIHHG81_2_LC_9_2_3  (
            .in0(_gnd_net_),
            .in1(N__2957),
            .in2(N__2923),
            .in3(N__3472),
            .lcout(\uart.N_146_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_fast_RNIT1EN1_4_LC_9_2_4 .C_ON=1'b0;
    defparam \uart.timer_Count_fast_RNIT1EN1_4_LC_9_2_4 .SEQ_MODE=4'b0000;
    defparam \uart.timer_Count_fast_RNIT1EN1_4_LC_9_2_4 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \uart.timer_Count_fast_RNIT1EN1_4_LC_9_2_4  (
            .in0(N__3473),
            .in1(N__2593),
            .in2(N__2963),
            .in3(N__2917),
            .lcout(\uart.N_41 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_fast_RNILTQT_2_LC_9_2_5 .C_ON=1'b0;
    defparam \uart.timer_Count_fast_RNILTQT_2_LC_9_2_5 .SEQ_MODE=4'b0000;
    defparam \uart.timer_Count_fast_RNILTQT_2_LC_9_2_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uart.timer_Count_fast_RNILTQT_2_LC_9_2_5  (
            .in0(N__2918),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2961),
            .lcout(\uart.timer_Count10lto4_0 ),
            .ltout(\uart.timer_Count10lto4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_RNIQAJ83_4_LC_9_2_6 .C_ON=1'b0;
    defparam \uart.timer_Count_RNIQAJ83_4_LC_9_2_6 .SEQ_MODE=4'b0000;
    defparam \uart.timer_Count_RNIQAJ83_4_LC_9_2_6 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \uart.timer_Count_RNIQAJ83_4_LC_9_2_6  (
            .in0(N__3239),
            .in1(_gnd_net_),
            .in2(N__2567),
            .in3(N__3179),
            .lcout(\uart.N_51 ),
            .ltout(\uart.N_51_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_2_LC_9_2_7 .C_ON=1'b0;
    defparam \uart.state_2_LC_9_2_7 .SEQ_MODE=4'b1000;
    defparam \uart.state_2_LC_9_2_7 .LUT_INIT=16'b0000000001000101;
    LogicCell40 \uart.state_2_LC_9_2_7  (
            .in0(N__2858),
            .in1(N__2883),
            .in2(N__2564),
            .in3(N__3362),
            .lcout(\uart.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4808),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_4_rep1_RNIHBMA2_LC_9_3_0 .C_ON=1'b0;
    defparam \uart.timer_Count_4_rep1_RNIHBMA2_LC_9_3_0 .SEQ_MODE=4'b0000;
    defparam \uart.timer_Count_4_rep1_RNIHBMA2_LC_9_3_0 .LUT_INIT=16'b0000000100110011;
    LogicCell40 \uart.timer_Count_4_rep1_RNIHBMA2_LC_9_3_0  (
            .in0(N__4159),
            .in1(N__3916),
            .in2(N__2561),
            .in3(N__3827),
            .lcout(),
            .ltout(\uart.data_14_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNILS533_4_LC_9_3_1 .C_ON=1'b0;
    defparam \uart.state_RNILS533_4_LC_9_3_1 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNILS533_4_LC_9_3_1 .LUT_INIT=16'b1010101110101010;
    LogicCell40 \uart.state_RNILS533_4_LC_9_3_1  (
            .in0(N__3344),
            .in1(N__5104),
            .in2(N__2546),
            .in3(N__5037),
            .lcout(\uart.state_RNILS533Z0Z_4 ),
            .ltout(\uart.state_RNILS533Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNICRQ06_4_LC_9_3_2 .C_ON=1'b0;
    defparam \uart.state_RNICRQ06_4_LC_9_3_2 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNICRQ06_4_LC_9_3_2 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \uart.state_RNICRQ06_4_LC_9_3_2  (
            .in0(N__2797),
            .in1(_gnd_net_),
            .in2(N__2531),
            .in3(_gnd_net_),
            .lcout(\uart.state_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNO_0_2_LC_9_3_3 .C_ON=1'b0;
    defparam \uart.state_RNO_0_2_LC_9_3_3 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNO_0_2_LC_9_3_3 .LUT_INIT=16'b1111010100000101;
    LogicCell40 \uart.state_RNO_0_2_LC_9_3_3  (
            .in0(N__3442),
            .in1(_gnd_net_),
            .in2(N__2885),
            .in3(N__5105),
            .lcout(\uart.N_151 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNIAFHL_4_LC_9_3_4 .C_ON=1'b0;
    defparam \uart.state_RNIAFHL_4_LC_9_3_4 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNIAFHL_4_LC_9_3_4 .LUT_INIT=16'b1100110011011101;
    LogicCell40 \uart.state_RNIAFHL_4_LC_9_3_4  (
            .in0(N__5035),
            .in1(N__3343),
            .in2(_gnd_net_),
            .in3(N__3602),
            .lcout(\uart.state_RNIAFHLZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNID2BC_4_LC_9_3_5 .C_ON=1'b0;
    defparam \uart.state_RNID2BC_4_LC_9_3_5 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNID2BC_4_LC_9_3_5 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \uart.state_RNID2BC_4_LC_9_3_5  (
            .in0(N__3601),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5034),
            .lcout(\uart.N_174 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNIB0BC_2_LC_9_3_6 .C_ON=1'b0;
    defparam \uart.state_RNIB0BC_2_LC_9_3_6 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNIB0BC_2_LC_9_3_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \uart.state_RNIB0BC_2_LC_9_3_6  (
            .in0(_gnd_net_),
            .in1(N__3600),
            .in2(_gnd_net_),
            .in3(N__3441),
            .lcout(\uart.state_srsts_0_a3_2_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNINUKT2_4_LC_9_3_7 .C_ON=1'b0;
    defparam \uart.state_RNINUKT2_4_LC_9_3_7 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNINUKT2_4_LC_9_3_7 .LUT_INIT=16'b1111100000000000;
    LogicCell40 \uart.state_RNINUKT2_4_LC_9_3_7  (
            .in0(N__3828),
            .in1(N__3853),
            .in2(N__3933),
            .in3(N__5036),
            .lcout(\uart.state_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_esr_3_LC_9_4_0 .C_ON=1'b0;
    defparam \uart.data_Aux_esr_3_LC_9_4_0 .SEQ_MODE=4'b1000;
    defparam \uart.data_Aux_esr_3_LC_9_4_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart.data_Aux_esr_3_LC_9_4_0  (
            .in0(N__5106),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uart.data_AuxZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4800),
            .ce(N__2777),
            .sr(N__2704));
    defparam \uart.data_Aux_esr_4_LC_9_5_0 .C_ON=1'b0;
    defparam \uart.data_Aux_esr_4_LC_9_5_0 .SEQ_MODE=4'b1000;
    defparam \uart.data_Aux_esr_4_LC_9_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart.data_Aux_esr_4_LC_9_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5107),
            .lcout(\uart.data_AuxZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4795),
            .ce(N__2756),
            .sr(N__2729));
    defparam \uart.timer_Count_fast_3_LC_10_1_0 .C_ON=1'b0;
    defparam \uart.timer_Count_fast_3_LC_10_1_0 .SEQ_MODE=4'b1000;
    defparam \uart.timer_Count_fast_3_LC_10_1_0 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \uart.timer_Count_fast_3_LC_10_1_0  (
            .in0(N__4032),
            .in1(_gnd_net_),
            .in2(N__2633),
            .in3(N__2922),
            .lcout(\uart.timer_Count_fastZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4805),
            .ce(),
            .sr(N__3968));
    defparam \uart.timer_Count_2_LC_10_1_1 .C_ON=1'b0;
    defparam \uart.timer_Count_2_LC_10_1_1 .SEQ_MODE=4'b1000;
    defparam \uart.timer_Count_2_LC_10_1_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uart.timer_Count_2_LC_10_1_1  (
            .in0(_gnd_net_),
            .in1(N__2628),
            .in2(_gnd_net_),
            .in3(N__4030),
            .lcout(\uart.timer_CountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4805),
            .ce(),
            .sr(N__3968));
    defparam \uart.timer_Count_fast_2_LC_10_1_2 .C_ON=1'b0;
    defparam \uart.timer_Count_fast_2_LC_10_1_2 .SEQ_MODE=4'b1000;
    defparam \uart.timer_Count_fast_2_LC_10_1_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \uart.timer_Count_fast_2_LC_10_1_2  (
            .in0(N__4031),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2962),
            .lcout(\uart.timer_Count_fastZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4805),
            .ce(),
            .sr(N__3968));
    defparam \uart_frame_decoder.state_1_6_LC_10_2_0 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_6_LC_10_2_0 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.state_1_6_LC_10_2_0 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \uart_frame_decoder.state_1_6_LC_10_2_0  (
            .in0(N__3351),
            .in1(N__3276),
            .in2(N__4917),
            .in3(N__3762),
            .lcout(\uart_frame_decoder.state_1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4801),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNI9O1P_2_LC_10_2_1 .C_ON=1'b0;
    defparam \reset_module_System.count_RNI9O1P_2_LC_10_2_1 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNI9O1P_2_LC_10_2_1 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \reset_module_System.count_RNI9O1P_2_LC_10_2_1  (
            .in0(N__4400),
            .in1(N__4448),
            .in2(N__5189),
            .in3(N__4468),
            .lcout(),
            .ltout(\reset_module_System.reset6_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNIN3HK3_2_LC_10_2_2 .C_ON=1'b0;
    defparam \reset_module_System.count_RNIN3HK3_2_LC_10_2_2 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNIN3HK3_2_LC_10_2_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \reset_module_System.count_RNIN3HK3_2_LC_10_2_2  (
            .in0(N__3653),
            .in1(N__3647),
            .in2(N__2942),
            .in3(N__3245),
            .lcout(\reset_module_System.reset6_19 ),
            .ltout(\reset_module_System.reset6_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.reset_fast_LC_10_2_3 .C_ON=1'b0;
    defparam \reset_module_System.reset_fast_LC_10_2_3 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.reset_fast_LC_10_2_3 .LUT_INIT=16'b0101111111111111;
    LogicCell40 \reset_module_System.reset_fast_LC_10_2_3  (
            .in0(N__4609),
            .in1(_gnd_net_),
            .in2(N__2939),
            .in3(N__3667),
            .lcout(reset_module_System_reset_fast),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4801),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.reset_LC_10_2_5 .C_ON=1'b0;
    defparam \reset_module_System.reset_LC_10_2_5 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.reset_LC_10_2_5 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \reset_module_System.reset_LC_10_2_5  (
            .in0(N__4608),
            .in1(N__3666),
            .in2(_gnd_net_),
            .in3(N__3700),
            .lcout(reset_system),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4801),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNI38F97_2_LC_10_2_6 .C_ON=1'b0;
    defparam \uart.state_RNI38F97_2_LC_10_2_6 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNI38F97_2_LC_10_2_6 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \uart.state_RNI38F97_2_LC_10_2_6  (
            .in0(N__3350),
            .in1(N__2936),
            .in2(_gnd_net_),
            .in3(N__2930),
            .lcout(\uart.state_RNI38F97Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.bit_Count_RNO_4_1_LC_10_2_7 .C_ON=1'b0;
    defparam \uart.bit_Count_RNO_4_1_LC_10_2_7 .SEQ_MODE=4'b0000;
    defparam \uart.bit_Count_RNO_4_1_LC_10_2_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart.bit_Count_RNO_4_1_LC_10_2_7  (
            .in0(_gnd_net_),
            .in1(N__4002),
            .in2(_gnd_net_),
            .in3(N__4192),
            .lcout(\uart.g3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.bit_Count_RNO_1_2_LC_10_3_0 .C_ON=1'b0;
    defparam \uart.bit_Count_RNO_1_2_LC_10_3_0 .SEQ_MODE=4'b0000;
    defparam \uart.bit_Count_RNO_1_2_LC_10_3_0 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \uart.bit_Count_RNO_1_2_LC_10_3_0  (
            .in0(N__4163),
            .in1(N__4102),
            .in2(N__4004),
            .in3(N__2924),
            .lcout(\uart.N_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_5_LC_10_3_1 .C_ON=1'b0;
    defparam \uart.timer_Count_5_LC_10_3_1 .SEQ_MODE=4'b1000;
    defparam \uart.timer_Count_5_LC_10_3_1 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \uart.timer_Count_5_LC_10_3_1  (
            .in0(N__4103),
            .in1(_gnd_net_),
            .in2(N__3233),
            .in3(_gnd_net_),
            .lcout(\uart.timer_CountZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4796),
            .ce(),
            .sr(N__3974));
    defparam \uart.timer_Count_RNI3B101_6_LC_10_3_2 .C_ON=1'b0;
    defparam \uart.timer_Count_RNI3B101_6_LC_10_3_2 .SEQ_MODE=4'b0000;
    defparam \uart.timer_Count_RNI3B101_6_LC_10_3_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uart.timer_Count_RNI3B101_6_LC_10_3_2  (
            .in0(N__4297),
            .in1(N__3908),
            .in2(_gnd_net_),
            .in3(N__4100),
            .lcout(\uart.timer_Count_RNI3B101Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_7_LC_10_3_3 .C_ON=1'b0;
    defparam \uart.timer_Count_7_LC_10_3_3 .SEQ_MODE=4'b1000;
    defparam \uart.timer_Count_7_LC_10_3_3 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uart.timer_Count_7_LC_10_3_3  (
            .in0(N__3232),
            .in1(N__4118),
            .in2(N__3932),
            .in3(N__4300),
            .lcout(\uart.timer_CountZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4796),
            .ce(),
            .sr(N__3974));
    defparam \uart.timer_Count_6_LC_10_3_4 .C_ON=1'b0;
    defparam \uart.timer_Count_6_LC_10_3_4 .SEQ_MODE=4'b1000;
    defparam \uart.timer_Count_6_LC_10_3_4 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \uart.timer_Count_6_LC_10_3_4  (
            .in0(N__4299),
            .in1(N__3231),
            .in2(_gnd_net_),
            .in3(N__4104),
            .lcout(\uart.timer_CountZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4796),
            .ce(),
            .sr(N__3974));
    defparam \uart.timer_Count_RNIJTGR_0_LC_10_3_5 .C_ON=1'b0;
    defparam \uart.timer_Count_RNIJTGR_0_LC_10_3_5 .SEQ_MODE=4'b0000;
    defparam \uart.timer_Count_RNIJTGR_0_LC_10_3_5 .LUT_INIT=16'b0000000000001100;
    LogicCell40 \uart.timer_Count_RNIJTGR_0_LC_10_3_5  (
            .in0(_gnd_net_),
            .in1(N__4296),
            .in2(N__3201),
            .in3(N__5033),
            .lcout(\uart.un1_state_2_0_a3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_0_LC_10_3_6 .C_ON=1'b0;
    defparam \uart.timer_Count_0_LC_10_3_6 .SEQ_MODE=4'b1000;
    defparam \uart.timer_Count_0_LC_10_3_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \uart.timer_Count_0_LC_10_3_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3195),
            .lcout(\uart.timer_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4796),
            .ce(),
            .sr(N__3974));
    defparam \uart.timer_Count_RNI22NA1_4_LC_10_3_7 .C_ON=1'b0;
    defparam \uart.timer_Count_RNI22NA1_4_LC_10_3_7 .SEQ_MODE=4'b0000;
    defparam \uart.timer_Count_RNI22NA1_4_LC_10_3_7 .LUT_INIT=16'b1110000000000000;
    LogicCell40 \uart.timer_Count_RNI22NA1_4_LC_10_3_7  (
            .in0(N__4101),
            .in1(N__3539),
            .in2(N__3931),
            .in3(N__4298),
            .lcout(\uart.timer_Count_RNI22NA1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNO_3_4_LC_10_4_0 .C_ON=1'b0;
    defparam \uart.state_RNO_3_4_LC_10_4_0 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNO_3_4_LC_10_4_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uart.state_RNO_3_4_LC_10_4_0  (
            .in0(N__3607),
            .in1(N__3171),
            .in2(N__3083),
            .in3(N__3029),
            .lcout(),
            .ltout(\uart.g1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_4_LC_10_4_1 .C_ON=1'b0;
    defparam \uart.state_4_LC_10_4_1 .SEQ_MODE=4'b1000;
    defparam \uart.state_4_LC_10_4_1 .LUT_INIT=16'b1110101010101010;
    LogicCell40 \uart.state_4_LC_10_4_1  (
            .in0(N__4253),
            .in1(N__3452),
            .in2(N__2978),
            .in3(N__2975),
            .lcout(\uart.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4791),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNO_2_4_LC_10_4_2 .C_ON=1'b0;
    defparam \uart.state_RNO_2_4_LC_10_4_2 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNO_2_4_LC_10_4_2 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \uart.state_RNO_2_4_LC_10_4_2  (
            .in0(N__3922),
            .in1(N__3363),
            .in2(_gnd_net_),
            .in3(N__4304),
            .lcout(\uart.g1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNO_1_3_LC_10_4_3 .C_ON=1'b0;
    defparam \uart.state_RNO_1_3_LC_10_4_3 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNO_1_3_LC_10_4_3 .LUT_INIT=16'b0001001110110011;
    LogicCell40 \uart.state_RNO_1_3_LC_10_4_3  (
            .in0(N__4303),
            .in1(N__3606),
            .in2(N__4055),
            .in3(N__3446),
            .lcout(\uart.N_28_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNIGLM11_4_LC_10_4_4 .C_ON=1'b0;
    defparam \uart.state_RNIGLM11_4_LC_10_4_4 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNIGLM11_4_LC_10_4_4 .LUT_INIT=16'b0000000010001111;
    LogicCell40 \uart.state_RNIGLM11_4_LC_10_4_4  (
            .in0(N__3921),
            .in1(N__4302),
            .in2(N__3624),
            .in3(N__5041),
            .lcout(\uart.un1_state_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNO_0_3_LC_10_4_6 .C_ON=1'b0;
    defparam \uart.state_RNO_0_3_LC_10_4_6 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNO_0_3_LC_10_4_6 .LUT_INIT=16'b1111111101110101;
    LogicCell40 \uart.state_RNO_0_3_LC_10_4_6  (
            .in0(N__3923),
            .in1(N__3407),
            .in2(N__3625),
            .in3(N__4246),
            .lcout(),
            .ltout(\uart.N_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_3_LC_10_4_7 .C_ON=1'b0;
    defparam \uart.state_3_LC_10_4_7 .SEQ_MODE=4'b1000;
    defparam \uart.state_3_LC_10_4_7 .LUT_INIT=16'b0101001100000011;
    LogicCell40 \uart.state_3_LC_10_4_7  (
            .in0(N__3364),
            .in1(N__3311),
            .in2(N__3305),
            .in3(N__3611),
            .lcout(\uart.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4791),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_esr_3_LC_11_1_0 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_esr_3_LC_11_1_0 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.state_1_esr_3_LC_11_1_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.state_1_esr_3_LC_11_1_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3742),
            .lcout(\uart_frame_decoder.state_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4802),
            .ce(N__3809),
            .sr(N__4693));
    defparam \uart_frame_decoder.state_1_esr_4_LC_11_1_1 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_esr_4_LC_11_1_1 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.state_1_esr_4_LC_11_1_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.state_1_esr_4_LC_11_1_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3797),
            .lcout(\uart_frame_decoder.state_1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4802),
            .ce(N__3809),
            .sr(N__4693));
    defparam \uart_frame_decoder.state_1_esr_5_LC_11_1_2 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_esr_5_LC_11_1_2 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.state_1_esr_5_LC_11_1_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.state_1_esr_5_LC_11_1_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3300),
            .lcout(\uart_frame_decoder.state_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4802),
            .ce(N__3809),
            .sr(N__4693));
    defparam \reset_module_System.count_RNIP8RT_10_LC_11_2_0 .C_ON=1'b0;
    defparam \reset_module_System.count_RNIP8RT_10_LC_11_2_0 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNIP8RT_10_LC_11_2_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \reset_module_System.count_RNIP8RT_10_LC_11_2_0  (
            .in0(_gnd_net_),
            .in1(N__4582),
            .in2(_gnd_net_),
            .in3(N__4330),
            .lcout(\reset_module_System.reset6_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_2_LC_11_2_1 .C_ON=1'b0;
    defparam \reset_module_System.count_2_LC_11_2_1 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_2_LC_11_2_1 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \reset_module_System.count_2_LC_11_2_1  (
            .in0(N__3704),
            .in1(N__4613),
            .in2(N__3682),
            .in3(N__4457),
            .lcout(\reset_module_System.countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4797),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_0_LC_11_2_2 .C_ON=1'b0;
    defparam \reset_module_System.count_0_LC_11_2_2 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_0_LC_11_2_2 .LUT_INIT=16'b1000111100001111;
    LogicCell40 \reset_module_System.count_0_LC_11_2_2  (
            .in0(N__4611),
            .in1(N__3678),
            .in2(N__4957),
            .in3(N__3702),
            .lcout(\reset_module_System.countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4797),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNI10J41_1_LC_11_2_3 .C_ON=1'b0;
    defparam \reset_module_System.count_RNI10J41_1_LC_11_2_3 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNI10J41_1_LC_11_2_3 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \reset_module_System.count_RNI10J41_1_LC_11_2_3  (
            .in0(N__4532),
            .in1(N__4430),
            .in2(N__4493),
            .in3(N__4977),
            .lcout(\reset_module_System.reset6_14 ),
            .ltout(\reset_module_System.reset6_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.reset_iso_LC_11_2_4 .C_ON=1'b0;
    defparam \reset_module_System.reset_iso_LC_11_2_4 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.reset_iso_LC_11_2_4 .LUT_INIT=16'b0101111111111111;
    LogicCell40 \reset_module_System.reset_iso_LC_11_2_4  (
            .in0(N__4610),
            .in1(_gnd_net_),
            .in2(N__3707),
            .in3(N__3701),
            .lcout(reset_module_System_reset_iso),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4797),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_1_LC_11_2_5 .C_ON=1'b0;
    defparam \reset_module_System.count_1_LC_11_2_5 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_1_LC_11_2_5 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \reset_module_System.count_1_LC_11_2_5  (
            .in0(N__3703),
            .in1(N__4931),
            .in2(N__3683),
            .in3(N__4612),
            .lcout(\reset_module_System.countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4797),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNICR4G1_12_LC_11_2_6 .C_ON=1'b0;
    defparam \reset_module_System.count_RNICR4G1_12_LC_11_2_6 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNICR4G1_12_LC_11_2_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \reset_module_System.count_RNICR4G1_12_LC_11_2_6  (
            .in0(N__4950),
            .in1(N__4549),
            .in2(N__4514),
            .in3(N__4567),
            .lcout(\reset_module_System.reset6_19_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNI97FD_5_LC_11_2_7 .C_ON=1'b0;
    defparam \reset_module_System.count_RNI97FD_5_LC_11_2_7 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNI97FD_5_LC_11_2_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \reset_module_System.count_RNI97FD_5_LC_11_2_7  (
            .in0(N__4363),
            .in1(N__4378),
            .in2(N__4349),
            .in3(N__4414),
            .lcout(\reset_module_System.reset6_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.bit_Count_RNO_2_1_LC_11_3_0 .C_ON=1'b0;
    defparam \uart.bit_Count_RNO_2_1_LC_11_3_0 .SEQ_MODE=4'b0000;
    defparam \uart.bit_Count_RNO_2_1_LC_11_3_0 .LUT_INIT=16'b1111101110111011;
    LogicCell40 \uart.bit_Count_RNO_2_1_LC_11_3_0  (
            .in0(N__4113),
            .in1(N__3615),
            .in2(N__3560),
            .in3(N__3550),
            .lcout(\uart.state_0_sqmuxa_1_d_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNO_5_4_LC_11_3_2 .C_ON=1'b0;
    defparam \uart.state_RNO_5_4_LC_11_3_2 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNO_5_4_LC_11_3_2 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \uart.state_RNO_5_4_LC_11_3_2  (
            .in0(N__4162),
            .in1(N__4205),
            .in2(N__3485),
            .in3(N__3997),
            .lcout(),
            .ltout(\uart.g3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNO_0_4_LC_11_3_3 .C_ON=1'b0;
    defparam \uart.state_RNO_0_4_LC_11_3_3 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNO_0_4_LC_11_3_3 .LUT_INIT=16'b1010001010101010;
    LogicCell40 \uart.state_RNO_0_4_LC_11_3_3  (
            .in0(N__4211),
            .in1(N__4114),
            .in2(N__4316),
            .in3(N__4305),
            .lcout(\uart.N_167_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNO_4_4_LC_11_3_4 .C_ON=1'b0;
    defparam \uart.state_RNO_4_4_LC_11_3_4 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNO_4_4_LC_11_3_4 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \uart.state_RNO_4_4_LC_11_3_4  (
            .in0(N__4235),
            .in1(N__3920),
            .in2(_gnd_net_),
            .in3(N__5042),
            .lcout(\uart.g0_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNO_2_3_LC_11_3_5 .C_ON=1'b0;
    defparam \uart.state_RNO_2_3_LC_11_3_5 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNO_2_3_LC_11_3_5 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \uart.state_RNO_2_3_LC_11_3_5  (
            .in0(N__4204),
            .in1(N__4161),
            .in2(N__4003),
            .in3(N__4112),
            .lcout(\uart.state_RNO_2Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_2_rep1_LC_11_3_7 .C_ON=1'b0;
    defparam \uart.timer_Count_2_rep1_LC_11_3_7 .SEQ_MODE=4'b1000;
    defparam \uart.timer_Count_2_rep1_LC_11_3_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \uart.timer_Count_2_rep1_LC_11_3_7  (
            .in0(N__3998),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4046),
            .lcout(\uart.timer_Count_2_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4792),
            .ce(),
            .sr(N__3973));
    defparam \uart.data_rdy_LC_11_4_0 .C_ON=1'b0;
    defparam \uart.data_rdy_LC_11_4_0 .SEQ_MODE=4'b1000;
    defparam \uart.data_rdy_LC_11_4_0 .LUT_INIT=16'b1110000010100000;
    LogicCell40 \uart.data_rdy_LC_11_4_0  (
            .in0(N__3930),
            .in1(N__3860),
            .in2(N__4991),
            .in3(N__3836),
            .lcout(uart_data_rdy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4789),
            .ce(),
            .sr(N__4706));
    defparam \uart_frame_decoder.state_1_esr_ctle_5_LC_12_1_1 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_esr_ctle_5_LC_12_1_1 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_esr_ctle_5_LC_12_1_1 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \uart_frame_decoder.state_1_esr_ctle_5_LC_12_1_1  (
            .in0(N__4692),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4897),
            .lcout(\uart_frame_decoder.uart_data_rdy_c_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_esr_RNIQ0UJ_3_LC_12_1_5 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_esr_RNIQ0UJ_3_LC_12_1_5 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_esr_RNIQ0UJ_3_LC_12_1_5 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \uart_frame_decoder.state_1_esr_RNIQ0UJ_3_LC_12_1_5  (
            .in0(N__3798),
            .in1(N__3776),
            .in2(_gnd_net_),
            .in3(N__3743),
            .lcout(uart_frame_decoder_N_130_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_1_cry_1_c_LC_12_2_0 .C_ON=1'b1;
    defparam \reset_module_System.count_1_cry_1_c_LC_12_2_0 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_1_cry_1_c_LC_12_2_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \reset_module_System.count_1_cry_1_c_LC_12_2_0  (
            .in0(_gnd_net_),
            .in1(N__4949),
            .in2(N__4982),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_2_0_),
            .carryout(\reset_module_System.count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNO_0_2_LC_12_2_1 .C_ON=1'b1;
    defparam \reset_module_System.count_RNO_0_2_LC_12_2_1 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNO_0_2_LC_12_2_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_RNO_0_2_LC_12_2_1  (
            .in0(_gnd_net_),
            .in1(N__4469),
            .in2(_gnd_net_),
            .in3(N__4451),
            .lcout(\reset_module_System.count_1_2 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_1 ),
            .carryout(\reset_module_System.count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_3_LC_12_2_2 .C_ON=1'b1;
    defparam \reset_module_System.count_3_LC_12_2_2 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_3_LC_12_2_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_3_LC_12_2_2  (
            .in0(_gnd_net_),
            .in1(N__4447),
            .in2(_gnd_net_),
            .in3(N__4433),
            .lcout(\reset_module_System.countZ0Z_3 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_2 ),
            .carryout(\reset_module_System.count_1_cry_3 ),
            .clk(N__4790),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_4_LC_12_2_3 .C_ON=1'b1;
    defparam \reset_module_System.count_4_LC_12_2_3 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_4_LC_12_2_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_4_LC_12_2_3  (
            .in0(_gnd_net_),
            .in1(N__4429),
            .in2(_gnd_net_),
            .in3(N__4418),
            .lcout(\reset_module_System.countZ0Z_4 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_3 ),
            .carryout(\reset_module_System.count_1_cry_4 ),
            .clk(N__4790),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_5_LC_12_2_4 .C_ON=1'b1;
    defparam \reset_module_System.count_5_LC_12_2_4 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_5_LC_12_2_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_5_LC_12_2_4  (
            .in0(_gnd_net_),
            .in1(N__4415),
            .in2(_gnd_net_),
            .in3(N__4403),
            .lcout(\reset_module_System.countZ0Z_5 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_4 ),
            .carryout(\reset_module_System.count_1_cry_5 ),
            .clk(N__4790),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_6_LC_12_2_5 .C_ON=1'b1;
    defparam \reset_module_System.count_6_LC_12_2_5 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_6_LC_12_2_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_6_LC_12_2_5  (
            .in0(_gnd_net_),
            .in1(N__4396),
            .in2(_gnd_net_),
            .in3(N__4382),
            .lcout(\reset_module_System.countZ0Z_6 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_5 ),
            .carryout(\reset_module_System.count_1_cry_6 ),
            .clk(N__4790),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_7_LC_12_2_6 .C_ON=1'b1;
    defparam \reset_module_System.count_7_LC_12_2_6 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_7_LC_12_2_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_7_LC_12_2_6  (
            .in0(_gnd_net_),
            .in1(N__4379),
            .in2(_gnd_net_),
            .in3(N__4367),
            .lcout(\reset_module_System.countZ0Z_7 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_6 ),
            .carryout(\reset_module_System.count_1_cry_7 ),
            .clk(N__4790),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_8_LC_12_2_7 .C_ON=1'b1;
    defparam \reset_module_System.count_8_LC_12_2_7 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_8_LC_12_2_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_8_LC_12_2_7  (
            .in0(_gnd_net_),
            .in1(N__4364),
            .in2(_gnd_net_),
            .in3(N__4352),
            .lcout(\reset_module_System.countZ0Z_8 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_7 ),
            .carryout(\reset_module_System.count_1_cry_8 ),
            .clk(N__4790),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_9_LC_12_3_0 .C_ON=1'b1;
    defparam \reset_module_System.count_9_LC_12_3_0 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_9_LC_12_3_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_9_LC_12_3_0  (
            .in0(_gnd_net_),
            .in1(N__4348),
            .in2(_gnd_net_),
            .in3(N__4334),
            .lcout(\reset_module_System.countZ0Z_9 ),
            .ltout(),
            .carryin(bfn_12_3_0_),
            .carryout(\reset_module_System.count_1_cry_9 ),
            .clk(N__4788),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_10_LC_12_3_1 .C_ON=1'b1;
    defparam \reset_module_System.count_10_LC_12_3_1 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_10_LC_12_3_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_10_LC_12_3_1  (
            .in0(_gnd_net_),
            .in1(N__4331),
            .in2(_gnd_net_),
            .in3(N__4319),
            .lcout(\reset_module_System.countZ0Z_10 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_9 ),
            .carryout(\reset_module_System.count_1_cry_10 ),
            .clk(N__4788),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_11_LC_12_3_2 .C_ON=1'b1;
    defparam \reset_module_System.count_11_LC_12_3_2 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_11_LC_12_3_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_11_LC_12_3_2  (
            .in0(_gnd_net_),
            .in1(N__4583),
            .in2(_gnd_net_),
            .in3(N__4571),
            .lcout(\reset_module_System.countZ0Z_11 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_10 ),
            .carryout(\reset_module_System.count_1_cry_11 ),
            .clk(N__4788),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_12_LC_12_3_3 .C_ON=1'b1;
    defparam \reset_module_System.count_12_LC_12_3_3 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_12_LC_12_3_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_12_LC_12_3_3  (
            .in0(_gnd_net_),
            .in1(N__4568),
            .in2(_gnd_net_),
            .in3(N__4556),
            .lcout(\reset_module_System.countZ0Z_12 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_11 ),
            .carryout(\reset_module_System.count_1_cry_12 ),
            .clk(N__4788),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_13_LC_12_3_4 .C_ON=1'b1;
    defparam \reset_module_System.count_13_LC_12_3_4 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_13_LC_12_3_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_13_LC_12_3_4  (
            .in0(_gnd_net_),
            .in1(N__4624),
            .in2(_gnd_net_),
            .in3(N__4553),
            .lcout(\reset_module_System.countZ0Z_13 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_12 ),
            .carryout(\reset_module_System.count_1_cry_13 ),
            .clk(N__4788),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_14_LC_12_3_5 .C_ON=1'b1;
    defparam \reset_module_System.count_14_LC_12_3_5 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_14_LC_12_3_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_14_LC_12_3_5  (
            .in0(_gnd_net_),
            .in1(N__4550),
            .in2(_gnd_net_),
            .in3(N__4538),
            .lcout(\reset_module_System.countZ0Z_14 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_13 ),
            .carryout(\reset_module_System.count_1_cry_14 ),
            .clk(N__4788),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_15_LC_12_3_6 .C_ON=1'b1;
    defparam \reset_module_System.count_15_LC_12_3_6 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_15_LC_12_3_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_15_LC_12_3_6  (
            .in0(_gnd_net_),
            .in1(N__4651),
            .in2(_gnd_net_),
            .in3(N__4535),
            .lcout(\reset_module_System.countZ0Z_15 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_14 ),
            .carryout(\reset_module_System.count_1_cry_15 ),
            .clk(N__4788),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_16_LC_12_3_7 .C_ON=1'b1;
    defparam \reset_module_System.count_16_LC_12_3_7 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_16_LC_12_3_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_16_LC_12_3_7  (
            .in0(_gnd_net_),
            .in1(N__4528),
            .in2(_gnd_net_),
            .in3(N__4517),
            .lcout(\reset_module_System.countZ0Z_16 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_15 ),
            .carryout(\reset_module_System.count_1_cry_16 ),
            .clk(N__4788),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_17_LC_12_4_0 .C_ON=1'b1;
    defparam \reset_module_System.count_17_LC_12_4_0 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_17_LC_12_4_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_17_LC_12_4_0  (
            .in0(_gnd_net_),
            .in1(N__4510),
            .in2(_gnd_net_),
            .in3(N__4496),
            .lcout(\reset_module_System.countZ0Z_17 ),
            .ltout(),
            .carryin(bfn_12_4_0_),
            .carryout(\reset_module_System.count_1_cry_17 ),
            .clk(N__4787),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_18_LC_12_4_1 .C_ON=1'b1;
    defparam \reset_module_System.count_18_LC_12_4_1 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_18_LC_12_4_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_18_LC_12_4_1  (
            .in0(_gnd_net_),
            .in1(N__4486),
            .in2(_gnd_net_),
            .in3(N__4472),
            .lcout(\reset_module_System.countZ0Z_18 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_17 ),
            .carryout(\reset_module_System.count_1_cry_18 ),
            .clk(N__4787),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_19_LC_12_4_2 .C_ON=1'b1;
    defparam \reset_module_System.count_19_LC_12_4_2 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_19_LC_12_4_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_19_LC_12_4_2  (
            .in0(_gnd_net_),
            .in1(N__4664),
            .in2(_gnd_net_),
            .in3(N__5192),
            .lcout(\reset_module_System.countZ0Z_19 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_18 ),
            .carryout(\reset_module_System.count_1_cry_19 ),
            .clk(N__4787),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_20_LC_12_4_3 .C_ON=1'b1;
    defparam \reset_module_System.count_20_LC_12_4_3 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_20_LC_12_4_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_20_LC_12_4_3  (
            .in0(_gnd_net_),
            .in1(N__5182),
            .in2(_gnd_net_),
            .in3(N__5168),
            .lcout(\reset_module_System.countZ0Z_20 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_19 ),
            .carryout(\reset_module_System.count_1_cry_20 ),
            .clk(N__4787),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_21_LC_12_4_4 .C_ON=1'b0;
    defparam \reset_module_System.count_21_LC_12_4_4 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_21_LC_12_4_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \reset_module_System.count_21_LC_12_4_4  (
            .in0(_gnd_net_),
            .in1(N__4639),
            .in2(_gnd_net_),
            .in3(N__5165),
            .lcout(\reset_module_System.countZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4787),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_rdy_RNO_0_LC_12_4_5 .C_ON=1'b0;
    defparam \uart.data_rdy_RNO_0_LC_12_4_5 .SEQ_MODE=4'b0000;
    defparam \uart.data_rdy_RNO_0_LC_12_4_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uart.data_rdy_RNO_0_LC_12_4_5  (
            .in0(N__5155),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5052),
            .lcout(\uart.data_rdyc_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNO_0_1_LC_13_2_2 .C_ON=1'b0;
    defparam \reset_module_System.count_RNO_0_1_LC_13_2_2 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNO_0_1_LC_13_2_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \reset_module_System.count_RNO_0_1_LC_13_2_2  (
            .in0(_gnd_net_),
            .in1(N__4981),
            .in2(_gnd_net_),
            .in3(N__4958),
            .lcout(\reset_module_System.count_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.source_data_valid_LC_13_3_3 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_data_valid_LC_13_3_3 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_data_valid_LC_13_3_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uart_frame_decoder.source_data_valid_LC_13_3_3  (
            .in0(_gnd_net_),
            .in1(N__4825),
            .in2(_gnd_net_),
            .in3(N__4916),
            .lcout(frame_decoder_dv_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4793),
            .ce(),
            .sr(N__4716));
    defparam \reset_module_System.count_RNI34OR1_21_LC_13_4_6 .C_ON=1'b0;
    defparam \reset_module_System.count_RNI34OR1_21_LC_13_4_6 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNI34OR1_21_LC_13_4_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \reset_module_System.count_RNI34OR1_21_LC_13_4_6  (
            .in0(N__4663),
            .in1(N__4652),
            .in2(N__4640),
            .in3(N__4625),
            .lcout(\reset_module_System.reset6_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // Pc2Drone
